// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:35 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
I9NvoDT7KP0fmSyM7u0wsmipnjIhZGQGTNp6oRoA9cZx/kW6z2nqdeapKuCiu3ar
z/PVMXgpUauwb6J/LVUad/dJauh3fb/SJzf6qojdnFBTCqdi7RoLws+WgE+BlXtn
ufvbafBshnN8rCP66+wSYJb1UueCt1mXrpOcu5WEGvA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2288)
Hn3JQ9KS6rC+QlF8f3XrvLzj64uDl2PIncBxb8cZFBwaeVtj5moNp8GKb5z8FCOC
gy/L18oMiSapSIpgWfiPygdV2578dOs/JjitFaqOPVGipUaVfWk/6r3JA/PIJ2/z
+4S6s3DTATVOZQq02VZ5u6m20UsA/fZ1c/jSpoRvdMKvsEi9VDhsY++ZUzakNPrC
72XaMYq89CQW5lXnh+dSB6Jo+/qH18vTARhx/sY7B7klYQIErDRoWl8cOfPUw16q
N5quBdgVd80GI0qX9Fw+6AtxNeZNjffuXywo6yiaUh3t+q6nuhomoLbW1DsdY9yX
F/uwqStlvJKZ9Pel3TMk9eUu/nSnWLQHLJyISvrHxX17xpOYx7GpXR/tEkUz0psL
8RhwU6Tvpe5KQgU+6FSCcAtZ+h3f7CsOy9BdMIev0mPGQnxtsuUrvQrd3RWoDs+3
BBExsxDe4jVFdzD4AulWhTA8SvkONtet8xG3O81dVwsSrSCyVJ0UOWm7pKOYjgj6
bbITe+/FSR7FE2n7Z0cMflrRomAYBoKoJA6hzHesG/DIu+0GRs/HUIf30VBXus+Z
t30N9ayHyNNtXkiXWMycpGsNNicL8973qwkkk5uoWhYr84hrBcD9ozzzwwMRWDKG
D3Lry1Bqge1Afj04lHQpYL7+Y7wR+VKsR9KMpBHS/jHD8nNANBRDK0ZzqILOpsHe
10JIH9glV56LGeiko5U5t7bUoc7PLp6YO1eoxHHHh7RluLRcJ/zZDc1gIrfiGVsk
5KpepMrB0rQF+rJg8kcNLpXsYHZbdSRSjNjuH6noreGw5McNfAwuUR/85k463W2u
62JQ/Micf9azHYpFor6kT3vdMW/lw5Je4QFNH9YeZG+PVY4A9a0IMfDGpTGpjXzX
sZw3QejZBZ4Vqg6V2X7Ab/aHmP+xt2vDxjPoeocEVPFjdcA8rWuuOZPe8qDMt09y
y/xVK1Tt08IyCgvlYk7aEstFiOXuSKm7uECWDQCW74qWNNcPaVMPu3SyawLaWClM
3Cq0HZm6JQRZIbTv/oTTuEbCU6O5nKoztF/4AmCUreXNiRNs5nNtqgQug6W8fbPU
Mjhge8lFTyGkfhmkGlZDEUnFP4ZUwyxR45ZTi3Xg25iEu41pIzQuIn1HdJKt7cDT
NHtRYI4E4Sf38itPa85T1nI0JWPXbinuMQ1cL4fW8M5JZBXybb5Y2M8GXILhITc9
8Ge/q3Au9KdhqIoBtAl+Roco+nFl5r+J5hpslW/NX94AkxWRfCZMJlq39ZSagX/x
0yFj9WaOsXspayXYe371gL8hfFcR3oc1AciuOzTi0r8779F1eL3/fAXWf6IxgPOX
s1KDtx3A8gNx0b/nbwtPIIVK1huPBfQjquV6K+zOzl4jqlWaKzVc3VJIvgMxQXf2
uHwjOsQ9R2+aYnDdH5+ByMdIUte+twLWYqA7IGut1UZuBbTsnGTixt3FKexlj0fx
oFR26T31Jb7extXoJubfNz/3LNYuOKeCKrYZDT07GZFPZbLYC8ad5Tpfrqcdpou4
sRXM8E+oBErTb/9M9d52K1uLyE47EnHIAh7m71zBcnfG11ZmKUhaFIgzCE/UoH3o
aqbMnKcApvLr9MHO9980MQNaTEwwYJC6T1nftAVR2NCg4mwpotyCDB9vjDFPOJDH
zG2fkl4tI1tDKFxD3fdoNB+7iMtMspatXq2Yzo0dqqNZMRXaGOOMMt1qv43bnmWI
aPTJNOa2PbPLr00I4jTIUdDZmcc/z9myRlS3Vv3jbvtmkW1MG7/XWgOmOKMkoVvG
7V3zGducAtuWDNoVAD99+ZeQzj+riQGSGcO0RSqC6puMXu6AjtaSAFzPVnDhXDLV
jxekZ4GuinvtACjKY//dT5b91fMBUe+UVEMVJk6YNG01puaKw5DWUkoW+302c733
UCL1Wg8D8clj2pD0ePcb3+KMertIYsz9GcqQOTWdDEz3rm2QMsvuTVZGVRpYmQoM
736Oi84LDDZfE501KpqURaaZNY+TqilGYc/Rrr63FqyongPMoK5hM259fy15vdQe
GGOcNDLmttpeLilf8BDImCIf9QYNW5INVs7l3OoczlGrAy/xqB16oqBln67kfz4e
Wp+RyGDWmKHHFC2d+kuXvWhL3hW0Na/xpBrpeksamxWdgtrYaNkLt4lXS2Y/Mig3
D7ohgijp05fKZuR3tfHMcRJ/WF2PFkcHnsbX/+p4D5okIizUowRUTQbvEz5wNIpc
x7ZIdkIzy7ALQU92BwRDIiW8SYtfCzanTfZDpGkPsIj0gDpLlz8CS3L/+vQbuY9P
3hrTFWWvRfi4w5JPa5+/E09YexgCwrXTc8nfuk9HlmqteXK0F5e9YTBFwahG2C9D
fORbThc6wF2ef6obscAhkhb2yuoDbZGupdJGf9KPXQ8W98Wa8n6QoeLDQn75Lw0S
F6z7p2MOQkf+Km+6AemWx60VF8lmR3ZIF4VNbg6DXVsg9dbjegvYT4lLWbLpp+L4
OWQrHDICz6ltZzmneLJ6KCM2O4SkF1IuHMINAhehsfcEKU2X1Frs4v3BkiG1fcLd
KUKyNWUhF1tlMARI8MCu7Urex3BulFDyrFNiG/TP+EKFEGCm9qbchWWJu/o3qCqU
woU11keAIuNCQHDanw/kkYxKZ2Hq2i1U9/RZDEg9a093a/g3HXv6ksZ5dRLLQXny
NtTiGxxIIwpz4bZ1rMj+2IKo6Jomr7SxuhGJX33HBiTmkq/JlboGPB9XgYWvAxsZ
u+n61P9VHijwr0VTx0pfbY1RNyMFxDZkBBmb5kb14++x3MEXpYt+SiL6qRFmX6vr
f29juXiseP5N/3jin2FcDDA9wLqqakYAsRiv6goGypy32MskHuABX1pK1qCIMMar
eeejq3M/NBePzaAoPJvwUi6bamzudt5L49Euvhvzc6f3BvzFFMFCkOx1Ba5P9qwF
VvgAjlU48hGzqdYbdqAn7bbFmaWSlKHSTRk9YTx8qhZeGWHzEWnCZ+pYCb01oBfp
Cdu+mWz4LAGs0Fy1ovmSqitTshbjM2zbnnGtOuL7Ga4=
`pragma protect end_protected
