// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:45:24 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
q005oDyCDt22wmfAW5P/ZEHLRQKw0ZIrkSEOGHWir9fUPDdczwbMZ7PmKIEkJUuq
o7Uk+OnCIXUkaZQTXcfZHckohojlLhVgDu9PdFyio6A3/8clm9Wy2zFRxVGRhFfZ
wATbOOuA/Q4+rUjQBL6AVF1lkqcw7svrXZyUQYe8xZE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12560)
OM4Pm5jYl9V+ZNN/tkJf4Z/8XFZq/KUBikzqh+ceMRzRuDTijjUWyWCxBYt6NZlk
xN/YUDgteyD4Ifvg9eW8GrVgEcvi+voXGQarFwPKoxsndw0oq8f0+LhlBc1jQA/j
euichRFux12tghyW5RaCxfwiFkuy4a1SR2hS8uV0AaZCwZXysGzVnQfbsXPPJfnQ
JUM+ZFSQMlPtVC80nNViGVmYOfOhNPoOK35aEkCIiaQ2NMFvYFouN2Ui5VLASkn4
SHt9qNdBCRjcVELMBUZsJB0orB3ACrqKF2IKt8NVeV8llvc2ND+clcBaMp6mK2KM
p74HKuysO/5ND21vlkcTgQCV6VckaIPX8J52xoAMlJhrESGBdBM0ch9srAAq8dla
6yeoKt4Miw/byC9xjH18M8jgrjILduT/tUxsFmgTpGJkm28Mu/C48kxb6gY025qX
lnz6do9w2yF4DxFKM3Qm+peDJLNQ2wRssfOgx0SVUsm5JACowds8bNbQTMxbbG1g
6g+RdGIvpIFPY5dviJoWzuspYu7cEaxBLA+kXhXa8a0UINY3tOPyV5toK/m+bWZJ
P/ogiDIJpdRynDQTYIbfLfhIXF9dWWcmfh1uV+Hi7nMHdYOzcne2r2lqR/62qZ9k
tp4EaGOCxTxigUYGm1rAIzqLrFknRT2ee/8JMsMTyZqY2DKz4h67eQ1hfGECZSk/
FdQhMELNToGk5L0FJprJv9mFP8Sn8gNaBaw/YBoE9Al8Ri9N8A5K1ZFDRwwxDklS
aV5VCd7nNH5JRlj/HmlVC59qkc55Qo6ClDqkSx34uKOv5UiX+5oSa45TTKKe/a/W
ymHVMjK+mqughx+rkuynW3+2iJGAxihXdjYTPJ0br1ZVQoqyXiFBtkSZGKCZm2hW
7g9FxsIKYVCgMVHxCgSDqrlC2XI8LFBEd+oPQwVRYRbR6d+m8c2ryHYrpjGEdIhk
Hc60/G6YtZkY4W7aOdBpklc+3q1vpq/lRCXS+clFE2tqb2kRaCql2DWfXL+w+GO7
kPsCizasPEi/FKpXWvTJlORRle4b0ZEA0vTFsbyW+psw4P4nhsEyQG1SSlnm9x/O
knDZhC7nffrP+/4Hc8gNzepkbH+1ObqJxssBBNygxuaTfOThF6K+DNTNxX0CfAQT
pmLgFNuIJKs3CZLRRfBQqky1mEuO/GLkdzPa1OKTIe+TIN3IOua+GEDy07rIbFjw
Uo+xKbIWWjwB9k8kV/ym0o4Yj1Vtj2i70vzX1hJd+P63RfST+E617bvNYPrdBycy
g19dE9Q892HpDobaWE36DVTQUejQHbOd37FZCvtfohabnNoW0kz5Du8q39DAViuz
6tK47GqVQbpRqRdYkBXdi5DqEGcOw8jo919g1O13ROV0/Ol4hXZVPaGCVeioMW8i
mVWNP5gDGonm2DLlTajxDOqcqsNuEY33/SZB8eFfVNzTILCENLF9Jj95UibrqaeX
xGYk/cUazaTvDcBwrPiPT9y5L9DeWbiBtRyIips6yDqzf++1bUCfjn19Y0aLYZKt
6rVBFLLm18cZvC8jngh7GPaJqTU3rEUk0UgdLi13hA+6n+k+Z3e4clt7SgvZH7Rf
ErFVCip00teVDPTyvvyeRyRsauXbzIY4VxwZDoFZdZ7fB1MUKk/HJEau0sNN0zPU
tyKTGd88cL3tsqVelldud7AUGoUA58T7H4rx+IHtps8zYqJs6O1yBhx2GMgh+Og8
PB8cSF55kWx9fukNMk9ojnLPRe17pGGuzy3KaOgpJnlbGWmpRgJRTvORxgJpowhx
6iO5A/YzLLlndMGJzTqhi4YgjOnTAkT8fz26RDFs67U6DGvh1r99S4HYHLa3lDoC
1OXxXMT31bZgNOif19FTUrqSTMg7XCZDGnIj6Tu98U1Qu0P52dXL3IL7+IjnutQ/
Ky5yHzlhBhszDo3poF7klu/XOL4A2yWpON6OFSgA1J8VI01f9FUWilzhA+8oMNeU
TS1Gn8UPAwgIDfiyJZxn8+2J5sbKiLdv+/hTifIBp3DenMr1FVqNo+a2XL/akv8W
oKOVm/hHZyhsorMwFJmOG1xbaGc35vBiNjQrbw0jj2AtD3VIR/Z2nh6vdEheR8XO
HTwvMW5SzK1t3alcp/ci9VV7qKAF+7auHevILYWGqW/0yM1XpBb31nNKcsriPzeW
gYA/Ql3PLlNJ9C2FCoaOIPorC7p5kgVgPIFJoq3xOL1kx/eCt+9GbFyW8c1yuKUQ
moaOj3AmoTw6Ya2DjNTJu3B4xusgR1+W+MuuQT1wDCBHrcpHOCXx1sL90/RT4+7S
MuiopJ+Zvmto0ydBKUkOGYaIuDP3kFXIuybqrntCh5WF4AgAh6mbOtHcn+zR4zBo
CELtc6VluG00XXaYjla+DA9XkArWNNQr6mFag8vMrMXLKRqvzPxqUEarKVPDMici
gYhgzAuO5CM2u1jmgvI8V3iXIr3BZVcQXDKDrMAutuhGE/sriz3e6aJ5ybn3UjMC
UJcUmAW94NSg36TG3FKHL0WTAKc+BBb6mS1JsEmdfivC2NxcEocF5VJTDRMerUyF
CN6iB46I+OPJjpQGM15p4IvoNJBBKli2CDHagluK22HqSs9sgOIigaov4OdzSUKV
GkIYqubDxMc+NmNJvqrDoKqoQ3vka2lXFUcHJqPMvNlvLhWAf/pJTTLiibZeG6OB
9pvtm/u4RgRYoO0q/CWXK2mEeAvV2oN2qSgxmxstIjgcWDGs6ABH7SwIhwg6YxG+
nNDKdRfU/qiVG8lEndOwB8l5fYrkO0ln6o+mo3CRKbqor822tUYHWle08hQwhLi3
DlV0gY99DOLlMSSleawmPWpGCJMWMS5ByGBbnaMRALjyNqZv4VHD0J9op40L7sJ4
ioEAy9c26JVQOkGFN8o0UChLFnWKLiX7CMgFWmTsQAsup8bvWmsoEIhxxLqUAImU
Qix0hBWJiy3t/oHaA8wJiwDlYNdkPWCqa9aQ+smPH27i329rMheDpcsi5WkEs0yJ
SZ38NALnhiWlpgT0XHr0w//xqnom1RDs9sTbyfXBYM6K6baV7mF4ySt1cZ00QA5H
uP7X9GF0A5Fkz8Y2tHWGcNAZUkJBV9DHWmXagBmhmcwQttqIJh9hz/0FM/S0sYhR
PqZsKugyTXBc7RPiK0sANyq9EcNjZQwwQNwWwzQxDdhhzhuBKDuN+iWr3s9zw/5X
+FvcBDVidquSIlPU1ntFR2ZxT/v0/QXqo1Z+DjE8lb1HpCWRypeJvkbMl0/uZNMp
QD/8hfi4wjDYOZYawZFIcomDDhtYeoNGAl5QJAdoAH6u23NZwDKMn2WHCVTNhwjl
f35vj0Jdv2pTnKWugxGzb1asbs5Ob+FY75CPo4d4RlZ6THRJ/qowr4KSG3yQuZ4J
yr2tvmAsVuEwOBRac7VJaw3qAYmjWByI/oGS6yNQiAaRdS/umG+9ZpYfvh6NXbC6
evL7hus9Z2Dh71Z59n6BPwP1EYhCqtARGna//LIzxpgbCEL+Am9NnHlJOKEBDWIZ
YPWnkT9NIbNhEfPRPnOWvImGA8yJRaYu562fw+DuO6E3aRksAYdZ2R1D+xlHtiF7
qEeRqe5nmge775U/PklfdW0dk8akAZ+ZgdH2IgVuh6Oa0m8NUVdescCa57BKmLat
44E7KmE6N57+LTiFFPbxPHveba4jeTsuSlLoNZ+S9VFQyf95tsAE/ESG00oYdBjx
PYVRiOYYSIk8I8Qlm2Ch/WQDIKMhlAll79ygMBiJpLi74Sj2fvf/KgxB9T2+ZfZp
XmNIrCnYL+I7BIjjIj5jshTyIXW4C7kR6dhQNklk+19DoZ8bw2B9WRIIUvXDw9oW
JCFKd+rL1jNdhKkkD+U58mTazGCkZ+8oxJfJrPnrFDjz9npsz05IkFnqql5+GGdN
DZKelbE7+Iv8ywXXacn7YrF4l9LQfQLU4CwZUAO4Z1J3fj/ZYNowdYko875/u5Dl
mvLahvk/CkBKBFOOOu5xD966wvrEDOLuQMbgALGPC9/0z0DMtZ8gVlWjdLJqx6ZM
aQEwVlmwtMKrXnum11T0IQrSBsg8eE/5dW0qJ+nSebmn7xuaoV1qaHogB/KMEzyS
FaOkeUitQWwcCgSzJLvjGZqHKqbCtB1rRKDjDxf1usTMG24Nq9WR4Ptgel9uVMRN
ZG/TCXEl5pdd2mutah/97GjjiQfOE8bbfeedPIpsizTq1RRFTaJC5Lc5rKrmU+gI
LSxsrc80XpuIJp9sBeRqn41aSU46IY+nwn1ZDN0tOD7+3OFX0kn44icO/EO55tcA
z/HCYPR3qunu8vE34cfVHcEQ32H7FB+P/LxMdjqWNVuLGA7fS7Xt74A0AuJ3hzgL
nwit+IaSBPdBN70wlsLkFGGSC2kBmBwiBW5yFhTE3gsGRmVE5yjUIA8CCvFpsm5z
Bhh4ThCR1r4fv/hjKTrf1kwC7v1TFu8Appsj0T0o3fafE9G/b3SUmzMuAvQLyIJU
wZ1+Dj5xb6TUoThXQYnveP6cwb9GGhEuf0HNVSTZ5KgWq+MOgAzhwxRoJIfjeZm8
AkRCZC6k3gEHTh1HjSxmDOcKqxLQ10Vtl4evE2XMZ7YI2x3yUZL1y8JxZEgxbAXE
Ej081lK3Sh65xiKaZqfVgDu+kZa9KM2llQ0v43/OU/VeSFYQNRBvTmFUtboHXmZm
3wDfWgmXBEKUL6/c8MM1NydYOoEDZ2DfxP5Y/Z69UtMMjlDpSs1v/F2VhG4rI9qL
vSKk+Cm7GnSLkGk+p1+3rdTbQmkQVxI7ljoZ56kIKQpkpSfhOIM2xpBTBUS+eRMn
jstBILUdgyC/Nf2EK+qQohmgL84cqF0V0Fl34Uvz+zlPzHcObGUPVD2j8yt0i/ZY
7nKbO2ORbeWi3GUWQEeEpwjvqHjmWB0OqqdL6C47eM0885jXpRvvZ3dtiYDuHbAJ
MmSkYTmm6QfzXaf/ognjuWuv6Fk0uVNwaI4TsI2MrvFvDGiB6l1+XZN+CHuasN1s
E3MLCKY43fasGTQEOlU3jPW1jrBUB4EQeoc+somQHZQtGn1lv4/IBJSEGFbrvhw3
OEBapKedk5AuFCOCYHkhjmEOF2QEXEYfH2VCjYHCog5Omh6ysVLqMPw6CRaSzKwn
KRLzg2vr8eRIiwlRArl6zle6czVnunlv1+xXY73i5R/HnzJluCNLbZG6rUqch/C4
Xl6L16VpxWe91bgpieHBlMCgZ1ulCOMwgUYC4ZXa2lUq6FbUJuQUoQHwMgv3RgG1
xOb2IcZCLeSUpTZmXBUxg819hozNkQWZG/rPGygWPSuKImL5lKZQlZPiZ6eXqfW6
V8RyfB8oAjGmvJp1RhXZKc2TJh3W4pCMp846oe3ZZef6LXP3G0/OcK0AgpiJQ4/8
/CmyyNPS4g4vPKmBnTeKWaaGEw/Eo4EAjnPsGUWMNmNBqjyyWg4KTUbC97cMe8YA
SvwX1bcJq/n7DJ8/7Nbe9DCaas0bLWbRVc/ekrw/YzQEoMZ+KO3/6pCM6kOQjFPy
QU5d6g3AVdNY/bdGzDrIg2k+xmOd0429tDadg9jZaKJ+hMf0pF7oPuMitTO3YTRQ
Z6jnK3Pq330u6PVYy4a2uDRTw4UIB5nV3Sy0Xlb5DXiUskaDjpD6UnhmkEwrkM0e
2m7oPQZz3lemc6j+UphRw25FZVrorS7tEb5tUrq2X6Q/BJ71gZlhHjFiUcskoJSJ
BOny5qdiwduc2B8CbjYS98PDD4yuFjG6oPKY4SZHHG3yTPX2lYyLAv1cGJ+mT9/5
oEmABBL5sVm5WYS7UKtnbcyt24df2LleGEvEaNSp0FIcN5OdzIdfcS+KTS7IlGHW
oa+XF/0Ppi+GrQvmeruioZe0S2H9nx+fdmn6IuPSMFTuar/K+FALxOqQ0HtauE7T
E4M1RfOEvy3aqq2LzspkhWfZUTEJofVHXA/2yAd6xakrKdyVNbiI+5i6zQoprum7
S4V3gxufshSch4iV11V48buwyQjWrtnCjDLt4z3RqaBge5FYBpzrZ6c9EwhQz9zw
ALwyFPimOs4/F5Ih5+boa3WEVYtvCZHXw4C0RvlViNk70BcIG3A4do2n/Y041wCg
DDY+bCSDlAcDCn8SE9v9LVKIe5XfEgQTv3onkofbw+tVHyXFrMA4gTFOjlPLQWQE
KUhOMj0EKVciwUjUF5ZZQH6cQyV3x2TTMzvsyXqzG1yCzfmDk2GuswNAipDNVnsg
KQLP8lQICnF4CDJOvDXgaJRNvc+UeLXodrV6lhUv2uESor5BOLit0cZfxsZ+R6Vj
vszH44luR8IlekMhmXnd9+KahduhHCukSrhBIP+eNMX6oaCcV+SKaSJyJaFkVR6f
MvWUxDz/x3GuGexcGYWKPNujtijVJlDFCDq3CM65uPmJaSsC28Fy4NrKNHdCq0/T
zuRLwhTAB/6Pp1oPC6Zy2Fcg4ND++cG6o2xeoFpT8MOtzNowg9sn0uVLfksIrjv1
Ol5cZqAFdB/LeKsO4Cfm594zRzm39zemhNS7mmvNL0sngF5nreXrY93mNeDhyR90
kjhTYtS8EHN72/T0oioVhciOdpD6v/70nujcQrfdtbj/gWZ3CqEfFnNSBlmIFUp2
3pDHh/8OHYB5d+Xj1LeD+kDIXYe+dvigoPumBbLyPm/O9GlJTu+S/5r867OO/QVh
TGoEPFSTkH/69sJhZtTcGPxw3x9ZUMJxRT9YDehdhG+tG59zv6+8Y/L++1jcuGrj
L93AgD45swTOCqbT7QvCoZ1q+YE6SiUkLHhk5AUOdEyTVwZ3AhxaoyiPIFXx7uw7
heEw5MgeLVyciu61ZyBBrzirpXJpT6wGvuTN1MSy3V+A/JQVKs69kxvtMsXdaiGU
Z6gd1/C2KK3uEhBniWNNyaaiVQdAzKoDeRvsbLJpujqj6M1l4a9y0XR2peXFjqDh
G0nznficWEOKHXWDGTChq3FDsFGyGsI26k3FvSIbMeI9jZPoEKKt24SH+k/8euHe
hfUTp6fJdV9Y/64UKGru2KvuVCNfa+XPRFdFcTV7RfU50QKQFumpoIu4u3NNUkQq
A6Y8bwumFHx6TrQ18ZYkSfgnug/3CiZsHZJ/0yXu1qvHVh1a8KzWcSJn5BVewOMO
Ze/JbBAKVD2m2V/nW3eJp7Xhr4Mk0fn9CofGe4/N2+u3OVg8umzi44YRh5v8GLN/
buleIGVue269oODTzOV5Gx7y5vl3QeSm5oJTVoqmL5rr1nziLL5gNcYvAJOHhB2p
quxmG+JyqS+k4pQfbNpZvrVRVV7vE2nhWMMT/Yd/tDux4CBOjB2+niOCmMBPXj75
sNKQzIQ2ys4guaYsfuiBjHb0OQG4g0/VrJ3NXyb0E7llot7HPYAP4aNnsKF2keSi
iMr4H7GGoQJl2txBdwvl7/C+V0wxoqQdoL31jHVYblP/s4oFB344g+bI7Nywd0NU
eee2EfKn6WfB54Q2cYvHvSNOKjPEEnKGHXd1PZnZMYB6eZOG8g9R8nydrSdmTip0
I038uY0d78IxeZUebghreDB1pSN5S8YXivQQaT8jZ4JGDb6YOu3BNoaX38s/eqSj
oVBCe8aJ+senEFtAqPHad8Zv/3Xc1NIu84IeRsTD7lKCsiFEPGbQtz9VMlH1awyM
xmiWGRoNYTDO8MDZzWcf1W9Fxjc+NHvxen2NcWtFiWNxTFrE70fwQbCmzcvT0CXy
KlHjEqhKjH8AwCs6M11eq+ebIvIP2CwEhJBgdewJNpg55EOegfQ0+WFFX4bLB9Xd
mh76dvsuvff6tXWt6fUGbtAq14Pq7bsrdbe5WOcUn4yfaeAsk2LA2ZPPPF1GPtDG
LreK9Jf0FelRJGgK0fElWtLzVpvL96phkjG3X+a4qKT7EX6u1hTLLmmTjsZG28Op
Dph0RM7w1OEdEtmAPdSlKcscj1LwLjJK3EW2RfzqBsXlUGCIYZPEYWFpfl0yy955
/AEa89djib9wjpyo7163pTjIeFV1bAElWStKii11BzWDHXfA+ir+ssWTfTgWl+L1
rDsjFPfkr9qLCZXtmFfAFG1Sy0KFLnYkOVnlBJ6DTdvoO2fzTatjfkLrMVmnnPbX
ImefHQdXtxKlcnnMda0BnYfM8P0Y+s+ENuNq32JM1AO5V+oXwd17ZYTWa3eZD9TY
O9vFxhHGMXpBRPxGTNaWyX+1wb/7zm226gAieWxR+YhwCtEfoV80QI2ATCrvCdDL
mWwM8uBMWPq4Sodfhk9EnKCao7onytTtsHYEHR5Y/Qqll9SSnY8zZrMxOTdKpBwp
NxLLHoM2zH+jNgOXEFYbJ/nsO2m0GRKYYSr89V/m/ZgdS1lf0UP6TK+CTuCOaE1a
rQOzpc8gQuJnLt6Bfl7+PpTy0KyYShiqDAneyyTjcjsDqNS/sSpBEZQYClbJlcEm
5MUJRSNhNfuzJE+jKx8MjeWq+D1U6RnKQFSqJ0aBi8CTW3nhgnwLjVUNWCkS6ISO
jlWQL9U0qc9A614WffNmmfbhInl5h2Krvf+simU83m7Ga10NPNromCe265L3MTJy
S/Cd8MzuRRatR3ePib87XN0ThuE263O2Hc+Pa0a85HKheohkk9NjmrXSRgdzBUGg
S3qcpDmnMeJFDS02trJUQmLBelgD5giB/ltQGFwRsmcDgv6ev33hBx6bd2kXd4Nd
wdR/sOIviiB/ECmikLH12VGezNuhl5qt3q7iOx/KyiU2nBqdPWwEN4nmV1/DQmbZ
Uuf5vb9kM815hut/Si4rk1114Pz/TQNyh00zPqkOSRpL6vWsUXzxe8HTNYafglKP
eCs0gZU0GuI3flKdIhV7U8GzVlHW4c83UnUDB04xEm1PlkmQRrZgRiT6AzEXy/Jb
Y9Y9izKECKLYq962J5fZ4pf0nz2UZs46Y33REZBVMA/4xWG4q82ld02rIki0uNNT
5/AYhPUBvg/TRS/3Eh6GCCm2I9jH98KtRnbWjl/VQ+fBrI2F5rB+ac5oV1JbU0m2
ZJUhbZp7Yli8NKuOW0BjWD+Ca691bbodvgaFnnQgoZukOxoLpJaGmVZ6m/tbyM9o
iMEWkP4eksv8q8oZr1upTWgo31t8lh9Quuw/4incGkiGm9SztK9cy8f/1sIJnmbA
UpqUH+d3QGY7AonuJQjnuMFOjieyqbcqwnUgTmiyetzdVO/fbeR9Cz3h7MMrJBL1
84u25B+7RmaUvoPPGGx3gwjfFJYdSQNrpiDmAWynfkGnfrmjdLr+i1rS+2Q/LY/W
H/g55CJrmIkSXKw855+PjszWdEqQPqyZWh13CNDOPoyqb4v1FCOLUiZLsQklhuBd
TxMM1j+/QlBaaSYRwLnpDWkoXuXTMfykqywFJvsvoG4TynnX9dDIDQc+6uFLNxsL
4gOrWPOOI+wIhm7AM9HpPigaBVIqy60iqvx4rOXIYkzJuKejlv16W1pkbdbTCi9d
4Tms/88Lkdyh1kFvCyjmZUkTSgWYLODkYNlcxffVjZ30iROqxXIvkEbS1VJqCT2+
bheFLHxnZIfHMFgxrXhQOIQKhluRE9hQmZqE5AwolMS5fbnpF/GCMDH4mT9zml5p
IPVVlKB/5aW4Y9wY55sTYj8XYsnO0FiwAOzKZ2o1sQNdO3wiqpMOBYd7weVWmMRF
Qkk8EJgAqfzLt1mwDvBGTGVZ970yOkcf3kn+O0C2/NOTOegZTfofclTO3e4m6fap
tvKCNDgIOnW7oQ8C8UwSOyYLpuQXcA9sRgaMNM4+h6iAQ6ULRxL0GZxw3LD7W5xY
TPmHaocryh/RyFyCsZLsrLjUUY+2MNhPwNtIbIBLwbuKL2R5fbfmaiBVkvEd4aC2
s362W+ew9wApMAZyOe9voRtPnAvwn38iXfeUrUgNjYhktF24K4kKCcI3NURr4tkx
gBIqeTHGRIdn+yr10ofoN+ih08/8+3UZLE+0YRXR6HVe5R9fHLWv/w5Wrfj1BUh9
0U7XzP/WSl/EaGGE7XkKcy+TkehoC5WS+mjQy1MWG5i2lHcS/MReeipkQYjA82hf
CaO0IX+cPP9H2sHBeJwUdXMwwPyrtBEHMAkA7i4RJBJQE22vtGTx9ZxWpZ/Mm0T+
mcE1szLPaWRmOxCZUHr05XDTOVfJKNZoNrg7MvPs+nmCUjIxEqdKjL4H7Gjx9gcz
FvzN7Fxpg75RBZ6fkr5HwmY56R00gWBVGH9fXe5I/Q5DKJTA+xbDY/t4CoplCsHt
3V0YIgIgoy2gBVUKPnTOZquKZZ0NAMiq5wxUkiVqaNmoAXmYfWAnN4HvDhjt99u0
Ad+T7O31HEyFNjJHlLyw0XzVC7/eWw77dChGXcREdtW+us0grlS0e7WvkBxKifqh
eKFhWMJ2XNSRH+QyFO1U+f0V8HJEusvI0CMO2q207hz57/cGEeqlX+3/rzh6HH4F
TFDAcm/UIrQsPxMN2BGtfVZQ4EowgmvOvZJGD9e13hkSuKbqCNsdHDh+15SDMBZX
2mGOQK/Vcexpjy1v2drB4SyLrPSN4mUVp2CyWGqM2HmCirSz5Ru6wyeja586INz8
23S1koG22Vmftd8lmade+7vsJ6Rw4BiDoB7k7upT1EqPYqBlqy8MUG48rV4Aokos
BxZGhEfvOBoNHzpwVLdclGPIZlINMUHlFA3xwHsOHLoYNvHV9k4MSaIPW+auQVUl
Gs/9PEXKiUJB3AtWGJ90wBABIWhvFi0By5XhSf32L1CXmFjtNUGpuK4PWPzXm539
qWbEwryujfKdC1EUqxhJ+TFoIZHzdgkG91Vc2AyN95qosl9HOp+oSdsv3pS6d6ff
B5v57uMmxLy7TA8Ln4qFS6GhaM16SJ6Wg1++ORqD3Cbps6X8Eyc5sC+gFAlegmez
0NokiitqTJ+Ih7JRzOpHMnMJAWWlmbSIkGoZw76f466NOdM6uklLjSwsrG5/j+Ub
RJ/yCLqyBkdbuuKfk6E8wb8r4Fwcs0Rg3RleLhNDdSgyfVuo5mJjZ8QKaIVLN03Z
SqNsDJs5rvaqqMkOqpr7JHLGdbuk3nnZ1QdEI9cvmrQnhkeYMhTm1rLvvk8MElfq
rQN08rjbyH3ZWodORhss3DLBPe07HtKp5RntHvfBrhGZvtRDwMcfjq+XUA533viM
rwT04YmVY/5RHUfHDLAmkgY0l00SSsEldikwbu/svM7FBmEjqSFRqd9qLHxntgm8
9xreK16lKUPmk8FmT5fDHPPTJcnRNilJCJ90O2oQyRzrQ3iZTEj011o40o6CWGW7
rKIK9rBk5J2YVy80cfJJ68YmG0qzSyL+HOgoKHlDJId91htEV/+BFunMzg87Ecgo
TXrnzbXNQ6yijQBeFmuSeNQzKrthfUqwNXkSfxAXBCrnDBcZRym/32NZn5LoLmGv
oKhfNiXX9Dwa+eSiq+1YQa2dfTRo1bPc2TjzAGckz6BLuqb0jO9uUAewERr7mw7W
mK1u+nZJlYjWIhjBCEaSETzD81TGQ5C9Q+2uwAr65mBifD7LYHBj1c4M5A70pcro
G4QOsn4FzrIcugUN8fv9kYHHLJOeLl3t95LoyTttglWEtp5bMX66QDgdqWbm4amN
kHgTEHFCAHmtfsGw1BLsSKsAXOUdiymGwlLfjqlWJKbNAg79LrTt8775xDqfSs0E
o98oJMNH1bOrEdbpp21tMPMFtiF+CDiEagOTGsRQVEDJnnTujy7jhNekeBts5DpH
e6hooeB898UzDyLlO4l/5Mk+0rVoSQQLjN2VbJi6HURfZ7uIMQ+r3vmjKq/HP8PD
4k+IqLRZbxEn9I8874HX0fDXQmsPDGBSgSsdBm6EBcZzY+JHuYdpilW6tMUVGPT2
HjoG5Ahf5X2AsxTHRSpt/1PZlwM0oLMfUSwrqfxepLYop8ua01YZKrjv7lmfwa3r
50WwS1c4yKLqAkOV9YL9UyXwTNXTlKumqac5N8mNdQRgeiWDEL+NxxAhhextVbGM
VU1+oR9b0jfg6Si3fdc0vZb8APsICLoZ5ybnFO/2aM6HGEq2xNPqZtGPKwf/Uct7
Vv/OcpBxVCuvLSUcE9G4rKQ6Q6qrpCzTEyZkGIDsz7hOfxWHpIsOvKau/V1WYnPP
huGUJHshCZA52lad4gMALMVEqdOUc9MYXPaSjK422Ox90xXUGCr7u/EpuxMLurS5
2AE1M2Z6yZeSOd1syj4bMzQfAGULYpo5DX3XHFwt25h9g6raxlfcofl+tBO1ITkX
V+jNTvB42e8h1yey1RxTrIFhNj/sC0P2Lh5v8PorgjzTNbNhd1O2k9/dL/mo+mB3
LSLw7pweM1mUgrS4QLhM7rEhEB38H7/WjWQ4D53WKc/OyjsPZjHRZXTji9Y81V2/
ufFT4il6S1JRovluSwC5VWkv/p7KZJgSqDHq344LHZiEwNDm6W2301AHDvbFAJR0
tCCRcC06QyFgcHbc7kLC9o4ZFM0VFhcwimym1uyxS5dOq668ArVHfomXZu5qjjvF
zVA2TERkB7caJSU+WyJLKJ1ChhvaEn80s5ND0M0YjmJqsDGKKwVPNjzrtxph2XHy
/Fq4RkEu978pQaA7SDUIkHWTGofBxLRZYB7v+CHP7+bcl95OLnSnufutbcKf9fMU
tNYE8gtTlx/8C3ljVkjZj9hZJoFOt50AaN5ir/uHWSIq/RCaE/OTJtVaO8Buc/Dt
Cuib2KECjG+R45zGfnrDJhqys5DslDO9YmGrqkLzvGm2Y6RyDjW7fd6Whin0R5MV
ZVZJLy6/4vESHfib44UH/0YhVlHh+59Uo2SHI/Wwg5MZELaiut1gL/kc1JvY97l+
YNFifcRMr8gsFDvxaKtY4jEiZ9vZgKc4HG4Y5PjLDHwxjV5CcyPFbAHAhQPlSSEM
chBD60+Ct8hYVhONU1O5IVa+JieHx+w0tVTzF09QIBIaxOWwu8Ex2GW1GyhoALei
3N8akC1B9XHtzXj0khpSelqq+VNup0N3D5IB3lAU889GtleqZnmgVwEdbjm5/t3j
C0dvX1YYO3OoIkizMXe9a1gPhbGmIwhDh6Y81uvFqAxA5IdTC/e0B14NzsG5qG8L
i8lGrbxzWGOTTkKVGdx3qcNC3xs23GJ9wW7oxEI891MZwQK8s/ZcobqpB0xLDgvt
WE9u3+zx0sL01BZOkEqrTgUNYxxJwc3Ae06ddg/0LStVwOgZ1zRU4AG8IDHiMqsk
gUrYIBkf+3MEZKV4e7VHS5tW0KJSfoV5guvsczxCnvsxTFtx8VNGenWTbwNrROHu
AYfGoK5ODCuLiBdapjd13KrpeGVlVs0Hs0ZNOHSWCyELa6m6Ad12+V/qHJZCLVod
JnKzmKyWUlk1/eG5X71OVNWjDDZi8WyfeETitaXHkDl7xrtNlecc+VcczWUrNP7W
s4rc5UBIYiojwNVvEh0HJKeYxeDQRkrTgQu4EV0UGLUUWizqNh0579BmDSIZCRfn
/ujCvDE/knFFarEcGlU5rL62ovYoUZELhpD/RDnA0X52MMl4cqpnekAw6bq9zEd4
aGW1uu9F6j7SBJyDqqZpRYI6aI28XRD94DMLZdws6GuIRzikHhQSG6fc9Vwh3R2A
mtrb7dOGo7eBS7/aBhr6k1Lzjo5XG/4Yh5wcbJy1agyc9w2IWaRTGEzLszO6xdX7
WQFQr7D3O08TmQqyez6AycrZbz9M/8xQ8iIiBu/iccp5ATGciBGRkNOMg1qnZYWk
4Yz5z3XaPTi8x7xeYydEa2A1Xya0ztO7bH3hpTt2gNzMZzV7Tm5JGanB0AnSMogx
qVDPhZcSLutfp+fB0+oAChRkymBHjt6ZHC5Euzz3pBpxyy8gnbYATys9SV6LZbtX
14hDzMcu39w0DPzAMZ8z9wBJCoBtMiZGKQxIhK/IKimTzWU+8L2OI6emqXfThRys
CUVYuSEk22VpYxzB8RoOJeQJcNjX4/lOoToJD8PguA3HkFpbnUuJVzjSjNM0Q7Fj
PmMDRa6/Hw4pk+xg2UtbyppZqHMpEbsa8IuwY2LsQqE5f40LCwBy155yEK8vZQJ5
jwhOw0OFbR/mVvPRy4DOgYzru4UaqIjiXBK9s8T9KN4c0NQaLO35NVvs7YXycprD
NgR19sE6kHGvjZkFPVYfLJ9GsFUisOydQjcM6062fVxY73zLv9/Wp/Z4IFvfC1ZG
7Q0GAhLKaA6sBRh2R7veIGMhGCH6yJ3beiZPgkAWQrbHqIMLUe55gpDBLejd7eGf
BBPLOOttwQw75eSFDWGcZ2NMm+y2pdOAuRdjc6J3SPw0Kc9Z9/slQuJGJU7l9XNO
qU2QVxmsLYkwgnCjRF+jyYjhzo1BDGQQ6O0+WWV6AADJxx1Q4O0i72I7wxO2YcLP
UzjIgMzu0oHiGCOl9PWvICgf6jYJsDKNSOJlkxnXXk6qbYDhgwt/kiqFkLfnAxdk
JlVUHG/v0pdDHTF4bg/pGFYuWxS3fG2Ht73faZhyt+MXQzWLY4ebjshI4PjQhIZA
zs+t1lWy0NOksj1Z6TsSERMBOeExOibdC4Dspa9rOdVSYsbU4KjNmmJ3PeLUeKWU
u3RE8psGohhaHbfr4Zd+1qaPjVW1Sckj6efqjSROyoGumHgATu1Wwk9Dnki8k8EG
TvhDOehFEKNlcJ4ELyFYutft1RD2vX+LA4gqkaSu212tHnVg7WA1Op7ic3qoBsDf
hSmgJQGD3bxs99irzhks3hcxPN4aqSEshDkvReCj3sfU0396c1B7KOLSnxwUzDjg
yUQBBIGSmJagbiRM73dB4OiPo1KN9BpLym9nlOyR1VxygeOu9ui+Tg/Bo6XK4P4m
ThATVIkDrMYkWs2Y+N+t7VRWROBztxhNG2mCuJftqNYGOeeXpoIiy2rGYZae6Jg/
PEqqYIx02JzZON9xn4xx1ZyS8pGROVDTJsLUJHd40NUz6zAASAlK0IYw2+IMak6j
fgDMD7uNchfvW0fHz3RPKlJ+Y+i6qYFZg70oxOEoutt4rXUoeNcdH3FRSx6figwI
awhAAAU2tYNGlLR/2Wus0YxczlBncm2Gfe2/IfzvHYCKMuhXGMgCaATKHAu6MAuo
Y8apbJlSLZAWrIGGdDu6ukHFC7jTPUfy3blwHB6j84wEIvB+aj/9FGdXdlOC3bJy
KA8xRDx+koFRIY1BLtKlpAxBi41K+vKd4BpSDFnPR3zrjfFgnhGbwwOdq9oaJQfK
yO5KB7pJutt+5GT5ncWPVCSVyHjyiOnR/rXWqhPd+zz0U6WfSJMStidhBC0x5Fyx
DudFZZ7Lt1ugX8Jth439DVjcrJBo9CaqmHodC8cnZvhygRUht52ISqII+AJX1Z7+
UD0se7RgiRlm+MTtco8P9blcMSh/FJSb2R8fGTYeye9gAVJfxNfSUyQBk/uRpYaa
nsxeOPDojTeQ5FMYrQeyfWpFuYrdx8LW0vd6ZYOyvYbrUJGgp8irSGrYMzgj9V92
0sD0wYxDuYkQ/6Mb2nrRVBzAI+kKOd/y+pMcJE+ufr6obnwBjwwkANrw41IBuzc3
lHoRVyPFWtHcynZLT3r/Z3OPMqr+5dvn0QBynsdGoLsznrBJMkeMPmGLS6ppyBsL
DVLYDO+x+hvsairgDtSyltw5fuI0liJA+2jHDOd1CgJpToNzObRHxVbg2luY/G06
uFIlIwiDJiFPgzJ7gVeFwsuxTSoU+vNIEkT/Vj90fEwzEVIz/1O25Jo+DA9mkZR0
IaZpuetrFfSRJiy5gjVK9FxEkQijm3hkJxDX5VHmO6CvT2fdqS72lmUxjo3z8UIr
Mcq0iEQR737ZnOSOElMc/e1VyBpjVNCrSujX0ndtZOlMMPqG/wi9Y11/ky+0J3dM
UKNkiLHMxQ/zRlGO+TcJr/ncfnQZLRNJs9FpJSxNynjZm70QHzRhSLlHnrHWOL5p
kCSgyeuNHe5L21T83pCwGIOUYNGpYXVFe/D99NL1ONwcTaPMejI6sMSMJAjIk1Td
sZ5uLVj4+iRtlBj/Y58/rQ2ubRuMwdA3ldJNir4g4FAjK8ksIIA1zMWUGb1Aj9lO
6VkWMo/NZq/lkKXqU4yhIqyshvXdjFEDM26dfrmh01zFfWamZ7XO3DOpRwCJR7o/
1+id0p/Uthu2WsuJCox9+lGlgwygh6cBlu9272nQrBheSvRKJKHqnDMItoofXHQn
xmV9GW0OUmUEBK4HYgVM8UWJ3DUcOkOSdK5MriZEwxRd18joblzTApGJA/TyChbV
z3csZhiQETpBIyOrFFSUHe7siIg3BuCff1WaljZghR15q6x3ipBgbnMLSZ/zJ1hx
VlEw94c4Z5fiNpvgqMwNwvI0AnwL7mjkPvtiMt3AQN3E6qIhXENtmIUscqcUpBiC
2YatdhrKz/StQJwwEQulgwJa/wFwGtzgrBMWmhdKB+d4SPBKeiGyNDu30Q2WeMgY
pHtkdqTfYTCPk30OX7S1i7kgA40NxE98jqMC+KSrUDxaRLPUZFMopaueHO3bUaQe
c6uCUUmzmpIIL/5RJzqe5NnGoWZ/zsgk22XAwZ1dpBxpW4RVInBRyewjq6BaG0ET
3NE5Yhnmg1A6Fm+siIGVA04bAQNN+Wnp570zHfuQCJszzj9J2crM1u2nhKA6kxxA
LdO8owc2j+NDgdoDle7tYxah62U8JeCN4yK20XTkP9lkkBVjHEHPk3bolu1fCmlj
eYaTisfZuXgu/gstEDekXUVbhrIaEIyiMCwffo3UEfRnbfG81KJdnZqkN8ZjCOXi
X8puaWPu9V/uueD96JqNn+/LiC6FERNPRq/ZQgrDqghRRriFxtsmUcPhJQtY33Vq
+XQjsV714Jqmja+FudLlORCXMBepRgUYskuIopik8dM=
`pragma protect end_protected
