// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:45:30 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sObCHO39x0KCVr01xYhDYGV/YHg+RsBwzMz9mVSMPz4Qwqjhoh4dDpM0PXIpHR0b
PDEWSQ02wOvM4+OyIl9kLglCPKXOCS7IYDHAlvWyTYw2iAYgKDyNG8xHWrxeSguN
iwC+eNWp6pmtLgyy1qG6ezCXXl8N9rL1W9xUMHcdYwQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22672)
NG7n4Bso3Zm0cI4n6n1b0h1vbDsUl1VKu4AwNQSQ4TejM8BZbUMn+QTFwG09/R2D
Jd+8of++qrKfQ9Fq0YMZsB4NfY76HA2XOYBGvz92tuYG1LKES+QmEfBjNLKP+kcI
+hUDOo+oK9lleP/x7IRWvjdl6/yohFlOM8w58t3aGma3Lrn8E1qyzdm/t4Kdvmve
N9sYOilQUFYHGilPpLkiRaDd20JkarNA/xGd038eamiLTo/dSiHXFmsWiQRVNMZv
sRkfM5h9v3BQmZJpoevyT8K6BcKu4iBsAd/KPJbF5frUVd7v9P5hZ7WfPIXQLEFT
Vwl5Py946xbk8QdJoD6b2vbhaWL8M5tBfEYeyBWKuzoDX8dbzWAXmyddlJvgzH21
2SRj+Sh3CHOnmDIureP68BIsZ91wRQPPJw/JBCxm21PfaNxPbcxUMyIhGbAfcslD
Ee9Jkn3WV4v4tFKM0XtFLgw3HfZ6Lc5TGbd1KVkxtDkmnXIZ9yic/YDigQuj6crf
cE8ZvzPdJ+R3iYmiHwlFqtmBQjyZLBh574inHEDnzg2IkJATI6Xpgnf2vPmaVe+P
uhuvebazAEGAmvWBcbUhpjPCcbBZAd/gl9889l38hDjtarJ4B2g573DjSXSopqz4
1YPvkOzTq3ZQqnsWdEO4T5JCRTba7VO1b3potdjYAad5TuzlzzlFXmwJlWu87TIc
WZlnEIvZ7kMR09aWRfPpM+C+U5rdtgWfjXQ+CC0dXDZpoorrmKY8Hh1cKppJ7dVc
YWFOvCgy/6uDtCeY+ujMKYrP6N2jHHU3eVQRgh07R0CUunyZrrx/YPXHwF1UcAPW
OSBx8aM6V49DmQkqsug6B87MlK808y+YBln6O4kUHAENMVHky3FQ9upi6mOOG5fZ
l5R6fwHgUawCYtCv6e2fnPRkiujTk7CHrl2wmiFbP43+gESq5qXuVUViNht6VHbg
2AdSMOnglxXsi13F84y8ytVWa4JM7CerpQU9Zuo2/WnSWTpu6cWw94uzz7ONGkTJ
ScIzOk1zCS3DKvhHQ2RuxmaW2ru8VB234g4GXYAWGwbinwwqFHjWBh2SqDKGrG1p
jG4l6WPyyhhnynjIXFnZSJxkX+zG9Bl4M6mt30LBZ0DGG95q7Ahn0H3Xkuwi+55h
nINlMiVKCxjVzrQsbQoAzEjfdOk19cUs5qEbzSwMIvif29iiLFVkjxNS+jm8DA08
BLzIc9WgF+D7FYcQqECFiWAPRABJRDqxGrfoHmEo1jmF0jpK5NEGD7AeH6dwFZ9O
e+0LLT9pJAmFt1aj6ohM9UHBQnbG2/YztUlz9bPYnkKJ1zfwpeYeUJa0xINWbeoZ
bI8gY9F27SOqXj2tsj3GaSj6YOxv69Cf08j8fRSepRiGylc0DKJwcxJPQr2RoOXe
l1LSNm7JyrhtS8kHX29DWRxNZ/7x6IlWYis1wLjRXV67mFs7H15G8x6y10X11Xxz
ZDuN+fcluWEcqY74Tn+fzORjesmhz5FHNbtxHlqcKRK1Iorclq6HTU/DZ8EtIYEG
tRY7k6w0AVxt5gU+1u8g692nl+vVwLpabejBjNAF4rLj/JdVlBjmb8P4WDwRIaOu
xe+vcggrPnD7dZRfv4/XsN/3zP9zAiR5MKfVlYvq82EOKU5jVBWcsBUnP+CY3grj
hy6KZicDFtTwTMF6BClSEltGFXjNDtbljhBnS8rJTrxUkfXwOznPgShcOpCTWjFo
YuMV9XsmUtS1s1urbOAg8WbFriWojXmqRuJ5mmA5UY7AhmSEPVukXNrRESQnBIwh
Iezz5mMcaHUfxCjn+pcgyFDLOwZuaNBvZKhuBSGTgNjdi/f5W93M/qWcVbNonB6G
FpnZ91lOgzlqOyVrEIZ1PNSRHST7vdJzAekE3WSDN7cAfzCy36saNujbnCI55cCz
lx0w8CpFlx9EuBaOM1iQWnwQS1FpZ2mqEZCH88ua8R+fHX9ELfUxBRz02Bsnrn2v
lDVlvR3v3ssJeXkGHcRzCyFLUO4FGXbbSW0gJK2w1dOXuM6/+XWGE4ODIwRcgRBQ
ETttMUJhAHRCZ29Pb8ZYBZVXsbsGSZc7GHwOah5Dq817ryIOE+IphMNfAk8Cmk7F
0KZetkZDy5hjeUh65xMJnnjI86GmV8XPlYujE7bt/+3yOD23uy/kqQU/RgiL18Yd
DJm0OLGfczMduZK1hx/AIKgIax06G4JM45vUpKsMqfCpsH13wOQbCnTifCsiiaZ7
vcXY4TOijZGmDwQgzooFaGhWOg0xqd7ZvO0zOkbwRBn9lSwuHYwOMlP/FNsFyE+Y
NKavAash8hHK8iAy+JysuSb+E9+lK5fRlX86gr1AbWJnvEYZ2v8MXr+soafoMdmC
GP9hMlTa2/oisGxEQyb8kdonbWS2y0LjtqFJyoCPnwFO50V9C0RS7OV9ToJFO72F
gQhjF7F7po1M/Jh2MN5pROtVlBmfLPFPgC85LHn+KMW10cxwTHGNYXwMjxMX5l7a
7yLRP+bZRBJgEYmrLuo9cqq5cYcUxG5aEaKcy0o14+TK8p/ujXXjQ+DJqYCQFlbD
Lz3Nvg/uPjBwlyNZzYyGJ98If9v3v1eRKix31PQWoMXaHUqCrMGIl2R4SDZmMP30
FlBXCArorunwjDICcfEauGF53xlgoE/jWXV0T5sYpOeJrC6URvUDeOslk1KIbte7
A9SKDrdBw8bZdHiqq0QVZ59xU66/J+sdZo46tLQ5cD172+89vc2zYcmHku7F/3T1
i0v5uNaQXYOdwMpAQvuFrdUk+pLlSJFm9uJgU6THVNJ2DkEYrXo0n7xne3W28upz
m0mW9kuufPdnU0yu7WBKc0VOASh46bvsVb/2QRwtoDKDpAV4Zr+RyYomLPphsKq+
9nzyb8oXHtlueJUgQ8h+uX9Mq0rJdUj8MjFUNtdPVzolsRW/qkMGYLgv4sREa5fk
sxXmcrVcE/J9+/WUTZdI6p8G3cHF2kwKWQe4SsJR8mZhHThIo93BE88b4LAPuFpd
9Hq3OP7tJ2iiDFBgWd+89fP+WyaqZlvvxhL705fn8oVRunmAd6bDtaCTBKvgwBmb
TX9oPts72nn0iAaUC7/k+yPcpO502nQEUiZJ7x6X4dSKtpRZfi6pkUtGY1JZFkGK
Opaef5D4tyvu2PRN4493KIcpNcJS+Z7EukGVu0cbDAncTu0dCsBiP+AewYVn6ALl
5FPyS8qQ3qzsrbiq+/33ehe7/+pO4tw+S+M/ovj3bqOs9yurmJfBN1Ij3eXPr4Qs
YXLqcwyf3Twl90nue2sQ2JCQEU3qxRBIUnCCV0vXTDvXBcxQsM4j3krJ2YmqfCN+
6PBWO9NJ9XtqcI83YmzZAnhtU6hr1r5pNLdTaf0Rt/PLqQoODCVBd+/nc0tKF3PS
X6zzC+4lbw3Sg9RZUipJ7M/SOOR4w6nLOFLPi0YZ/qcJe8a/uKG2S5yKQCJca+LA
5N82TQ3ZsqE1q5zmq1SZPnp/Tsbshw+xGh8Y3lh/rTC+S8An6jIiB8jq4oyBDXyf
Y8obOwgyTi4eIkMjYMabu+6uN/1COy/6O3DyaHdc4dZkjiIfq5p1eY3SqEVPUo48
UTGVlWopLQZHnGsPExudvbelZjlS+FQgq4pF0LwRPruzU8X6plBxdL6AiW0De44Z
koseGSR3p+POhFieRwaVCykH1w35lK2ZSYIhx9SF3Axz+qv0MWEr61+Y6rqx3IDO
XaotDPZ6vtSYBnuUICvV3gDi1u0CJJGP4mgi7Q276Cuqs/4OHuEGS0YZckgFVNUg
irTwVOEt4zsyh5WEkItQOF9Jd9gn359gxwatayycf8+g0zZqqYbYRGHdlLEDovWa
opwfzipbnceuc0j37ul1kEdSzrCDhKA7CxgrElJdK8fFKvQ7kjYSGOHkVb9kw2Sa
Fo0UWJx8VgAjP3RVzn14idlUOVu0HBjTwZ/F3HR0FrftErCBqTpicCVCvZjMjEXV
5a4jbkEN+dKBkfU5RxzuLNLzizAXNyW/Fd35avQIi8ojL+Le/Mz7cmAM/yiOnTAU
0G+fEa6r4BsTzg57SpuDXHZHRmdHenPR5JwoDVmCZgFyPM5n/kYt86Y6jVMjZIjT
qjIch1w8hQneqU2YKbLIIxplFiAy/5iDGcNfXq6Ci2nW4itnos1HKyatwNCEx+GP
G+1Z4Kdf7ccStRMr4328iARMQCVgeaSNYUlVpl9wZsQqPZnIbAeobvqr+xVLc3Gu
ZIAiPMxfiS1++/kypoa9yUmJ1eK/Ck8uuw5oQp3rjZ+V6euTQPpx4lf4LLSdiJeR
SBAc6xajvpj3p8Sgn5B5FZ2eRwZ/NlP9l1N1aVQf8w58M6DC38xF/mdlc4bJNIuY
ZjDx285NSEcXaxcy/3JdRwC+zxWtflxFlabIohK0fJ/6LDUSmFugOKDylDVaADgu
xAoS9Jo5vdrPiCGwbqkSb5k6BKgfTEL1dG51O2a9CLsZT3p67mq0AeDPb9ityeJ6
rAMbn+N97n/x5Ycl7bitvpFVJF4YCxmjqW/FoKywDKhCfUt7d2qWFs21yTgxQEa7
bMMKCDajoMPGfZvT9SHMioivaWErEKjWJyP6coy7bhhCGKw+V4/lXJqVBxe0+sPP
lb7Zi9jXrsdRGLA2s64GGvoZwrNB0LMGWFT+cECTEtUt23s93mKmBn4EERs1Nm9u
Hy49w96M27Uud/+Gd+gh/eOSlIAfe99PrC4Tm5zAwgHiVxcDYOgptdJ1fg7akeHw
Oqn1/fLWj6UH8y9hN2qKL+ZNogPI33H9NYTM9R30B7iHjPZVpie2G+gPC1PmeIU9
bFEqUOgW3siu6Bofweg8Gs1gKxGqd1WN8KJbP5aR9VxALFFG8tYgr+DDMlTdNvCK
k/mvfR8g/BgKhRzI0XoGxMKp1qzTwNBcmeY11y7o1k/YUXMdu2jM6+TkEnqbo9jz
9Imj7smh2x7OMVNSnhE0Qf37TwCzp8YQXzDEPwRz8lVv1Qlxn3bK9xhw+0s2uPlD
gqoPN9+3b9r1eNxOmPvVLrKLaQxb/Opg+0Kr9h1DuZvcABMZqgNveirAhlcM2Wcq
ceQKmwd3W5TiiyKws7VMaEjjcMoXoUw/LfH3mmZxZeqa/yUZE8mQBjz9T5OdnNMZ
qDcc/DIh2ytcHBLSTBFxaUSU7RiEY1C6r/u6zVYWNz5/oHeznHV2yP9m+Na47VPi
r4ZeeSVdgke4WtHYVPQENyhcLhB9Ke8BTJY5WwsbhhJcK/9MfjMzlvc/VMXB1VgG
cA5x7Yt4Oz/LG1oQBQbXy/gPkEBxcZkWu2ajaZSn460NTCAzLmxqbfvsUSIooZmf
96z9AriYD4+pBe79LIkCG69CQ4gOOeKzY8VV8t5VXDTSCQ95KiAPDnINHxB5j5s3
tqQSR0kJoa2e9zUi21fizDnOZoyAawVwyKT289OV61RPdCE1mE0yg1mTMPz8ueh1
rmwfjwyUakcWgdSVl4oYr6xNFVcbtRFn8DsHdIWIkJ1x5aPmWO9REHHIqbVi9vXv
Ots4Bdk5BVgzPgiNu7YAKr99o+nX7DZ2RMGyaUrRq7lh1Tc4ToOvKKEZq1QM99A3
rzUf1lXfdEKtzUeFpmTZNzf0NOvG1PVa8syXIGO6zn6fI1gcb0uXJa+QQooWiNbu
1ZNGKztbZNc9odJjUsM+98s2cngfc0huDPkhOqC6wACZDJ5E1jqyxvDMTr05GAAP
dSTqdXbd9ib5Au0hRije5t40y0MB0QAuP2YQegUCriozpfd34o5ZjWBjwRM+RnJo
/oEI1DOdG3xwAlq2KUvlLvhoIzAdQr+3QZ2QJDjy2lQ+rJGMV97B7YnSBOXITjZD
3Bz/BbQ3uKV31566OMMb0a39y0JiLhOMzJARpdAqrnjmqHj6n0zGTV2ZxR5Qaj9e
EgcL5hjC1XXf9i26Mmtpqf0qP5bl3Boc4Dn0xDyfS2YAALhudZ7+bPJRchRyYuUE
TAwxvKecB+mJTSzJ/Cdu6bDrSr3t4PJViZ/xZQK7BqYESwmREHTD/rZ4JPIKBaD5
qAddaFCWcRebBoqVDN3rn732u1GcSby/SgnUk/DHoPE7acaFLRo4J4ucKPS+2bsZ
B20GiDN/M/knSjjWQoOyoMc6P7H7DMycqbOYgipFBQ/J8X1Ya2Thm5c3GggTBGFY
WVTqbArbAqRh8UDuSyP9ngpqcZZ4sLygiMFQoSBhNAl+tMmQptvivUo3B36L48ZZ
/R2xXYzjxPyuyBA8mMkXLVzMadcrTTHIyDJiQacAH5JgMnpz1Tm+s/g++3CzClXs
KJ9ft5cGVNgoYn1xC/JhlTCSyuIGGyKWAlKoHSqCVwGU0r7fyfz3hv5yggV6GZo7
ghQIrT9QJivfTbPu/WxnPc5i7piHT2sJsQQUqEgoUypD5EPep3VO0/G76SwGrnC4
hz6vTH0I+/o1Qmv4dze9qmiWGhbwbRimfP00xwOKsoXLLpsBj9bJSkOQLZJF8BHJ
ycpKJ39aZCW+KxgJcBsEFYnoJ3y4MZ0wyn4jdM/iQZE6pw1XkOBZFVYtjDhBmFSk
o0C9rO2vnKY0ktkkYaPA3/Y3ARSp0tr2aYWJxy9hjm44H0dlag8j97z0Cdw/7z/z
75x+J0k0FL0SBR0zEaIBIsvDlTa3CSwO8jbyyIaAnKWLwtCZxTn6WW4y0vMlOtzW
YEbz1TU1RsJ/GOwOC2pj9FaYKAcCEU0Kz6kDrpu1BqTmBm33kS2l4a9NMuNxyqij
6s/t6zYI6Xvt91MrssoeeoAbbtJXWAT4utA5ho3P9jX2gDm3hucL8fl7Czey2k+w
Jt8Z+ZDAiQdgG2sI6pOrRcUdu5UoI5KXLijwZLIy8HqbElvGmwJmTH/8ZFQ9WOm7
tlrraamGBW2kKnYNWEn1bIcydtYtc0TJfkOP/MrfTkoA6dQpg6S+PJ4ZJuji7aAz
GvyPv6V22oWUlufJRUbqRKks3hXyyWAoHLq6jnojuScWny/6LU+v15WgRpp8usmn
bpKevVqACUF48eUn7SCVYIAMTge9axqGR5Ff7iud+v1P22d59LXP4b67826a5Muh
nx4RnZHlmSxBhOvzRCWJVHX7r2p78CZu/kzFfd048rRORN/z5g+Fh1OmFDBxayE/
oCQxEkzmm49yiokTKUwfIAyVR74uGHA+J0ykqbNETqSfABG7zNfdSJKBjfVQEebm
ulqjGk1soYj20Ok+VywuBi6Bw4LNfSLTNgMOhnckn8o+ON6R0XhlGUPL2K7qfpWk
NJ72H2x2wDUFE+zWWxBOZwMFO1Em+8TpyffcuiiJm40g2fFFG7a2Nyb2FWkXmuPV
4oxRZ3yp+6mGI8SU1C8jczF44HaOVw4Opz94/PoCiukEbNLZIxB3hPaihxaHWZBp
ji9nyUseh1LI2kxv8DUorAQANF8fT/hOW2jPfaeFjh6LzT1EEcU6atBFpFqjHv24
glIKuZNnrdNo2SLpPENckilgwiuHpk5ftZu+wVc6T2lDPiwPrm/zwhuWZW620Ye/
orfQjLW1+hn2CmT//tAWqNezmEN8Z7KOqQyVJsA+UynDTF2loPM5JtJXcElb+ETu
I8RYRjG+Mnj6aNCO3PCBab+pJA3AkNxIy2p0GdTb6Bo1Jc3bLW9nZFR8HG0+qM6Y
ldFN4pbjJH8dsAE9TtLIMoc5mCPGb0urdZhY9eEQzYPNyZVH2gle+j671zkShuWN
gT9ybetPdnxMWaB3fe6swboJ44RNIJpe51Q8zbYI/235qelmi41RZ0REiyrF+M0L
hAN5hAawGP89G2Ly5PrdBiiLU3/2yES2mMrXw6QecAtOG/K2Ugnw6RXLHgdNP0jG
l86+yTx/CYjJIHjlE2sbv8osrfh2dv2GottwyPJwDuc2jAuLxIjIG64zxynthPQA
bxVDRHnRrVSScHlSa9B5GmGIUfqi1t3Y8sSwhMigRl1vnv1ygeaIsierTIbGtCs4
sYKYqUN2wyIt+DrY0vTP1ndDwom3BlXVuFlyPB/B1ZG8svTcOAtgF4q3/vYTVfSv
6NPY8HYRDri8LSxADqs1uW/ULyWhWC7lG8hHKTIGW9QzmOF1AOwBaCfmy7xagOLs
5TUwDL4Z+YSCYLWpMvnK+rBgf3m1Fvg5oigVyJaNZwNGM3FJvTpOz8Fp9jxIfCyY
RAUHRZQh63cF6UrRqMi8NTjlgftzcWlBG/dL8gNtOTqN13N9wS72SMCew1cG1ly+
m2YPDcIQPSLeRm63hgdkiCAzbgwFKeZoRaNJ9cuxxTVvykgNRaj7ipnxWAMTP6ua
rfVLvq/UfGGZUsowrcikgkRiiJAPIpFb2tOwVch3u6a9T1UlmeNQ6mtFzsbn6mn2
xTfKbGmDXfEFpoJJhb6u1b5Co/RxQRR7KK2jaZzSWlA9Z9P0JScNbsXnL3HGn9Jv
CyTl6lPJ7FtBLDgY+AD282Rqb6jivIEBzxb+lEfKco3Fqiw3EuETzbMIqr7mDJZN
z99E4ihxn0k60Sn+aprPSsu/iY5F2CieC0O/YdUwmkYJiP4yBNuUZuXktkwfQjYC
ddKwdwXSjo62FP0MnarfPagDhOZeYDHTv3jAtZ135u7zv1uvpd/JrNEjif+qQf2y
vk3W1ZkV6sGIAW8d/Q2ChtkEv4MuGcB8GzA1TLVjNwlXBWiygBwdQqSv1X5YaxR1
zdsw8CF0u3sphHO4bBoFRnDsRscUqyCcX3KFS8s4vBfkdwBzlyaPtG9sycOxIzDB
iArAAbwGlODy3SdTmASBMeSgYMqlaYA891fKj8AWmU1+gmd9hYc7beJLlFdJ/vpr
Ht6I2PBuvHS5w0E3E120BVjke1OCV63DFuJiBj2H1dbTVJxaFwsnS+r9Rplrid8k
TXy3d3YSl/msubsQyGxm3wu8jGCJA9i/uhNngrGSHdGj1ijtjCr7WeS3ufcwxNuh
7RPHC4a30pbsj/x/MYwUUfno++HSRR1o/uSSgUiqdyVxzSMSJujeeG31Bd/o3gOO
jkO7xL5LSPOLfMh24B7HHJrASoG/Sir7IuNU4mTQoVoOi/JpZbM9QduyZTDAgkqh
dto2/1VDfoqOsuP6UWZt7/QyAkm3LVycDy1/+A3OFz+NWeSgwUH3WKhbXAeFWGk8
SKacnwojtQoYuWEyfW6L34IiUWFLePUoEI6z9xvZrBJ25i6VK0veN9NJIfduPbed
XNIKpo7kNJ53qIju6GTKxypXKR/CUWcQzFjr0b0wKbNETEuQtHgiOQJ1DQX/zBzt
M/KxKbPOlJY05rpvliqvAK6DQgsKqaTZyEQUm9dQGCpzRfB467S2RHS76iNGJ2xA
OcW/Ub/5lFsfbCZxhFA26s5kGDfL7TMLft8Q7R0CcJPLIYVjLrmbdS3rlUC/UMrQ
3GYDuXK/rqJ/lbTFbwpxmDqAXF8/loOoIhpG/hhdd6A0OnihiSNeJm03cusRrI4/
dP8d7f4TfcBBzCbF2TCY+J+tv4HYoGiv73KuuEpVV5Q8+jznR9xbEg0fK5oepet5
Ip0fQCoGTvRFZuuFLrLDNtaOqe6X4YXAczPJvrpNaJdQT43cBNIlBE5lEyM34k1x
MO7WBHEWa+Ry3oBOfnpW0cT0pkqSx5arCYf574hhOtBv1mLrnhQtBhGlxgrpR+Rv
Bloyiudz65VN8oMaltPw8f/IPyGZq2hfT764myn3y5w8X+2oqeb5KwBCrqp0e1EQ
Sh3UpM8noRV3WVX3F31/T//GV63CBRCx9z6OpGg9AQKb7I5vzaZTt5aVUaBP9U6o
L0cEJr+YJMaum81JosiGuhAH/nuc1t1C4kbzuJ6E+6SgE512xGXPJmbktR+OHeTs
4LEIUh5XznYn9xCODcXFNdSpEdgBz93JtAZDfPSNby0/Z7c+WoVFr+0KH5rApgVc
Q/DMkxGlc/wmzlHgP2eZJj55mR3sKfohFCXXzosDb1QZ8jtLmDJD9NxGPg15SdGc
IM41IKVTF9NOLN9MkQiJYcKngdbbVxfvcQpX5oogqymLCCmcRQDkr24kxm/5q4Ah
1DGzQWYN9yp7F7C4ELcncSrGl3Zd64sUxDHrr00AioI84xPUO52a/zL0vs4pmymT
YBX37w32uIXiyp/rUE6lQPdBug9Ig0ThRVKSCdaUuak1jDCmnsPV/wWOugjDVaW9
03+0sULDSqTfvCZ7tyWRwR4BMIUjoDba3hkEb7yRC50WXm2FSWIoCZUTvN6wFwqf
7wT/aeBCiAzwoN37szVr1hzd5JVzYw68g3SHXorKlAcRuiAxfCq10xzN01VKPfhj
x6xsBvc3k6yJOXh7Fb4Mxe+tCfV1N3k0exqu9QXXgDA2rcedjtzLdE0q92yhW010
5d6EPXNQXAUKTS/RGDgccIfISKeAFL+KXsZ0eaMQYZYRo0x/RdNrlG/5hbMbjNGf
AUeaPoy69P19YnGMTqe9Sl/TvX+Nr0PAy2MR7eB9meBY7bn1m4ZJXLb7NQlf+rPz
dBwje3V9ypN2AOB3SF40OcVIaL83g0CGlA9y/WXBYsWcHWK88uvFPYULvzOjes6o
3C4+FhKnePTOxn6xoVN4L9S+W2SAHm50kvUxihEMbXzt88pErSLQCFmunrMsb0hc
cfwJwHQqURXi1Ye0RbxLQ1qN1fhWoVlfb0Kl0sVnDEsAP7jCYmNzRgjFxDhKnKNU
gmGFiH5lh4bJ7m0og09Hzc3WcCu5rNjdwR94fXrS4XMeWsR5lHfUo8CxrUnn4IH5
sb0arDw4cQavxwGBNmRQFRGK5igi0uOSx9Ts/rJP8bdBIA6id0EHXACxK8g2Y0xW
3xAIeWhpfCxNlarSvKvLWvXe/ZL0M9S18kkbWCQjot03a5Gugwdau7CoiBbFyTPU
8K2/HJbi9taQskkRmAyvWOwuYIrVdXlD1EyUqFroddcb+xHhIKQp5+AnpbJZhQYp
tkPOBPYKnfsWstrSeg7hDrFD9GynTzQu4FFM5nojJ5SzfqTiSC+aY6ZOrbmn5bnb
cfYqVPJ22MSKJB8qu5/3bhO4e6RupwHecHPXxOq0g2IFhILgSD47vUuSH4+fnBIH
nMJ/mTX8R84mNTkac8rxJw/w1FFyHczWxjPmCWqb3rST1uaOVQj/FlHvl00C9eDN
xYTq1OD7AWyocv309arr/ei/ocp+FQ0oBPYbcBLTkiNYDI8s0q5xFEBlYGorwzfC
uRSpOu25PyYSaRPmMiYQqhxhaZC4CfrJ8PbtimpY8krmeJiSq6CmNbB38+3f28AE
uC7YvbNMifplTKB+WEWeFI2PChJkuXebR8NPpcCTA4rxM6eXcmOwUI8dgNXRrdLh
O8sGY2DPh+kN4VShINEoPd2ZRQzYuoM94ei9sS4BZUjUWgMr6zONwi5DoMIQbab3
SDihBxs+diVJeV9dqLYDhEYYP/mlbZCX5QgU708lFVXWy+Lv796LesAQwoRXsuPU
qmpZcujrT6+B5QLoOa6xqxECaui5wQhK6jLgLadbsHc9npUist8AFqBea8tWrNCh
b4i8afNmDZHPlgqHUJ+5EQ7pZIqB3xk+6tg0jYdmOxJM+SEVH8N4roxyugTvPLsE
i3Pdjpco9RQV9N65ZpqrHvlMfcyJEHEpvcLg/QqAASlfn03PeQRicTbOp4w10snR
60Y/JUSFyo81woI5DVFpJsDel11rTcctejAXRWk7XQ8A+7NSZJWrTyko319kUS8e
+G+cjg0emU6ncZTq5TEpYNRMA25OuJQXTScmXalZ2gBqvX5B/1WE+Y0BFWQ/a66M
rwyCCeeVfQTUjYAwGca/yx7BqP5nvLWAIsf7GjryuxCr2nMUwGXbIGtWk5K2laZX
YM0FNApdUQH/kMJMvqEahySTnwX0H5VHT+QeduWtO2nDXJ6e4Y3celJCIDle59i9
n1MwlXXGgSZBlmzsmNL4rYO+f1YOwBtc/pZlw/uVyIh53dc0fG3ep+pI3dTY1uwj
HsaNPFo3G1N3OO5MFeEtR+Q/ELuqzC4byrcCYslMBKmuNvSfXsDHUfnvUBJIyGZu
fI5P1+4yvElh6pn2iNvYKu/B71qpR5AKBhxyrIXuoHnH5DGNBQRJIppnMVqmL6OA
b1R/9LBzGpEGYxt4BdVNyd/9iWkpIpZm54Z4eysUnbOIi0YnT+CfAJLy4jFCSGtR
OGCuNn5w+BcR6WvNjrnIPHaVNPXqly70rDzsVgk5lWUkq6b3/3MTvH5kKADavkpk
3ajjQOAOXvwYUcU78JDus5hgjlriTGYianvOcZ1kaqYsdri8ATCfdeNlEgz+DmwV
/Ji7744s4BpCy2ENttBMnt/FzqRwDLyoqxf1PzzNn8FB5uFlTz+eRMzyw9AW3Dez
Ixx0p0DacyGJ7QIPWLtQUsDHEEykiiFDj3rWlvBXvHNPWwLyJ2Jjbp34MBC4hMLp
LmK2OeNcFeqwaMPBb/3UrdfCkJCOdfy1a9vzyKiZgfOZKBAOgBoU0UZlTxg/OXQt
1j0VlWC/4SG1DH67OAn/I9P0AjQOeFVPKW7Vk3QUqpIIxHZKkQ5KUcXnaI/DbBVk
3d0wjziHSeI6A3Og9wVswfl4lBWEw1JoRyxuA+GUPoKxBaWsu8kLiU1Tc8xI0l72
QdUc9Nov00jiaL4LcD2D5+Vzcucf9cwRU6iiW0FuW58BjGFdnzaQn0H3qPFg3sSy
hC8ht5GDQhi2fByVOcdHaXFVgMj/VqISKqyHXiZAOFTEqqY9SbvQbtWP7J4G+ttC
XGWxbetS65MOqCaKtF2OqVoVw+OXhWtmJfvNdWT8zisGEJ2AqZEV1vL3l0uYu2w/
CdAi3hNfcmeHCYgYYi13GsUDkfShQjkALuX2MB9ExylWiMhL5CP5TQDbx+0H0jmS
08U/Iew74sz7J1LMqttx3YV3GviUlGkiMupt9bBGHzNJ0XPNtCUPDd7THg+KAQT5
Dw3PQFF5TcCxFpTa7uluW2a7ra5E5l2/0yqiXhndQNevvQ+LxDOcQ0rRp8FgFWo7
dJtlBjLqp8WwnBj0THAOImf7blVjs/+ITEdao0+dK16RBrmJisxt0P+n3qha6dtK
O8356N2+GBxrujOmwUPRR42lv5oNX6A2dQy/keOYD80klQDMVuI1Q8N6SGuaqo2t
i3DgV7RJgs5YY4JUboLk6UAPGqCtf/9OBNlEbxDCRR28DJArtg/BxRb48vxV8H7v
GEex1kbZSy64Pf3hHH3XE1lATgIMcoACDpTM32VH1PWpLcDi//zICB5huRE9QL89
m5olBOZbbZyRQgBC1PybBCgki2XkQfBEceFEqUWYuc1LxoB3UWTYbfIPSWgdp+hq
K85MnuRA+EGGr+U4izTkb0+RID3wKMgieDPm3ENXSIybMhud1Wyrz2YWufbB7MjU
h11ebem4w5vfUGis5ncstansSJRq7LCnRT8+Xs+TH7TtpliM4/gOCPjo/AeLW/jW
a1Vt3FwYuDu/O3hShGuBWtaCpA5xm8LIz55ohsCJNbUy1S8wK8lNg/TCQOwEpswu
geg87Zl5I53YEx+SA3vfpYKmKaXrhAZnngypd4mmZPhU00irh3jGijjTRwDFhboo
jfYIDUWnLq85ALj2z9zYtcLmOesEfYYL7Po/aAS/SG3gkrBd7ZOAENKBZYjAYwnp
BcJ6KeiG4L4pedfp09CmDlz+JQtjjJnla4nNLC/KSLMsLYwNj1mX156qW5ovlPiV
J385jeoxkgYriDRMWpHyckkLj9tKhqGN1gjcxcyupQTC9gMH2gluXx+HeVOPBNBK
fu7D1HLc9KmS6cWwXc2etxXNAkMp+7teeu9w+Z9UqGg6ipX6l46JLLnoJLOv7ZcR
GZdqUbM/Gv5djQOswHuxs85hh9otOSUF7JdMHOtCD6gzuzQf2NUR4VMMndRVYzlm
dXBtmLwH00kiijt5dKx+uAVDrntzZRlHneAWTZCqRq6/+Ct73WwqHKXwsqSHrRgD
DuT3aHVW87a8a1YDvXtih2sW7uKGr4bQ3vQtcwVzMiiB0vDA6HZzYMTDLtHw32Iy
1349BDJxNcU+/H0Ve1TpWAugEOhXryGCkaPrgwPSV4MgcjhSvys1t2SebyKvRPzN
1lAvxFrrV14dK+2TqG7cLRlza23IuQJrDefxypb1fkiH7PouW5t8/qZWhaS6NGmL
BEBuHiJspxANUc5HRY+Y0cYWHNSbRNt2whk0RHegvX2IwVs1DkSmRzANtypek+MJ
lYKFQSlseBY4uESgqQLjlaXiQ+oZWRGOgkDmV3atqDcIDy2dybzIlmJHaTxwXZGR
7IJfW2x22OpV5KDthThut14l/QtqnfR5Eo4D2mQ3pAmRkschGywN1G/A8SYkWTh6
IJTL6gUWlEvwzY1UMfEiYaKh0WjkzDHiHD6ha2F4HnLGhhfwfO4UPzyNUjWf5Pip
7TF+1q1DSy3N9hnRRuSKX+p+kY8fhwjn9ypgPT2OjtSsaGdN/DM4trn2SvIvhybj
wlqZtq/GeQjTEXwK5XGPHhNqCGeAOYA2Q+fJcSA+2zuqW4nasSrRUdfyiYe4xSon
zLPMgHFdTVDZLpp/OnJsi36i57XxezTirvNEo5v9+XGVebE3KqYmnbJNPxRHOOUp
r0jWM8XVJEhURhgyMDmKv2F+nAQrJeja00qo46Rd2CyI2gyUIm7jIYRXUnbBAFpf
srpCP1xorGswLM8QkmTgCssocXl7J4VXitXjdgsEg7W29IaZsjvcKJIaXA21fud4
Wq3rCeZQJAbvyV8Vwv5oMtqIGT2oLC3uILU+06S/kxtPnjwyDXKM9W56TOTUTNMo
wH/lsfeZZWKetA8EcPJRH2bE5TIgjOs+tFUdMJlpNWoW3F+GyoQYSxLaz+7o/WXH
4VtkU8QfaTGMxBzuw/WfbNveL8BsgPRJgdcHkFl7Gi5gapNF+o/bWV2wK0wo4j4d
iQ+OiNGbdSHYDM0l2MveCdOzvA5//ULFLxAP35sdq4q8cx8TmVBZM1QQm/1MgM2G
VZsfadRmTGW3Y1U9PakteGaLIFt7Vra/CdiPNS+6+gtN5roo/WSJH+xfAKnSvZhJ
oZSh4RO9DzJ6goTuu24kt17sX84KJyXmczBwSvYSvRV8J8C8/tTdnE4ufU3YoPLH
D5uRXnhb2+j7yHApRqCM1iGXums5vSrILCRpRHF4LJCoXYbiWMsmGG6hSKcXpT6R
5fJxiE3Q1/5CZFaNrHF4PqUr659aK48skcwlmR96e3wTuaVE+/ngGqEKYGiePPqT
8Q8KonQv93Odk+lxJtH6IFwtWtZKZ4dUqsjpzO6Q/iwAjl5rXG15zwd2TJGiHOk6
cKJrWrtYy8HP9+zcuQkoc5o9wyio+hbvOcbtMGGZvC4fUVx0Chxh2EpvbMg0vtwb
d/0tS4wYRI6BYI+F6iKuN6piyZBXPyVf/CcWsZ1uvcg/oS2Ud/uDR9bPIDQ/eY3G
I5Y5H0NEAzH8fUcYAwong/ASvjksVlk+YxeM9mbQCMkpQ1lEHMII/l2ySSuTtMtc
gnpkcc4I3Y4hW+PI/KFNrJ2elMyBdJSdXdpggUGhoP14Cf6ClN7HqivMe488mpw7
SUXj2r/wHJbYc5SccghqPjOOvIfr6G4N5fGOJwlV2gHDvrYoR94QAyErvBINu3cl
zrvYbAiqaqbwQY1ar+YRNIEz50vDLuN6JelBywFLApBZMMpaAAqZBkCbrrq43qlS
xuxrnyC9b1JooNjrLmS+0+TAMF3qYjST/a2cMGJNzC1Je//DEUjH5+jyhm9ZZ+WH
N3W93D4IXelLNlo3zZQPx1/57k92MfB8FA4rXTL0UvUJGhPTFgRMR73HK0DIiBqB
dSw6cP7yigEkMNsALKndD60F9OS9ejUPS79WSKc4jMaA9xMfx94rm4kvkoBJOKlC
pHZG3W0Kltq9m1G6t9EY2wQqgOWcU0+UowyKyMbW4ZZvtR7l49oI0tp3WSryF+sK
mo8Dd4R9KG1sT+xjlVGqj22Ag/xra4jTIUSbWrhsRFOCud6Fn1WGS9fTVbVmEvbQ
CqXKXMX5IOf7hbD1ZsupTT34ALhWsmaSv3GEx7VuPJzuqr5I8+Tni2PHocFF40BQ
XJowdsOLeI8ziiYwNoI6GP7olbiTgQO3zkpE0vEHjVOuqil/tb0+DKFc2/ZceqYZ
sFYb8sJpTpIzUrV+TlI5EAjc4zvz8nu5Mug/ypWcSeCxagIe54vhlvjKaImKoW3j
rAQXZaNepNZoYaY5xagbFBhuYhGjgjQXzMyN5poJde9y9jV65ejmgF1vWu5ETIfa
DZs5OjeeTwCiFV73Jp4GWoMTUdiiMEwf0YOS/GHNuFf37oR+WbsZIdpRRYrbsa5Z
6fnjw3ZBJffU2h1tpP218UYFgc6GPyUYBVMt2ffKOt2xubi8fYfLIqk5FE76yRvk
RerEfUB8fAU/TC1GUclVbQWXegfg6FmYDNfpnc2SC7qDpd4a1BIecTlYpydoqGrQ
BYcDSJFdMg6iMKDtL6GXtAsZ7e/Z5KmsVmZ3wJpAHyTcsecAAmTTDdZk7WMo4st3
BqcP8t/DNGfbvfzT1ElHT8uynDVjSjHIKLnQvWrs/NTpxFuJxg0W+qvLfTcKaURX
TQu19Upy3T3v8z02ckBhsj0Ea8b0NbgxgI+QsBXv1Iug5vE2gJ9akSsh8dzabstS
kiYVS3wStlbgzRVEKXqbCJT6rKfpnkAzfkmoYrhQFOoVLBj/WvVlNTRF+dzWhhf4
6w8T/ZLc4a96KRIfa8FuH40+kvTgYKyhOcLOAd/d8iYcN42SjvfC+zxsgAs5+bmL
was4qDAUIsTgnHtm2BQTBaresYhkwv7ipBcW/XNl/CI7KMk2HvHMj453+oUt3YmZ
kn3NKTfHgjYCoHUC8O+V4uYwY8Z5pQuXYKxvIdq7UCaS8JvyPPwQ5LObwnL8Sx/5
zXGQzS3zpKjEm1znXc8Ja08axYYNG28W5Ms5ljCPH+EjZhygDhUgiPU7JuvWOARY
/4nXtiFH6uBRcs7JBYksqi1KazwJhos21hVqmJ7hFc3UUhSKF4tNDPTb1jg+8pPJ
Rj46dudoYk/HUCChWm/6Xlq587ssBdu61IVv+HeBE88f6V+B3TpeMXBpEqpG5fj1
YfFlUXot6Av50Cu/79fMWIS/4o+O0hvOE4Lzd9J6n9oko/1Bk5KxE24dueyutDpH
sHn4mHLaZ2ZnEKvuwQfPGTzPCOk2VbiCN5CHqp2a6JR9yeo7Bf2DUNteCCnXK5/S
o8EC2Zj29WCYtPkE3kuwjhUsemV8AA7aOSLOpnms9lgLOehf+Kg6qzk4L0SEW1vW
xl5qHRBfOjhuymbzeyun6CR363r6kDmto0wqr4KXC/JwO5g0Hafj51hgIdRz9uTV
4zNxD1o745geSjLCJl6zivk/fcGFXkQVbGCoMmxf5PcN9IfL47M3yARGAi9xYsii
dXRzGzM/sJ/w671+QF5hnMeZphInixrJR29wxFspiAsFnowidLnOiDwb/YTFWo1u
CSose9inz1OIvHcS2SZlmXf9IDmhxrFmTZemHl/FXhuZwS6Vpb+L7HFjqhGgxxsb
os+snDXJx0miYH4a4dh+DN9y+67jhDXnKQY4Exttnv1i8pn/xaAhlx3LGbI2HD3X
TD/osj8sNYue1Iq+6TMQyLouKet4viILF9LBw/niSRrZb8H9BZMGmsmxmkduEuOB
8OmkzEUTb3PqTu8HkvCKHsIzkzsRHzPl79ZKccP0sBsmGsrCK7L0dqujr4AcdkV6
YVPl00nEGS/JkDTW0eFWxl18ULGC2ZjMXnK5Tp3jfYVZvVqeSe/n1Me5BCny4iwc
PZ1n+FlOxC73gnZBJEQ9WNx9HoAHaQzAFggefancFfRuiEHJyM4gzIUny7J/gzfg
kza04nBWqGOM01VUkWodcWjkqHGrojW5wzRR9TR4QSADx19XTMf+ob8nsbVqAUuu
ABeJivfY9j8qo7bzY1UAwJT/OyQXTEa16zsyKPr5H5+PcvD0HiccaxGL05an4QJ1
J36jWgfGSrc002r03QRb9q4LAJOJ/ikw+14hIBT3ea2pJ+MvrldnFPYcZFDCa1ge
kJojlO0RzLq0rvh/pEYFymzplxzxk3BN+I5v66IzLN0PPErDCb3KZcOJQN5MNTGz
+UtZjEqQk0OuqFox36r0XJvzO72H4CXBUqE5OYvkSJOb4HPPjRAoGnDvp6eBXNzh
iEXkgzT9M1TC4N3ecB4OlPtII6ZwTORJ35QVn/6ldvEtzvaloE6/RZaeJuMuoB5p
4buywlHtjjVqe9yzfrfPHoyhcTQWl9I0/X0dzarOMzWkw55NUyopl87GzoBpCANO
Zt4jWG3OaZ3KxBRjw1uvgGgXkbmNI+SJZlY8ssWoGj8b0uZguzDpAQCF0zOvlcJK
6hQycy5KhTFQlL1kUQ+XNFUbItKcoClJWBXkzZ7DWYy2YAxvp0qbjiqPu8TZ3znC
fZSBF8TVGa3SUgjMSqfr9UjpLU+GF4rhjy9pntjiffPLu6VMU82p5C8P5Lhxxm11
4pgrICj9iJ2JP5oDncPcY1mCrcgcFlL6s1oQsTEaz394DTsReYdYlme923/9qDSJ
ot1b7in32W1oKI7mcUkqdZ0sDUTLjfpaEpWrcVedi6F2KWJmvmGyIRRcoIEsjpbD
4qLden1yxdhZG5Y+Yck0eNPQ8pK5iXFk/38rxncXS8WsN+zN/wQ/M1SoS9vIUNra
M8zGACH+ajX+4ep3v+7xirizILuG41wf4Cdw5p+JJSDpoZwbSYe61WQAFD1/gkJi
lsn/B1m/8QAw/xsxycgpIf7jQPpcj9Keu5kCRHOqwB6RrcXX46wuLlFx4D1UZWmF
et/F0v+ztLt/iCJbEMPXah6O61OM5wmOuQZXzk+Tn8tncMPiDLSkcWQ1l5uY2wJN
9laFmsRc3vLdG6SwKMSUrhubu2Sg9liUAxbX8WChQrHjD6xqEfMU7ZzQoszRSh2d
s1y3ltEkLDqoWLP0ZSNuc1u7Uz83QWV2532aB85fk7W1ArWrtuUSNXsAeFcu4Kgi
POD8kja0ghX4og0+XaEOAQ3iORsoNbJ5hBfOKND9SHasPde0EqUZx74t/clIq5MH
Xv04xvf86viFl/VTHcoaR0wOzYARJMEMfwjcalxKMprX6QUy9tPdLtl0QvbZwSjY
Da+UjL0YQyNTQ52BocUa4rV7hO/NQVSOh4jhTcIL9EzoOUZyPKbnLwz82Ghgy1Vk
QR1SDqT9CUeZ1NxockZ7waXY6lTQZfWfOLYzijik0RkZ1g6KH2uXuPWGWeyjzFz8
1eWQVoJatMbP6RxETC5++on0FZr/C7+JCv76Ql9ZQW73oh1Rovu1JhUM4hDIWmyA
zJiB3R3JmAv3SSltm9emMnUCdCCI2f8vi0tBJM1WYsebq9bkWAwT1PDR8vtkz/pF
rN0jUJqJBQxks3BL9Vmqgb4EGbvFR1ogKxhArESzzqAAUluTtYlUFuOAhion4Mmt
Ko9Ar+zPh9Zr+zFWdCxgMdtBqy4R1V1V4h1m3xz9BLmWyDOPr7U+0R0/oxbWPI82
g/2/23/rJlOp/wmLrwVeSHOq+zGvU1eknRjcYt29HxDTgRaY33fjwNQuXHAwaZAA
6lZCifih+dUKjltGqAiIP+pmv7pdbqasA2WLJKD5RmUwWB+1kcEeQrhZ2TBYtVxy
0ZvAdAtFXmHxf4C45c/XbMDomiXZh01zUUeCsd7S0wdkKTFfns/JOdnUSl/1/UDw
+0LtGwNFXxkZ7XZBUY7Wg+AoucvbmiqSffgF+IkGuhE2d73lKgithcexqGjI6r3C
pU/A4ImyGUj7s/oecWszvjf7dcShmIo4hGCi1NxE4c6oTEETaSQFuVLHnKg4tHSL
NebaHo8s0ihqk5d4PcjoUdUdd60C6nKXlpC4d5EgMPldjL9vNJ42TLAKDOM0F3gV
LlGFGLZB6lbhObP/78QlQSBDxKb+9WdoE1GhfzNz7oQPrElpf5t9oikN62XTTwxr
UpZLCkZTlPwZidF1WhJTKgSbaoS2ozRTE7nZSXAm6QZuHnPDXEYWQMUhEfrwrpog
nzSqnkYW5LbC/2U+COPLqsh+9xPwsT/mRk6y9Szz7ySF3tTPLwD8g8LL8DnwRWsa
rg8ppoXI0/agXBA+J4/g+ZO+Wq2YV7LJXDkv5IMOW3SP2QxzxM4DvRXHBjoRUiVq
mZi9/tVNP1sRMAVAP60i9X0ooo0Wo+Z0pNb8nYrKK3f3B6cA950HS9yqzT8foc7X
7birkMWyauGtE5F3IpJj41PTKBZmcYUShJe3WcF7C/MABxPaAc9qNNzjTeBIHvPO
mO2LhdretPcR4yzAgVv/iLTjP1fBrnhYSeCudTyKLYuPoWAYyE5CQV6JFzzOcSBi
fmfwU9yzI2hTi32bfj1RBvrhuNxOZSjDp9xtUeebbCwPCNXaeAKGNTQNfq2+RoXF
5gXkuZ9smSEZbJc6340aV472lWXvXCcTa6nROze13TjtqWwchaIicuYKT3jKJ7la
QEwfDwHq5sVno07W2QjvAvBOEMz+qCFlQ425qPZLrPExXt9SjlkKMjufabsBkZJ4
k2ICgx9ISPHCUUZ8t7XZbpwp5LPysrZijrhC2IgzATxU1BOM/FfV0zbtC0DZuM/q
JyE0vWjp1PyYmGw8UXoZHzlcjD3419X6qQ5/F3J9ag2vQqyw4dkdcX5uo/ztOac+
hHCldTVcbaBVAuuGh7mF0MEbHSvwrcf81sD06ObjppLV/a60ncOpD/riRlGYKCFr
7HlE0xFK4V2Ra4QLbmujQVMbQC5Ry1Rurk5Vdz18XjpbBucj822qB8WpYb3BNX6Z
Q26tE9pnC7TFx0va4i3seJA60rkIr+Pc7ZlKorvn6iYpU5dnwkLo+JAxeVYJ4dzK
xD2lCmGJjT7vxcwmAIAig+rwJm9RRx9vghMr7Nvv5OnljeQ3BHb+EIqksChx+uSi
0fzK8dc/LxtYv1DhdBqZR5iyRa1HNBbuRXv+H4jYGLNIEtorfnzIYKnkGVxVabBD
nEx9WlUvlDMqafkIreu56Fwzz1tqZnt38Z0QJEUgXD6BxX95l8bnPn9W+rCwBZHK
gNdZtUn3a9bmNBIGf5WMXzuS2bbRvIA/KlW3/ZVmIOzr6uh6IrtZQJM7zIKSAuJ+
VierPxpZNUZWIXuVjSmqtx1i2lVvxqwBDqm9yX2I/V+rfGIDIHoz/qtXSN6pmMa2
NXo5V4WlneEksz1ybaQe3FB/WrGk4vJRRreuQrKXdzrAR8XImMdZQm32+BMj+u2s
5pJL8s0TyXDtcjxsrGpxNkGtpb/7zQ8ZxforiJWwERLxfaGBWDoJJYo75xHJ8i+h
YdJiqZXJdzbmMCCuA1ZJgKH8M0WYdliIybeUIruBJ/PArr8Ak2MIOmVXZrzgTfN2
K3moabjmrocE/HiV1S3HiPtrI/06FnE/pnJQBr6DY+MjByPZS2XD5M1MmC1jKWQR
a1rK3DbAnD2O98sxh/jHdeNYaTMqFkd2l2hU+7mMpH0nU8c77Xcse7mA67AQSSjQ
gBcwrAUpfhA6GrPbkvdibbc9jUlWI8eWoLCWAFzKoCK1uk5JGwyX8IjiDEhCByfP
8E1skmAAc6AQ0P/4lC5Xvzsz4bEIu5w6di9A9RwDY7OKOFjTdW8sJJH4owO3SkX2
uqRDN+gZuOYrsdb4/uost72TXzlXYJNXezdiis/USmm3BnnxR4f32zNrtUGpqymF
1bHTZhUTApUDmKQzIH5M3ubASDYRfi7HOqF8YldTl6Qlr7tDNS9vYF6K4YJkOIld
NnLi8oATMPSjnx4jdeBr/gDujwkuvGUAdsxpvJQ11M9tWmbYOMupoMrYi4HPBXYe
BIOTBO35nEidLhKM6h5HySfNN7NUsOLvtcdFpiXrJu6FeFxHdwhwSEGj03W7NTTx
6M6y7Luuy8byTv8yEHIkzU+ikEYXjexE0K1/yT3ChnwFGESH4rKLo5mMZzPXcx2L
bYPA7ZTpslqSXF4X+H/el7DXwMIS0aW5uhFnTUUMoV87Jn58GkZzID117S4RJ29j
X0fBh+ofige+G7I09YIB3jGKvttN1Smic7M9oAi6NQMq+dVlo9/RhdyKpeLtNdWy
V61eqFHIDqhVEpqCC0vbpxNNBpWN0XungxOj/sii3X1rKYiTHWhLYRBvoOPHzoDK
Q6g1UAhdX+YxC8kilnroYxhh9Ti7t/I2UeiJ2aLhZMly2jHf4VRMSCkhXKxnHyOK
ToFaHMAL6RT5nGXMqzi1XU4mQm214LYLWicEu/U3ww6gLKbBIVmG43YYVLGK3Xq5
FPYCGGAQiA9mGxQHldWR7gLpyT5hlxXwV2yt0HbiulmEyPtcTErK84FF2GRd/BIY
VOXGjKMDsXjzkDn3G8rO2knf69g5s7UBPucgDfUSZfpMMsrWn5rpiOX4paDxLmEC
xalfCNZuoh2QkSybBis32tttx2CkZx4CoIVv9BxiTHEIonqAe9z7ZKlKaeXm5ez+
U4C3O8cpzdEz/NlIjmIHmlQAkb6HIq0yWikD7sbMNSa8CJ/Cw2kgicyczTfXl5P0
kPQmkq6lKHF69mjK5g6YDINcGr4z9mMDG8qqBEA3phC6GYZwd3Hf3lpsblLl15+h
O/lOnPy7xnn4iAcH5rjaJcQ9N4HeS6Ds3vTlK45GV4EcvC/Gfa66QwCU8Ry9gCoK
UUcsPsVxxgs1mvNtEL1wVYzTAWu7pn6omL0wn05MZZEubD6bxB57+qAlM22z9asX
V7bX0sN0Z5Jr+EvpujNQGciEEWcemeCmnF5J5XOF699mf/FuVj9jzRMQwUh0DIKw
D4FcjEqCoNCNkVdsuywPKAmLHlQcfpjZQvSzzGQVB0G5IOYS0fmX4oPBbdP7x5tM
k1CPL0DvFKpUKhKEf9oqY7ZYt+RGmHZzelqN4r8sAUrOLXdTxijy9c5l5nIHoBlE
3NOzJPVJr9+T0bc5syFm6DIXJcNsYrvwiaCIs32rmEKYCt2Ce3jxR58rmqlf31a/
kvkijaU7pGrarAZkIyEJlT0HVCHXBPjZCYumcxxTOJyK9CNyVFfcFn/44da/3MW+
7HBgTYipJblBo4FLghrJtRbpwMChV/crv7ReIH5cBGi631OQ3zxRVphStuKmJ1o4
kl1OlTyxI8cZ88ukmuEIl+fWuVDvh3X68XlWFv5YQFtvC/nVPsAv+mXZ+45JLwxR
rlACcVSSPUW3FXXSVRRRI9QBu08zx0fEius51kpjLYOFA+HaojgIaxv8EwgdCSu7
stzanyTX2SM1b6J6+WBKY7qyMqnifUorpZM6wkXm/jLF+NjbdGjrTvSXmXrNL9Ra
620Feg4rDGyiPC4DRtM1L+90+hnNMbGgJ31YjI7MBr6UPgtVpCAVDOEMyD3oCFKg
b/R7aVS8ovMpb3EenQsR93HUojwQeV7lZAzI798KVPwNxfELRNXS57wV4yDhFQBY
F8qtHDYQs3DJYr7zZnTZclEOajyVOccQ01mdpdIJZKkuXcpYSB8X/qtfBXhEQKfa
l818XcWHOtUwRRU23xaewSm6c+BKTJf1kWc1Fm2OIzg695uzVjQ9tTyT1i6jcHuL
ARIim1Su9eFoHlBonX94zUfmLIUG2VgE1KF5giXNBw9WZLK0dsLEF3/u9fGnuh5N
Hm1IWZG/Gsc540HKkf3JlJbpURiGNb3VYcEavqJrn5hNQP4A1z09pD8q5obIY5L/
1BY5pM0XC2K5V2q7uxJ8KkvNYA/Zymxy+RU0KjR7fvbIRwEWFyMP3pt9kHE7EvrG
A2ZzYg291iOfaVUrpmY/4kVl0C5mi4ZuBFkVCJtXjxnnxJtpT0cIKrnNpksdFJnX
oM3vHfPWkE0GLiPBoZiV+aMeBwPOEiVjShcoxdw5oEPzLhTbzA+IXFerxmUSldVE
P2JMVZpG4huIzZ5QFvTtd6QdsTRFmcaM7UClaXCgL2ZMmtKrPqX2AYlg0MjqVqdp
hfh40f6L8+koryPJ729pw+mmGCXhwzhZMJsVW5yi7z3gSoEAZko19liwf61OWGTP
jmi84r3X5Jn9kgAFWB54SQBmQxo/Ar1//oRj6IjI3RFUrhLHgqGsur0zxpsSCAik
htc8E485RRWb1Ensw09ol3nfkJAt/24wSCbCK403o9/tnqIyJILCO1BHjNv3fQv+
fLuEfNiHuSFuIldDhCqhlJn0TpcM4ndsBGh8JUP/LjTtbn+UVRJ4Z1wJ6sqlcnzl
Xz/ihxaKnRxBObSqdsUZUpZAipyKU2MPsHs0iZh3LVIWuCeBL8VViI1QYF5p1dFy
1iOGmZkAPoj/YBf7MMhpN2gC3+sXfQdejss2x2dh/bGd57l03MGOo/0gKYTnzLpA
5+FdGRQ/BMY+HD2mA93YaAX2xvCrP5PB2PheqYRL01cxygrBO4YFW/bcigrsMerN
FDG2SzdogTlR2RuAoIzUaCpxARdmqhpiuq4spXSgor2W12cfyaELOdvRG1HSy08R
6W07RT+62Zoc52LA9VYiDY/UBAHmO/O02MQp1zLuwZFX33J7prnauLrHzrf86SmE
s+BH6/zpHjgfm+09lHbldFL/t98Aj+/jMvzV+o1/0uyUOZCwie8iy/n3VVHP23QO
H3cxn5MBAon3nUs2kTUMEdYUH7hCtafVI0ygAf/FHnUWWZJ2PLef/1KOq72VHa/x
a6O1h96U2ytrvgjN4ypDfCxhBTJmIYoXI2/VPxxc/jp6U1tDDaxYsgYCkOq/7HLI
oZhgzlPgIqFY8vsT3ydMzONQQEjagpDOu4KVVGXSwQBOIPZbxDAZUw/VEzEa+2P9
/TiCWH9J8+UZuWES4/Ss66JZpbud9ER6fKga1CfXdIhq+WS2yZ9TtW8RZ91Tak+K
AHfEGAnpIGMJHsdmADYHkI34Y3vTaWj73fLSS/B2qZa9a/Yt8jLSXCJT+2VWqf8q
GRJQAJ2NiWZUtQZYQoiuIJzY57okcGt+ybO5PiblvDr978F9fa/0shkDCB7XQbBS
iVV+9lt9Q/M4bhC9fPSpGwXZJELtQI6+ZPczedZRyqam72kgKH6qSiG68qGlsDSL
wvPkaJFV85nQYXgIXREpZTQZUBmFh1IchWXMYiTzMJ7Hxk000AayAlTJ2oaS7O7L
0kZ4/LS2u4MYWi2RxV2XH6QD5DXbz6tDieiHPXZxw3GJfngDfQcVYOkVFx6zJ1lY
MU49P6VJxsXKdaGYzbWFBgjWNdZXQzDdsExJqvY6T4SqOjub4gt+P2Z1ls1raqBQ
sB8R6LsFQUDDDZDMRT6FoMOCuouUIo4WF9GnKYI8daH5SuWYA7f57BQ2B8I9F+Pt
MhC8sT3wer/0S8AaJ3T1abSR/WY6+529y45VlaSK8UPodRJ+Ga6T+YtvbSBVWHe5
PDo67tfEESOmybL2UadpozmKwl85dCT1Tv2ujgIIJ/9OAu3TAKG9oc8R7Of2joCp
6I6aU80Yh4FSmRD1j6blpuIacqn9dYUKp8ckMaXsMPLI3CHXzjPWBsdFX0g5dTR4
1H5SKGkbdkVnkmihcfoVb3kP2x+nZDGlNcQYcITSpMXgwy4rcvEUZAhpnqcn/954
2gu7Z8oNOZUFvhv9icjJe758OR6ExXR4pi27wx3u863rqy6RJOaSwnTV4B+bb8Kh
s29cmk91PiOGcuobr06pNwiTGL28+ob5wbSb/1K4JD3zTZoJAr+GWf2q3v8pi0hr
IpbsK3Z2Gr80OWqyeVKcM4YqqPuhq6F1ruH5VJeYUxmYBkOfXy2dKAX16cToB2fc
p0zZWA2uce0xWdjKOvg/zoAuYg+CDP75xXxPoQsF1J9Z0AUrNn684hFLVEgNIuQI
fBOHpB72szSK6mSqDdOEwErRl56HurwFSRFpJBb7R0cTVmm7HAY9EItDSulUYdcy
OayMyq1iZx0wVPLKFYNG3x1rZZ47UshYEm1/z7H72ZcdbiEapGJuNfeecoIGIMuk
Skt09qorYAt0oswkb9HPJT0gDeIB0EBG41v7KMXl5V+FilPwPXWMmOKOphVlUuSZ
VYmdFVN/l9iOvlabjpMYaPZkpndP/fixVxo0+GVJVwFb+W43gAC2vUuETka6WM5B
zFZBJystjC39e7zbDFegYhM2B9tlyjcnYHsLas252xNe6Topra2LfUDxQLOUnGke
ldaMES5ov1+Ucbbscur5frn7QeYWo6QfjtCw6LaWhZ+dE3+wk2rMQqkHDBiq6Ea4
tta+hUwfeXIeSUqXqa3sr808R/fKyImxLuhj6RE2dvfjdugzhfWiqs/gW97ef1LQ
f1oGG8B1TzM50bJPIazkJ31EM99UKhw4cJ8E8K+rDzcD8Bqq7gBdF9UsgO7ePiXU
nD3CQ+jMpqm/CtUlEpa+HrO20su4J9AQII5hPgD3Gnt8yD/b7UnB26Mo4WrBxwTk
7JaFD0Gcjj8oZSExCeF02TkqwI0lueWfr7+yt72bHeLlG5HWK+XlSZT+WnWv9jcQ
eWnl/RR1/VUn9JzZy55VhkBMMzW5qpnugZNVCB592OsDNWpXyduAIi+8Lc7Rx/P2
SghHazjVBx3eFMWvWJBlGcmWgZgAXyV/Cv8dVrUmi2Lln6Ef5PWtSaInmW9x+fOi
4y9k8zCEUT03tnxcQYADz49AAlS+Dxr1B3YF57jQHhgqSXS3oq0WrA+091/tz3J3
5qBd6mPV/GIdvDIAFH4WnSyJjnlxMJbt7Rdb8NCjJkPV/qy23M7vmtcVfnwqbCs9
pFuSZRu46PAs0kC0LS9mXqgUnOjDk80wugIung8WEMFbmGg50Q3Iym8Ftbo0F+Ru
qxcqTYsoqu9N3craxxrfWXrLp9WI3i3XY3eMaLn0YchmWuHhyeKkpmFHQZS/wdn3
TOHfkubBoghOI/rswl5YSpc+w2SfSbpQ7AIggcOumzKKjrOwOPmkWSr8vZWbO+Jm
JWJEZ0Ajnr1HopOG/OTf0cAWjpqP9x5fiHktSVMxVJvzcm/Hfw/GGgkhoFrCedaQ
qBWJn+f5Wc7BcBemV+KFqWPq7D4dFu+zt9ihPPuHk11yqu4XUUjD6qCXOkMOkPB0
KWP/dyzHeqGHcd1KR0JKsmV0y8paym0TNJIzhRA6Y3CXUEQR7Xpz5Se0AOahNPo8
5ogfbvE6OiBQH7KG2fXV7yo1vHDCn64ovHiY1+IsOOrvNyia0Pt4DLsrdeMCrLXC
OSGfOF4DOxYjKZnKTUtbq4UMi4qyWh0FJ5GPcHUrIKGIAaaOQqh6WReykVUExC9s
K9ddd5iAqrp/zy6FRiSKivPCyoMiDCJemcG17+pwoSoWLlYHMV+akfRUBitULmj5
m/oXOda03T9/oJTTuziz3yVCnFKmrwu5zHGSQ4fq6YZszyYwMMYwfLTIeIt9Ttsv
ddlBPoie6roSMgbd2TL0EGjVo08GtjIri/H3iQ9NcZonouX1wt/iaQrwiaqYtMk7
ukG+LWafSc+ZT3Gt2HFjOM7x496lXQuwl0+en1qsJTb7d9WsthwlPcwNCKuMB4r2
ffdnqbW+NwkNLv5IY3+spcUM7mcW7X8OtZYo925117NI2Nlt150ebnUcOfgeyG67
PvyChM/eh735GtCSeDu8zvzmM7r7MpdQ48W2VlSj8OVprv5Ti999rjtt6SZPbbWm
GGyTINo5MtCbM+zhyxA/d0wy81fdKGjPHR09+vLzexKOMia/pmek0wpfysfQn2HK
rwsev/4u6XuLJsZDtl1nV8HdSZp/Gr2/jEpJEnsvVYvcfKG/G8Qj4AhvES9RWact
udo0e8arKavw5+8r2rVSbWZYAcyzIYf7yMdeEqIlFSpdu7ZRMIO5Qouc1BXDX7yT
QybB4pEnX3Y2am2GEIg8X/WjeZkTXEFFPij5HkQ+VvPrn/EGojKxnGkooUWQ4fno
fPJAy3/S6j1zrWL2bKQebyRLaelq5d68AH9/GewvH+1Eu0q5cWt2gfWgDlMeIXZ0
erFKX4c6qvd5w8lp91kab3mRmRk1xlUbAR7bFCAvgAjUO2QtSH80UmzORxJVZD3L
79YBBGnZ73UbTy+/soRUokyVpUNDm78yBC+QlyvhqGvIHJhIMUFPs+VwERzI3HtF
qPcE3qExg0FccF8SCerbWgAnuHayypXuI3d4uFcgqHQWyIYWPkb5qt6X6w+U0zh4
1ifwZisZeomnax9tGW0PnZzMeG5FCZC/qC9xwGyBQm+DNZrA91UahOWEdIba/WPN
bV8LRFhYYla+uZofaWfF4hUbhoU7ASf5DdSsHHA6en863rIsQU9gSqMxTvPkaWtt
cDn0QzM+ANw74io6yrR5/SL0aepq6exOGeKiYOECYiiwdXfqhMi5E3/oNkuBOgp6
RoPdieAV5yoHE/n+Vw7wIcrW7ZvXk81fWLeFGdPjZMLgJ2R0oc6R3tmJnBB9/8R2
6NboCBPyCMyT8X2sHdaF9Bn31xfawVKS096hjgEfXfOC6Cs5FANTCZne0bNX3xFS
nsdrBz4/hCjv3rDdLkLP4d23YI/IRqHqhewGLeVq/KWQa0MURGlmMygoSP0IQu2C
UbNg6NlezjbPkNVs3+5fX4cjEIK0NS9Hu0nsYLWS3yb+vE49w+VrP5GuUnC25gaU
MD9GiLwzCpOL4DnDvRGIJscCPD5+f0lmD80kMP1Igc+JoatRWc6RIEeywIsxYusz
UF6KN/yk7431VCRgwCqUj8xL/wXTe+E1O36ICj2/Rx/DJ5l6/I688A3M+AdGfwFR
Hdhf2eo3+RBSd8pdgJyRDyNDayidGZIOynUBp1gbruLB5AXhtannnlQLqPG5Sbwa
IFoRqPqdNQKgQzU3xKFa0a0Oa7kNfL00wpapqMsbFFCQe2HinH8rCWgN3i4G4JFv
fubUf1hTZcG75K5vse8iL2mqpT2cA417EP4bTzQTH641XVjz+mKyPPcoq0O8ByYH
qZqthFkgN2YEbzNnWmQBX5okYn0lwNAus7J3EZxNoMD4MVdjd0gWvzBQ5q9F3mTJ
As9YqL+Yp1y3OuyO7eln9a5Q5afI5h81nmh2GiEvEdwKuAMuxRxfFcqL7xZKfFbG
Ddlak4GSO5sxJTMR+W4MCacrQlzpKdDxNY64obgTsYHNaM4eDNkPTPSKKFaEBeUV
hXPNEk1NJiOT6JaXzF9n5z7ayDIr27FkKXFK0oy05SXp3Wh1CCpbX6u+WNaa5nKS
Ua5QgZ+F2M2qzeFi3NQ4ZJTd4YukYlitLq/pQpj3cF6xxR2tESdz2NdM5CdQ92sx
gy7S1dfT0Qll8BQjCLUlabRePNlSuVFP+oT1N2Nl7ZHOHkaQS+owl6kMxr3bXkra
SgzMWOh75oWNI257iM4xPtHwzzGqtFZLJnQL+BBNcDx+Zxn6rkdKM6sSoRAt3sYM
LrQeaICqptoP+N86he6hvPx6sAqGuX1qVNlsoUlF9woblnhouI7Gm33TzXvYwj/0
Lnzk20nYlhWbkOGDH/dtDTZQe8vUMYjhFtr1dtcu3E6L7Yxt6TYI1eMpBBBwWvhc
7ge4hCkVWKTaeyASp3Xc7IXGEgCeAOzdF1Oc5Y5mwwRD8nLvkkX7bj6AM80Ndy8q
fBJdPzwOg9QHlNUBOSCJF3cGtVYrQRKpQw7lVZQ/lH3VyB6WFvtZ0rmD4sgNjINu
ESGuLe4AUTgdlDBkXmcpqhcBVhZo6XJ/vRGGHNvW4Dpww19lW5TZ/TnvqpzO5S8i
wUpVmBdmc83BXluWlHu0ySLqlnI48wqs0ikrCZnsDWUAbs0pHpW7Glg01/cumGjQ
Lk5dOwJoAs4pGMkBhC1kyAkpbSvQHIULObl5CbeRszbERFNvqtlwcl6ohbgj4Jfl
25B/8FWCO76WvhvfNMK5KBG+NVozC+ShejxniW2HAkOYaPVo5J9Z14vaf3d6+mt4
Q6pquzwBmO12bYNQdqkLLraN7KoJBcm/gWTNs4nBbvilaVxC1BWUpNi+79KyzIgN
dkl2r/KjPR07DCGqDJYp7ZL0X6nPWOw5AnU+YIX/ZLMdAl3QF7ht/hKQKcawX+pa
n8dz/SUxkbdmH9LSUplpyj2GZtQ+tlUCIr/zYEl+sg4MWNwENaWoDVm9+Yz4XiDl
DEnX3LW4MhyXIlc9R0SpEL4OorzNctl9GGkDnXc70BGE27Ae8BbAjzE7GbP3geFB
YAXrNyNPDUfWumUTcQkhFAGKBxitem7g8ipM+QNtnwRAk/JzbkpSFS8ZH1mZhxtf
I8PAEdieS2D7Uk+ij9d0DtybEeO/snGpXilizeDD0s0z3FCQYZRgfem3fdALOwsY
wX1cAhMpDW1zKV8nq1Pw5Pd3gvz9BvSHkVkqANVzkAutGItXV+8W7tfAdvLBDoDh
X1xeGxs5tCWPOpiUWJOc1w==
`pragma protect end_protected
