// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bxzPthPJ6Qa+LtNWN1hE12lOE/9KnvZY3iap9/W64tnenrtaKBQIYVAq8aLIctkh
ylhEwzi+7bjrnNNQm0vVcWhfu/dLsk36qyL+5opkOamYXR18GRQNY4yBkWsUY1Nz
cNNWhm7NnK3rfjqBMEBXM4Lsi6LDWNZCuvc2/2JAP1o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8576)
ZEMLzEnKmMkS9yOw+oXbblFj5M8svDh9Urb2YUvRyfUzyiiQ1SVTNNjNkP8wcEk9
ZCB7YAwT5J9Ae2lIwAZDhpll3usbWPwztVcfvz+doHMfpexYPWvNd9y53AIpTHbY
9JMuP/mpXPqEyQKRYq44UME9LX45MP3MXn8igSbgk0Tbr4oYQ2UIKMl1v0W8pwbN
9LMb6HjH++QKqugTDCF/+XDK0nZitnSkkyssih/wDSmS8VJS3XNvDMU6GFRM4qMV
B3xuz+ZCGWn2LmZinFVsl6VuNWsNwzcOR4xCUiWl3lcPVkmTqD/9j3DR+Usk4qcr
tG2DrNkvZV1SkVa6/7vJdzzOaG4cG64GrzQzh3Ni2tB0XWILaGoKW/4PI0DaHKyU
SW1xp4NuSL2OxTFqeMyQVsZ8dSyjfqKbG6wxM2w3vMBO/E8WFczpCsvWwdd8amXm
XBDspmCl2BavIV1YhS4CRdlsmv3Y0LZNkoULhkD5eJ/A/X/vELmliu4eijRosuH8
J84oAedTokINTbaX1nkkS9yxvkj2MjIneWZNI4S/xvhrVombmz7tpI0aVfLjmVQx
fNn+HoEHXq4ja91NM8t7v+dUeUyXz6cZoyOZOSLKpxe+3gBWZjcp9TI5SUfNcU+W
Bt3eNRqLxAGrttjZPkn1sea8eHniKVpiBcPq+L6+JIf/UN6SguWXgDuZSsSboI3Y
NTpdX4K4JlWAtHCp7cr7aJ3UBVWgbMVnC+GvTq2tHHHjpnPfZnzffgErsxgE/9mp
WwGcLl3H4I4NrYQFzLrdod6HPoTw0ccDILIYi7Z29PKVqd1ts2HCYX8ZyrRYn2Zl
Jpvqdk69juxk4VLmPIRjxqdK49/FxvmbbDZWMt72Tf50wW4J8XIGxQzTPIKCRMR0
uI5Qhw0h74xlpfuFcNsVRmEj6SicmdyT9HA8yKWtKBuJOOPC9I8bLxfKTaMZi3br
zM4VCj7ycPo4RcpxgVGUBJ8N9scZFJdRzYrWgG5+j3T+piaS5cF1ouKfjziRhl6d
hSDu25TPvOx5jS4/K2Lcvv7BgxD/fik9xZblim3J0PuMorOrlwF+cgipP8thCZST
6RLJSN1qybrRjTrzInv3hRstSdMeryClTXq2AsYCt1Q2MCX/jFNIWiVpZnLW5h+z
e9RGRcMM21Pg5p3x+xxpjgsZzinenW4gGx97Buw7+wuTVNvd9Y0IVY5A0LZh4WLp
O36UdSB7G/PuIG+bX12jE/aUNekeBHQWIfXX5jTsZqxjRny1Wo3fmgo0RrSxHCMW
d0xiFBSzUDb8dK4sh0AG0a6aUFMk0oXVkzmIsbx+KIiPmX5HNTzwdNgv3EQA32e8
+aFAvcwGgbgOHzAw0Ck0WCc1vUKFHQ5/5H8uMKBXXySa9TU90Z5KhYSxPpIeJtgL
mV9BD6Y+Rh/0pswShdBcPlJDuGArOrqZvvyGsEL4Yot5L1VI+F1rrTVMn5xU20Qq
+paRY2fooqlN34Pt7M1d5Me38MisBb+7fVVCiXq5txgBv1xUp5ZAga/AVv6HCk5p
v0ehHcqncMTYfHg59lAlontW67VtvO68Susn192hkj+4oiZf8FLMEtQ0QwAkVUUl
1SJo9jGUYlyrm8duyRUtKi2fcsuQZ4gO5jCrH5g+iuJIpUXt9lOQgcLevS5gfnZo
usvPGQs72uGpFSFz99thBEZKZHUHe9wZVdmU9lcWpJZSGGxleLMgPJkC87+SpP6T
Gmd2aj2y+iSDkuYYuo9SNCrg8Fmi449Xp64adXXkRrjisbRocfueYHA5774KsUO8
+WIlvFUFAHTkBWGZDE5e09prCCG/g6OhCCtj/f789C57Fk5KtlbwkkEXXgzdhQxo
afSQn2lAylxaxnbaaIJRQ3dom7xU0zt5c/WFV9Lie6dYoDpfGOAHOR0/HbwaHuS1
WXppvKQnezddoVxpA5d7q7pxHYgIVawQLx2WhtNWJLgfVhV37mwJcjetkK92JjlA
ftLJJafOywso52d4sLOhNSpSiceqzIiAK/RXS5y8rL0uSZmKnfr5krR8DAbhYiQH
9bs6mo/LMUAUye2wBmB1utfjyfZpKITqlK+YLU3vpyGConGsY86s1lBs7yXgZKzH
qbXfEYiOigVH5Tbeacm5Bcp1dNQyR2igAKy7yYeIVYPegPGae/OrG24lQd7qdDxt
R71x4xCzmMWJYeglUMKMwdATFG+g78kk3OXUDzA7Pj9tI0T1gCuQLdoRc8v5sMf8
YTzOr15gOYgIkV9j+yP9r13FYaF8Kf+pjOoDL3PnxcVb0z4YaNQ8BfOYAP+KiPVq
W7J/MEMX0GCd4TUJa18BeugGk9MYekvitde2rVCtJqfYdq1yBJRXeYbgB8ySKzSX
rGiNnm0YAbdNLhv1aHuy9oEYQlyYfhnR2j6wKIp7U3FqgHPvE7sxtt4OLWVZrVS2
tkOeMCOiSGTCAdVOXEYd8N/zO+51GYP1sQoT/HWt5ly9I+aZmZ7CxVyflNYX2bcw
xlv9bQgAWO3qmaEEZaxCDPU4FcpEJim0anNpXkE2S11VADgr9HraVbS6jsS/OpJ5
1Wuh+Gbp23p3m+Xu121mK+Dfw15S5j/Eb30HUb7weYZSqvJzjKbONOfqceYeGnIg
jFMy0aHKp1N/Wu5skgEjdbBs5WIPPcFffsNF9gyuA/NP99EkpJwvh0um6fy10thN
GcboCCDBcvEXlEGx92vlIYZ3zM9awfaF5B/8GCUloRrkvAlgzwsoOWh5kS7OEOss
kYRoDG+g2RFEr66rQb63omdu3dUyH5nKPFh0wQwStcD8klRqt39p4+x5CTbA9IAe
fJSrPPzUsUQAFwZJyULAZdV1dB+C/vnVNIgfbJW6wH6jXWFPEBcAS6w3oExhcN6b
0KvU1Y4JZ5T+7vA853CkfD0d6QnZmDq0gjWtQs8kfa9GOc5H3O8W7jnwC0ZOoAiG
dt+ko/FAN80i4rB4yMTzNQXKG/dRNq7f3HJTR4M/Vf4Bx7ILsHS+JuKc2vDV6yuN
yvyx94vGHFGcfkJYMNG2Pasy3QbjKbppaR/FclTt0APMTWiGvt3cKwgXDmdX0sgB
JwNVU11xioe/BLbMxDKTnd6pByaOYScTOzm3mTQ8M3Ml9sIuqVJw8/yi2cDepunk
SaW4IaYLyxV8rwUY+aj8WbSQ5Otdsy0gJCkY63sAa4eZDcUzNvfFjxwcnCenXM5i
y1vCqQc3urCxjTZpGyHhMBezdyTROsW3UKXgCPVsxr7qvNT0c5plecMXOPqIe8kz
7WDUBd5dDSzn48WzFfBW7uluIyN9tqtjkfTFaFPBBbADisFfBqN8HlwxH8SOuRrk
udgtDiG1tSqi+RkEDr2gZ9ZTqS56MM6f5A15DDM62n9geQIsWUDlresDdlwQ+wIb
3IwbosX+6ARKqN/WiqtofbxsnItAaVnizvz+XApy1dnaPj7RYP0ZsSBfBXaMDrzz
aoakYMstL31I/EhGi4FLid2B3cX1Kxy1zWEDgrj+L0dmuE8H8lEl3CE51opNU6Jf
kY7sKjGUhl58FjFbPTOoQZtfR58O604VV20BR7b6uxlWM85vvlvnqGt/5UnGyvZW
3Xz9fEMDreS7nq9vkjLAtWTGBMHs0K5JsJj8wAtIJ8kB0OMzLTtYc7paS21fHATZ
MGzziVmQnvouGvcpZLneLahOG9zAMz8EstMkzANQ4UF1PFLZ/SJv7gOOCmW7nyUB
gfuhGptwWYjaP/g+iCt5v78SUo9hd5JCZU8o1PXtcdb7xncB0j01JrWCXzJ44Q0K
c5vU6W4a7r6z8XxJjxggTQ1YPVWndPkVDueb6oCksupsd20Ezz97ilHlBoBZeedH
DJxlpu/tyQzE18r0aVT++9mZFxTIzNt0vN+PYq1yuPjXPvboJ+NsKab7SXj2lK25
+SGHii4wjsFaP6S/QNjvVly1fDYoXggmNA6lYklW2JCzC81IrPCFGf0EUWuuFPLX
gBQ23/xu3+Zf9Pou+1tWCB1bNoyvjGLbKkYnvuYrynmGEJb6U/ufzI1iyb9aan6k
tc/enWRCNZVlWS7q7JimG6mKGIOPoalzev8DNaDMFgWFw+w+78IQ6PY4jbPZwuCo
toMjM2wQ38mwEtO6UqzzdDZBRaxMtiMKPiuuY8ixFtOrucORQu3L6Op7l0+2KZFl
77qJMBFdavd688dG3MpwmZ2tcCJZc21bY0Jv5aLuYtKBVQOorN+wNgswbf1eTa/d
ZWl1EYrfZcrWFGGe2CxY+feCkGjOJ9nxrhX20nGnSYMnAh2TVP4aEcNe6UHBh33P
P/RFKpoN4FBXx8CvgoYALoLLiiFvVTKwwlOAtHexFXsEfeHevVs27o+1lvXxHWc9
xHruCOn0062GOH5NLcdQ6YOLAsZueNyE1KoHTieuXzclB/2mkRcyuuMy7FdY/u9z
QECh06P3UDlKTBvt3w7p9ZM/Sb5j50hNvS8KtmVnp/0Sr6XQv7UFAWvSNa1hflSs
ku0r5JGS/UXUPHOUUscrvO8jM3sQ43p7nkwi24hrZazdiKVqujTKrNhTaubEgyg9
YsIdUuXPtNKTynlOKGecmi4yB5qcy26kXtSn37TzZG9KE/NYz385E+65GjTRvPHp
Z3iVBnRIKgTHJ1prd99N5rrLo/9mRlfr798+5cbbrNz4Xq+UV2YGrQyLXjbruUAf
vj1VLZ1/MfdUDRKw9iOXFK1/cWMJInuzYWY25lXzDxGF/+qy70PX0/rK+YOJ2sOK
XPfOHYcnpQQJ833Xu1c+NOQkxFqbMhKfPUgNMLRgzcxI0urt+jhfXwxbUtYdfI5a
Rjup1CeSOchID8gajBs1LuyKQXJQVAh00Xr7LBSB7pglkGQeQlGt1iB0+G5G/Nps
ksia75863JhO6uxkw1Ehwb3/FW8sZmVMsT6rgoJE/SLC0d0Ej3DeqBF97T/BpdLD
bXJMEsFCQuo1QhxNd5O1dwQQXhpLjMtDGwaL5js1XKi2qx1dx5JWkH4rfhGMoMiB
nUvwZti+i745jKnC5NDC0UTYiee9MVcoCGh+5nH1On0cuaqusKGDuuH7DHoI6eis
BV6q0XOkRGwJbYNva3/wnBtdwjB7UG7jnUWkqk0t/A7NtdTrFTIL2z3u8uJayZdU
U3uNTcsl6sWUANj0T8EC6w/j3gws5W1SAVObz+ytX4gs8ghu6m4iAwMUXIGj6kpp
2sZwnhGdee3NZa9xp1jChg0jhbYnTS1MxYZMjAeasLqAaoaDh6bvpHRqXJRhAWUx
opJYIc/e8maZtLb9HqqBJo4ipHYXmQPbYRtN/PNR+XI4nB8ECam3VF5KWyMenDR0
XZhe5tc02QJMcLbsEQWvEAUikMjKUolXEZs7vMaU1W1utcupvzYf9JhFBMd7ZDup
T0nBRCajTC/MGqE3U+CvJ9U7CrPjqngEd+OV8Kh+48QWxc/hN7MQYNlWT5NFtNhA
c1xu/0vUmP6zF06WmDSNySsChXJ77ktgwcQnEvNlIxpswHqnUBeIcnzgfQSQbL8B
+6oEp6OeuRAk1zOaQaDENM5U9SGbMEawO1+/4S5LdDq3oq+I2gxDtAW6IksHCN9f
QihlD5+CqH13ze6IRwhvFZKFjh3XYFLwm5Cv1FkTOHYUaXk3TYfbaXQuHroa8EVf
QsC8aCoMyudyuy/pLmUpD7LBcSncAl4RE4G7dH2Z7oBlnDww2TJP2n0V50gULTVf
MupoHrX3jS2iy/dKNTBhDAClOy2fYfT+hi494RYhteAwhAMuOvBrljgfXhMqWcL/
ot1EffsiBoQMP8p98+Heja30IgTuZ/rIxSFhgD2gVb76pwHAz5Jfo0DGj5gB9Hmc
c+on+DEatAF7GspluE4DGfTHRMk7dYTbyN1qK2seOhBXHOhuYND2mOALeaFDUjmF
sm8ZSaRET/AYRn+AHMZZU1wDHiZyopWWS+2yKGJ2cumOvMTEEj1/wEkBVSCHfzZR
5D1a0yCli6zP+Ps+8GJyjZDRJ6MO2J0m/fnvZ01bUN7Ipef2ymVyGLSGx+6+wUTY
JceWCO8nwS2zIwlbsA7jn+QNLVVLjoiK9J9hh6r4Lli5tfEHNAmEYJr8H61M5ex1
bGXPlHBkUTyYhun3fhjWjY58neDBqqPUDXqCXwaZzikg81J4miMWZdlM4cIZC3Nj
HwHwjxxpNDSZVGurdDuZdGXLQDdYL6P5H0GuukXNLoiK9TFBM0cHj7XxdhFS5rix
OzCPq1jpEWVDcdqaOQy8SQbCqdFJkptwfNPN7wgT4A0sZkhG0/LX8PRWB4w+qTM9
AgXzcG+KSju/nRU/nPuZNbFdJpD7aEIYY+cb80nLchBBpjc4Pu/gVmuH1kZlHjil
IxHFtsnKd4Fqufbo8SdNUUeQdmUsQ7mjOAMp8d4NbQDxyeqmN5dsuAqBySaAIGa2
SCwXsWpwixA9b9Ng4jPShZ67dyGTG8C1MC0jMj/uYtbxNgfgzMp5Suo7dG38ulIl
YyMViDWxfXJ5wiBINgrBFjXBaWcfIKtkJX2IAWVe8dYU8euTcEtw23DDCzA1hbG/
e8VheJ6w/VgaWTe+Xa12GPEvMZErp84n7a/g7ba61jsfYoPaEfV/wdeGAX9agGKV
hjVTXz2dAXu3JVkHgE3DuJK/JVcN7WEVaODwMmFLzPibbr5mDy67DGn5xonp3NIH
yHqELxYrjxnF7LH+B4FnTFqkz/0ARPYfqdpDSwRL6h/tEAG+bSqC9vItCbpjgT5k
9WmmJsZyhqstcOcjZatA00q+sdX3pWFK3n3m9HU+qcxWWBHOFKnpICa7e1aIexHl
69sWCaDZBbDTzzYeGgJuDbiNLp5CkPkBwThugrcNdtaveB0QCDEFpGRogzC3ySQl
p+1ESREbY6lvjN0kojOAbAgbmv2AMRHWinEvwbxHsWDBF1jPtTc0fb5A2Ti1s2cv
VpD7tGr++1AUkswcCF3lzg6zXw9YkCR/mUFVWUZWEN5z+2efc4u9pUpTDIT0Gtbq
srRFct68rbPyxSjw4/T04z0WS0wxDz/tqWCpRFLS0a5jcu9Wl9ZGZJZhjsM3SUOb
i3El2FsCaUGxwVY7sgX75CGRSBHETlsqC66/x8ZgMujopawSr+mahRA5IU4lQaoo
WcJEXXiXBBVbpkLHh5jZK2F7tqcxLA5PCAyHvOiE5t6BeEwCHT2aEr/GIElhXkqJ
EFUDlv1hq/MyyS+XsbHVt6yimn37lDkcD/0FOMQHp4AKD1hnyro7hnQZF5sccgiH
PRMb841F2RO86ngPeaq9ng0rTEsr58tYCARiwkvpArkBE6AJ2FZcXFMXih6roLoc
+ZAUaZ/5AhQgFWl5imrxDxHk8rbLUgEA/2UgMcs2IKSvxb0JbiaAp8eQKNIi+hTm
Eskh/zuWQWDdc9tDSq+1VMhUIqkSdI+KJgZJ3vc6AUUujUw8pCqyVCaF6xpQvGD7
ZyFcxaqCzWYziyw7RXVfn2G9YwZwTY9AG8DPGlXXMN/DhPiv/yRr79yP2wRR3x5S
nLqJE8ACUg/Um8XJ6+67U4mUMYBnW5cw1o5amDkdxg3MOXqpcnwjLsVbLZIEBvPy
vgnLjvVNxSSpZPJ8YDU571qUSNMzdH/dvHUc8rs4RvpTgSO0mCKyOOvNn/IR85Zd
9Jbj1MsVeJX1yYm5ILGgftWBk65MSt6ON6zSkSq8QZFupbUHNlB9mU3x4ep/D1CW
lh9Y+SBk3hmeYbHJsxNAHkVMEQe5fezS24cVEqdOYcWSFxDk59T0fRbpDy/A/ieC
iAK8jZWCUedXdTxtxYCA+vAjEezDwZBBTSnpBj0JVyQPPNhMttwl55+wGm4lNt6q
tjrVIkbRznwQl/CSqNj4XbAOuTW433HG8XoSec8o6Ihn+MsuanbIdfNHbcKk47TL
cRwf53KeUUxzKOFpB7gYzGSd29zG9ammEbvoxXxZ6q9W1XkavkaRuW8ZbozDInP+
3IbsODo+KK36pTYJYeztJIA7/KesSjlHJ2/wRPM0rqmntzgeRoIxM9TXYhw+Cdb4
DPN4lCi1E9e6v/1sixeFl5lvkbOCqkf30NsUU/2+mMf1G+hz+JZTxMg2y7qVBtCs
YflOc/H1m89Xcu3/OuBydUyVOLj0+ZXE0wFKdsntWjCILQmfOKzZft6cN2F1uUZs
S122rLVaFyrStgRmsBnco+Hk5s2UWx5GnOuAG9e0vSqNh//68DEoWxckHoTveB2i
VUj21WKjhQbv/ybmljjGLWrcgwyvtfZfn3aJYQc9dj64KdXO/j5L6ugBEHd6XGVe
3KNKYtpikPYjvpltT1qjolRL3zg3wPnJaKM1MCe91Lp+MuPPKueg1Ljn0oPeSj2e
7HL65O58hLCaO3joYid5hOwXMurqOFyHzyeprSyoAHvjOzjk2vQoiLXftjey24hi
MyxmlhVjLVWsVzINFYc1RqJOG6j5XzsK0fP3xpu5lxPUl757o+Rl52nMc+fEAAN6
+w+3040xYHSu2JWU5TlPBT/Q6LvW3w1rekd9X9+jPkSJW8RFxJvuKVaaGGAbC/an
X34fVxjbqjW5sLtdGHiLDAlynV1IvZ5TIzJGi6tWZ5vYmhU9JPFRUCSYLOMoiHPA
fLvaK9G8pi8eFh5y375wJrfzl9kSbOomYCacRErXG/RKS9Mzy0+CJHJ7dVCHbJ3W
bnUjyfS985csltl2FR3Omt4OOMhIsRq72ybx3x+C1Y9vquET9gzMtAPryeWGSPdV
OhbWDMxfmsy7wMh0CXA8Y2BYDjVtBl/rJiN2Nw3SxjVomJHUJZHKcbsGnMcEZB3X
puETKF/oOKWl0MB+772Q+gTyRfnqcZ1FeFzcC8QnonE4KsbvLZ2GVp2FkYSsUV7G
nxf7gFJWp0Onj9i5BZVQqHsguPk7o7lAvCNiD4u5jRfidcTIu2VMPu+tG5o78RYv
p+9D0z2I6m2wmA1Gb0KQJwJYg1SgI+GnlwAGEjX/Y4tHJc2fJJ1j9ZX1LhA6xsBm
WSedtSTH7JGwcxvAAUvytHBHBhjdUGG2DlLHHjPp5x1GiKAoYxazuo89ma++Yif4
sO+2ugbl3gydGxoMDEJqA55BUtmrikJbx02XPQW+EBTTzgVQQqjSd87BGA5uYRNX
4WRBtpNIfWA/ZBIEjW1DZWvVNeRrfnFePWxJw89xiBUVvcrI7u/ApvdkNWYNoDwg
+AKcoYz9iwTJjrqla4gQl1K/k7rP/1WSIYoRjH74KSJaCTVGZT30Zy29zM6VPRJ7
YhJ+TE03GWdv4/Unj+VJ5EOXp9rRc8kspZG3IHbt/zL2gprp2lpnWSrMS/3mYzN7
bgtrsUhMVT1XB9rjFvu1NAyMyZ5kXPKAFt5byYOWjyKbTRGgFVDWbUhNaZgx8lld
ZtebwkhEvl8QklPDZfd4MHMWAqPZS0oKbFr2SeS2EZNepSIuKpKmlr9KHRvTsiUK
b+VbADSpHYLCDwocvJdc2dgE+R1soeUQ8tbPtDFOdlTO+ggxtVZSZznh9zQy+S43
asCqksh4wo0j/8FrRsrhrCiho+2uXRcve5D8bIFxT4pDzv/GC3HuMgPbDbXjak7M
6oDU2MZcT9fkETCyVTNtW4Sk5quS4TSNlSCM731IfKblA5jNYrf1ERL+Jru1+N9r
CU26T7gjRzFYqg9n1WWGkzEw5vk/KWHkQGoAGHSzSkeKuxhCA7u/pCk/m6QwULb6
1iEv8valgNlj1TvlGUj0xh8H42rlhBiUQO4jOrWLnC7DprqtFlMi9a1piX3Z3Vdn
P9Qkx5rUwEMaaX693+FK6osPdSQ63kkvHjJ85D8vzFgfZoB1mTJTruHiYuz3uB4M
W5F+BULK50MSKxMTklmn6KuKWa3TAKz57e+NKwq82RR5GSzsONgsWEpdXCy8mESg
XfM6/4048SRUWGHfPYB0wNEZlXoPFPRF3MO6YVGABFUnKazXTc0jIPN+EGIQNpSW
TyrYJwnCSPrQL6K2+6xCVL/vXRGiy8AF911xlARFaf8CT3FOQ0LDzE0BdAaGwLTK
mpVZyt4C7tXqpNvVs6BzXPjA9Z8cb6MA0JczMQ9r489R40nKZzuLhk/S+mTS/+Nx
lFncuOrjSvleLyUj7HQKMKNgXrISuA3WpAQ0bpw4Ch9kRXFQKJLmZqpHBwZfgCXc
hQsinXFJ+gjSyUaJdQVCuX0TgtxvzK19hb9v+gP89sPTx8OMhjK/YSUoo+dxcWZJ
DLhdPuE1WWurMzFO6QzmXgY+Aigzs8kiQJzlH8g57lM3fSMYAeFhpFBwcdc9F3Iu
4fqP4pue5t1eXRKt8lUS6+tliNCAOWmpVpFWH7VJGeuhvUH2+IDaSqFrS4Nes56D
FGphVIQbACADexH4vw2HNx6BIo4DjqIgAgNjpTQJyWmpGRXCjxJ7Oo5zacjRI26m
4o+II/yNDpQ1+p9MIriM7SUSvHXpJrdArUZdhGT9ltG3Sji8D6GVWkk1BrVG06Qu
VhLeZ01RMw9lGgC5Qa+mnkUM3Bd3dkKNxV7QB48J6OkLytQj2sHNLKtFkl4gweGm
8kurxuVVL17OOhgZvKPMNJeXDOpCunGncFJ/aczfy2T9/fiwy6STmKBaOly3+x98
gsUudP9jf+LzTF/xKUxoo+D/ECdhAkj0tGl+sBx6swb6guGOZ5EVsMdA6mFrlg+K
Pr+/4+cNSzw8jmWipmwFLoNRkUzAurqPqvDji0eHeYtHGB0fAdKcM8sXHREVw5xy
IEHyEtwZ5B+ohoa6Fo+v9mKUCP175t1xpdFUWSjkQ+XPmWFS+kfa7ber8tIoa0cI
cbjiwUwp6tkiDQi1FUr9AW9xRq0HDuVOMBDj18FSqq7bQJVFLqI4fpXpPfAlBkAp
tLKUHpbQwSFxltbo0FcujPLCA9ahgeuvxBuJUqB1IS+c7vJP5KzrrN92WyZu9G/7
c5YOrF7Uoni6Iih0L/EO6NrxelKj3L47RyxUODBWaVPjzZmlR5QZKCrlriWoyQCn
8QQ4OtctYJJ/a7dha9I5gQ7zQ3GcnwTupVNig1Wdtizi8XYvn7xare6axOD0qas7
Run3vKXtzoc4AgznKMYzul2eZO+X6KRW3gB2rH2nKOfuEiXXFcBbFV54g2yXtpOu
LAmxDU/265ofh9BQq+fVcRkwz8o2nnF3MSuEw9hW3GdlZwTntwBr1BmTYEyPs8iy
db+N+Ws2x347yrqEkUjNGsodulq2gpiehkuZyA+X65br0lJwzeWRcKL0ltgUqXxz
T4sSydzJD6k/iwM4nA3TnXufhSpA4l7+BDioXpMnW4DRvMufaXbptuZSpqblI8uF
Bq7p1uJQxM7Kjxr0EmeWhE2qxLAd/3xyHlPUgUlRnnrwIjQK0ggrazmqEsowmppz
hcypdpI+47Mi39dzfZyypF5Q/aJPTa+LKS3yf3Q49tFYO5VY8Eqvxo7fV1jWLqo/
kdjmlJ9lWzp9KRQiBqMdd/DYb/YUF3gSZg9OBoaaysg=
`pragma protect end_protected
