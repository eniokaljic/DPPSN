// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GYNq8+JmGTkSYkWZAVEsTOA8m9122yP1sKavxb/iqnmnLG+a7QwOp3RtydQe3x+K
mu3OUhCAG9Chdz4f+MAG5TzP/TcrRQlOTdMI2qGpmlvBlcNqjYsDQfpltamRq49F
jbTHKXu23ECkxvPzGSQXlu9ocaWjGHupWFPtaGAF2S8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
18e3rQ8/sxiNqHymI57AFuTuZbMdItFSFaGkCE23t80sr1WNXsNApBxU4VXFpQhc
c2M/XVHahxUxqkz2xLplsaH476nveQA1ExM7r/kOKJ0aeKyV3BYMhCWBV5pufsy1
fQ2D6HpxPZkvNxroYsYqABW+RrDJsTOGYJ4bqsgrIOV6qHww4t34cTqaXXZ12iW0
p6nG+wv3SmQ0qOu+vt9mHX7pH45reazcKk9Z/08pLmTskWFNOjpU9AQLgpNJMMxQ
6URRBgCA9RQ/6A9xur3nrJhMsN2a6eyFcTcQyjrOa53i5R00Z7jVIH9MnINXizWq
lACqHuXqn9G7L8RX/+Xs2EAFbz/6UIhAm3hQb/zrtVBx10cfDWagTuzn4pHssKte
PSi9VF0qCXkPey4kLtJg9M1DLK5zY0Z60KDzf/pnTJsJkABuqa9yuqfxNw+vAOul
EiJsXantsPju+qPh6G/MVpIMwB3nj4Eev5+LfcoqbOsfmIrN/fBdNvinMILTEfXU
rIeVK+caQbFNvWyYQAMmBm+RBcAwHlKuzJn9QmP4Qtuejy0YRTsk5h6NdTQUHQ81
nkNCZVIkglDfg2Zu2+aldMoZ1IV5aN8ZvHlrVD0D2bJNeVgDt5Oxb/T2tMzXd5LS
e0ni/a0fJLxhbRUzv5ZouPjhJxpuxEXpqjMC+IOa7LsMTh2Izq6C02Bsx8kE3KTO
yNefu/bo5daYs48zBeqyL/JBm6OX4Xay3oqsOA5RyrP1x9YzcppH4BzdyVCg8M4S
ZYTy8YbIPzllRPOOokRtPJcZDsyEdwUSPKeSnEXAQVkKclY9WnRZfNF21+QyRR7T
TNXG6v2nFyS6aBFE1D2hsovk/hz37p1aNag4LhAyDo9AZyGZgKR8mKFYFTz6WkbK
Zi35OCItDKY52ga7oea6Jn/FaRhtDLt48SuNBchBZXJkYWZkwtUD4AaMoBDBNewm
cjfc4bPg8K0CtaPOMXBt8AsNCzVQu5Fd2NV2AFnZjQtPnNuMZ8bFaoIbbfgluYjS
itc545nv+8FggvVrMCsVgCwSrpwvzwwPVcu16DPnQBQ+hC5rFDwiCthJ7wj2uQE9
B6f4QKjDp3lnQEq8r+ZCjk9pAqV2DYoIQLvaGtYBordTm8Cvk6wiQ2zGAE/HetHy
09nkGdo8LU+ijPBPN+jQy5OoQ/8tZKLq7ZajiPj3rY5gfJ/yzhaOWgLncQ4nhLe9
FgLAZakIPX/mBS+RIUKIhNIjE9CfiTHJEY9rr6j0CQkUz9c7OegIj9IcQlH2sNRd
jXjL5dah+29ycL6v4dyIaqRzNMa0i+G2YH8cs4ACmrvGUmj4We9s0xAwS9n3k1S7
kimXZdkkfog8bz7brXbL5LNss48ozhKiGnKYfh827Y6wBHiqFimhwQknL5poqE/R
g0lMY3N4r5LPDNVFQhLtHGhs2IkY6c6MRKtFrjn0Rt7rnBm67NQV6SsO0i+LMv/v
aDcXDKRNflYg+SqBthvBIhPOWyqaWZFYXRYp9h9MKNMa9ywcSBRss71hXSjK5UQV
H7kcuNQi90l5Xf/y1NNza/R7u7oktkPS4IY9eO3W3gd3LgVZ5NRo5/4fvRDIhyge
VY58XDklBaRmrCeJYvClwyWp52wnG0+GE4A52zP+6/hHpqfWMFHxfbS79tFD3UK2
6HY59mfNBSSGQWpmvCAlEBMZafuEVQBYuz+fCaBJFCEIhiPVZI+VKWh+6fUeN0OQ
6vSDzRpEHfFE1oYbEWJ9oJKPfT19ydS9+X4WCWmVJnb8JDNOJ8hyEhNZVcwiTG+3
HqESVUVdscaFb9Nlg8OAF71cGuXAB6SQylN9CWRUIXiLwpV1TgM2EpjMj8EtRGSh
Vu8JZwCNKcb5LV25haP10nUq/71jsfDQvyyzFJIagqVfHC6xA1bZKZj4Z77J8H33
v17IXpM7D6hDGRMrzCs+31suoSdhGt7KLiQcZy0dheFSxT5muL58RrmbH0yrbioK
wEbut9v/t02m8kMnxbnP4KbGASwUug+tWGlo2MuvBHUNapAKYxJzWSZUUix8uStG
LCD38BeZO2l/+MNLHmcl+OyuyjbEwu1V5JmPERJRxRXy4kpUl73e2f2vrHhVw0Dr
0fFJ2uNuJzKKNWSs8CSyd9W0ZhPuJiDJi7fWUHL6ox71VLTjKcbEM+3W7OWWQfxN
9V7Ehpin+8V4Bf7mLfHjQ91Tl6RWyraLArkJ+kr+kK9H06eTTnU0T3vTkoSBRtm2
0kBuiLtAY8Tq0425jRtZ2/wr1vujo99qaQ3Ivc0jJfPA2x/RRpRnRwIM3u1Tx4M9
BahHBfVcRXi8FU96vwCqhptdcUEOQXT/wIHDKgqDedwZzFve7btTZAGUd5H5I/lH
qPnr/TREbjiUTstJhEllxUagTm3tfUZBjynrN8xiDmAA6iGAUn0KVrh8Lc4EbfNA
0CpytzTgJfu60UEFmSZQD3Ha7uWzzwd9hPJEb6S4dpXrlfgi4G/awM26dHAZW7sh
ff6eP3FF1wF4s7Fu2xb0AqO976aSTWl5K2M3PbjhSVxR92WCY7lRal29BWfh9SzE
E4Kqv5wvKaeSq0BhBKKYNu1O7jgEYm6iu4uDX4xzhhWEphllTkDM+VvezkVmcaKJ
tJsgwmIIfcl0lf/tIgw97rGDgGQ9s2ZHzabwlM94ToGINQKgWAXgRwwfbYBFG0Qx
4UCXheSEzcDilaOLb0eIe16nk1uwJyFhmLqUuJhN2UMLyJyu+GRQ4ESFloPHC51r
HrqwLK8z254XIcmzzWJU4CP9W/fGdNdMUx1fU6WDxwyprRNrl457qhK43C1i6CAZ
zuRRRIhVhyclq6UN5tFOI6gRDSMw2OWFjeX87m5dmoDDkWAoU9so6kqBNLSlW0RJ
ANMcnPPwrChMxGWTtGDhhWkIPhaweTXir0fdAesOVQaNxTBnQGvumqEiEbQD+fkj
uCOq+aNobDsVyjUL5hWVbMOBCuZ1WqZmCvRJUidaIYH0VvHBB1C2vyxlyK4Fyy+D
XiSFOXWd0LgtpX0c1oISZhZMoOV14i+qTnZIArqp+Vj9gf8Oym2FCSnw2h9k96WS
6fqKPNcSEnXdeaaoY/ug+FBbIeOXqqFUeULJShBHnwoY6YiOCBA8NXB2P5xMO8KF
QslTrULPV4P5feLwyujzfg8EZ1vj15mzMze7wWle/N3xocC17CRYIz5EMRQqowXu
i+1eCXR8F4WfTZ5vSHXrXeqQKgSTMgPOHp5oGuEe/zx+bkxxB5XcYu8ht39NGQVs
KbGtrK/tTvFopNsfhjqwfVjBa+P++jbZHmRBnsi/COX5maezL/baLxyECCdZCi0y
a3VXP80kcgoIOqZiIW7r05jBQMY0SCVq7xxqlNEblboMqGX2FVigUe0U5oGTR/kc
DuVPb2bBbcYXtnsGk4KQWzrkwYVYKlVN1yDn4HvC/MEVAXGOoy5R5Xgbrzh2IzRK
ugkqoQYuhYEjrM0JimSTCZf+lXbjkIk+/yrgqvuE9AUmq0CIcGbBhw5mtNFrhQDZ
0IghF6EQVSPjejyiCrzoP2bgIUCUGFJp5r/VX+csKcMwWTtExIviyaCEK+VCDpE2
pvb4H3QxLK8DT3rQWXlNYZZucIWljVe8+CWYDN7dAZ5/H9Oy+Ik+6kZt1c1I/Cjt
P+A2xAcP/p0uE9t5hjViJSJfvlgcZem2tAvu5JJVitmqhwWrt2iK7+C7vX/igcYu
LK4Cg+566UZgrxcV8wJfDJ2PiNNZ/2/7dY0ZPFNNltK5VVdJogTb3aMXkJ/Iz4mF
JlqSZernUoC46RmhwLyHG5pFqC0Hzn1aWHJDIxFAiJq9SzC5bwqI6PwwfQ9/oZdY
xuI8WuCgx7MfTvpnUjebwqQnsHBCmQsEY3DqKnWPrgIBTRa4Ucj/G1nLWwPdUy+P
E9WcVrz0raaP4Xf+SyuGnDZw0letCphurEWgvCfU7ZTIlm1ME3pBFUuZArlMhW0z
j0sAxK4VUtHndtvcI9Kt4Fj9Ooaod7/u9VdJxYL/UwiBiVrkmXzOVxCE1wBeOvHN
WO1RgYsOuUPHbrQDn5U7SbNWhk9ragggt2W5/VcUMdI6uPKShYoIgXSSlmp2prB4
RdPBdwDsEduVQrCCO3cdPr5FVn7SPbFhPqEYZ20OJ5i5kUDBOUUCa+CSiAgY2Z4j
I2eSZ7dgaaflzzm2hMvUCqK+oDcYfK7LJnTFA0HhDqwp5BE5ZEv9T/Xv62U2rkFu
w4RggsgpJGDEPJpUGDoZD5uzlgOGNOJjxGbBWZzYcwnyGNJ6gCkZ6jZwW8/42ejL
8+y1vKT4SV0wZGLmSRBDLYs9i4cLn6K5x7T/1W6cAl+lL84giF3S2AZTQ25oM4Pv
RTfiYhkRsfys0ZxFkRrFlaWmTiGG6ndHIufvuqMaV7yIlBlerNE2lEcr77dCoCeu
izs7Bc1WDE/5MKzjtBiYNTCv8/d6tUFaC909M41pjh85Hf2DhVSmR/wD89lGlVZJ
VGshchBbhD+cddsdI0kMZ0EuQrmSMNWihauJ9fce+hUPP3kKoIccpjP9RzGcmHyZ
mx1/YnvWzC5CcGlsc3HqtTQi9Qnagn8wbMg+qPERnDcy+pMAa6yTQOkz9+37ywSD
K8vNyNLmo86fHW7FBEgNdPVBpDGB3Xn9jUZ/YZF7ZnR/N+e7+Og4QR7q1PwIlAHp
EFEdYhHe47SgI0/Ip2diM7Emq3BrMebTYr2iw/I0LGL2JCxO0bIwpZU3G0emoA/a
BvtiPAwwoXpPk9GWmkyaT8DWLdetfZHybcH2owKgmmv28Ltnq8t6wV8eapNWqwzA
3btctXG8xNXjn5h4iYIeORgCb1tvPMnGxBggZqaQewBoIzq6tLcVe5GTomZKJ6QU
r6qugn/0Olhr6kMCK7MaRKQhdWrCJfTgN61cOqaa0HzEo2C9yXXdGHMVwlytyNar
KTkcbKoN2canOLL6IinhQ/FkN3Q/aT+Tb7RoM4+iNvVAQ2tflLWcwMsi7K46bX2F
OQppaaRKd7qFr/LfuAr011AFUG5A3YsHnZ/f4QVTilLz7iLoq6BLT2FZMiKVla5m
hdKZ2ZJoUfr+CF15WJuJ9GUCZnctF/G/UgOsSjeV1WacBAlOTLoBnZ/J0Ix2XC3i
dSdJUtCE6HQ5OqaamHCtlBhObo7WL7EKnfUM1Do4ZkQ/8MEej9KyRoduGNuBxNr+
kg39vRFk2/nCqIINSoGHJPkvU8khpDi1oc5HLYsC/Pf0BEk2LDJGIqAcLvv2fgjI
M1D5nVTOVRExB2wkZUkSDCAzpJKshDKDAfKkxgjlXJCogZk/KjwPkz2AtbFgWAYd
LoPP7b9xX6mrSGE88DCZ2JpyiUeqLLbw955NdUYwHqrbi0u5eJcuxSk76kYr20Vz
K5vZEc1l5XWA+Ysydle5T7wmEp51yCozJQ3O+OLakXRKe8FoFwNNfoN/sQf6HlRj
TqVSnq6SYdbSeCfWMAjhjH1Crp2Fram3Be+XoSd6fp2GKKLwzAtBF5NDyjp9onG9
yDU/Tduo47e3lTUWhufZsEYY5E23zaPCLcV8bJKQsu0zyNG3251m3iMsMDJUZM9W
yzrY4buOquEwNRyCaFbkhIB6lCQkAM3uSUfDYeAzVuaZMlAQMoFBTHD7dmyGTUDD
Q1UZyP+5qGov0up4G3jErjawlrcRw82iQDexK/xckGfBCl3OW+VCIhYohHgUsizM
PDa3zCpseELBI1Pb5wW6d7aQOfhs3/hud4/OOOMjDDm8/BpwZli4w98W7kZQQJRw
in01QIckGE4J2zZGQM0SB+nTnS2SFBkjlw3wK0jI9SVzh62tLtIYDFvU0GM5syO/
mNm4mIXHzoob1KhDzgb0Fddkk2dTEdYhlvVw3Q8UfpB5q60lW+AmzpvWuMAWctWN
RkQDEz6TldNea4ferFcjHVFdW4ZBKBnBJI9pMDDReztFFAoqD0ku7xwuT1IMgkcU
WcMgDQeOG5b/22nLCJgvJ2Czr84au+h3k76HROaJ49AmNxEfturfHy6MTMsiwf/+
tMICm+51Akfa66WUJik6qTXeuo0meKsq0L8JBltFPQKC8IPwKthDWQQpJNQrQF+9
AXfuf58C5Fh52eIEBeTwDeDaYm7zXpsjsFsMjHMZkhSYIX+B4keAM/kIml5GO8he
mFF4rK/oRcTt1z3+U24q3BEvyg6ZAyhoKx5uotpPdlr3B2Kr1YJPQ39oJM67LmLF
HiwbeuiUXoZ5of3rFZ1QQJMwTpuHseMHG8q9GfRdMyp3pp3pfZMoUj/mlynjfMtJ
LtY24VFH2eBCscFG36iGsBkPPT7ypPlzBitU9G8XWMam7s6f7V2VFSMJHT7wOU34
30eriUSbEa8gmk8FTT948Mvjny7lVz3Rw6Z1v++vrr52B64CX2ujYUgdY/+Ow4G7
ryoB1m4lPRTQeoA2f/2vF3FVYAuacVEKkXwFfvZaEB/jTs0ax8ttkyzwDZJe8LYH
QA7/56TuDd3qNyb/X20xesqrwnwfPvHoGh4Ii33GJi520n/4xkbVJ7NKEKLBwerb
0a1s0Tlimu4qAKnJ1X0MHUpBQEIyzpO39h3I4ycgzpkC+VLxDbFlf6TJTOJX/U8J
EeBTRrU5QXSKZ0TQeSS0GMLO9KD4wJRvnu1FmgWGqnfvV6gTddp8EhCnGh5IeH6m
CeXMCMNM2zCs7hXGmdwEzTXxGNnZAIPdeHqsuVGh2qRRWNNwBDjcLwN4lA0NEvoX
+UH4BHsTsUL/S7EzjpB/+S2Y7WcmRKaPpeyYJ36UwUlbrUETJL6uiBedgqkIUj5a
tvvZ5FpR0tteq7VHrclTXB5kxVAQvcf+SWRUPMya967EzqOwSfc+aKT6dm8XpIxz
GpipnGDjdqEQSoWO50X8Ok4BoqSg17tTPTFgYiKHNUQoK0nzbbXlCC6NfbW2p0G7
LVVLMiKgNsefK+Lnqff90B116uPQF3HgET/3FpNrw9nn+JV4hhiRN+VVcBC2rDo2
ovElyvki+jchoGr0YTbVcjVDV+rQaLJBog3zjRLNNG74fHw8nZCNUX/Fj2qhmry0
xA0SQlIrh2Ir7O4Ixt344Es7QkTtUecRJIR4CDodOWm7k8mj0s1MaluxyzpqcuS6
eDIXXIPAL24HV+M+V39rpVwnX7LjT66oic7031uOf24SmxzGMPiRN0/hJIpeqhdC
VBvQUJC3H6BJJue0NnNsOc/alQrnMwjNdoUgumB+Ro8=
`pragma protect end_protected
