-- phy_10gbaser.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity phy_10gbaser is
	port (
		pll_ref_clk          : in  std_logic                      := '0';             --        pll_ref_clk.clk
		xgmii_rx_clk         : out std_logic;                                         --       xgmii_rx_clk.clk
		rx_block_lock        : out std_logic_vector(3 downto 0);                      --      rx_block_lock.export
		rx_hi_ber            : out std_logic_vector(3 downto 0);                      --          rx_hi_ber.export
		tx_ready             : out std_logic;                                         --           tx_ready.export
		xgmii_tx_clk         : in  std_logic                      := '0';             --       xgmii_tx_clk.clk
		rx_ready             : out std_logic;                                         --           rx_ready.export
		rx_data_ready        : out std_logic_vector(3 downto 0);                      --      rx_data_ready.export
		xgmii_rx_dc_0        : out std_logic_vector(71 downto 0);                     --      xgmii_rx_dc_0.data
		rx_serial_data_0     : in  std_logic                      := '0';             --   rx_serial_data_0.export
		xgmii_rx_dc_1        : out std_logic_vector(71 downto 0);                     --      xgmii_rx_dc_1.data
		rx_serial_data_1     : in  std_logic                      := '0';             --   rx_serial_data_1.export
		xgmii_rx_dc_2        : out std_logic_vector(71 downto 0);                     --      xgmii_rx_dc_2.data
		rx_serial_data_2     : in  std_logic                      := '0';             --   rx_serial_data_2.export
		xgmii_rx_dc_3        : out std_logic_vector(71 downto 0);                     --      xgmii_rx_dc_3.data
		rx_serial_data_3     : in  std_logic                      := '0';             --   rx_serial_data_3.export
		xgmii_tx_dc_0        : in  std_logic_vector(71 downto 0)  := (others => '0'); --      xgmii_tx_dc_0.data
		tx_serial_data_0     : out std_logic_vector(0 downto 0);                      --   tx_serial_data_0.export
		xgmii_tx_dc_1        : in  std_logic_vector(71 downto 0)  := (others => '0'); --      xgmii_tx_dc_1.data
		tx_serial_data_1     : out std_logic_vector(0 downto 0);                      --   tx_serial_data_1.export
		xgmii_tx_dc_2        : in  std_logic_vector(71 downto 0)  := (others => '0'); --      xgmii_tx_dc_2.data
		tx_serial_data_2     : out std_logic_vector(0 downto 0);                      --   tx_serial_data_2.export
		xgmii_tx_dc_3        : in  std_logic_vector(71 downto 0)  := (others => '0'); --      xgmii_tx_dc_3.data
		tx_serial_data_3     : out std_logic_vector(0 downto 0);                      --   tx_serial_data_3.export
		reconfig_from_xcvr   : out std_logic_vector(367 downto 0);                    -- reconfig_from_xcvr.reconfig_from_xcvr
		reconfig_to_xcvr     : in  std_logic_vector(559 downto 0) := (others => '0'); --   reconfig_to_xcvr.reconfig_to_xcvr
		phy_mgmt_clk         : in  std_logic                      := '0';             --       phy_mgmt_clk.clk
		phy_mgmt_clk_reset   : in  std_logic                      := '0';             -- phy_mgmt_clk_reset.reset
		phy_mgmt_address     : in  std_logic_vector(8 downto 0)   := (others => '0'); --           phy_mgmt.address
		phy_mgmt_read        : in  std_logic                      := '0';             --                   .read
		phy_mgmt_readdata    : out std_logic_vector(31 downto 0);                     --                   .readdata
		phy_mgmt_write       : in  std_logic                      := '0';             --                   .write
		phy_mgmt_writedata   : in  std_logic_vector(31 downto 0)  := (others => '0'); --                   .writedata
		phy_mgmt_waitrequest : out std_logic                                          --                   .waitrequest
	);
end entity phy_10gbaser;

architecture rtl of phy_10gbaser is
	component altera_xcvr_10gbaser is
		generic (
			device_family            : string  := "";
			num_channels             : integer := 1;
			operation_mode           : string  := "duplex";
			external_pma_ctrl_config : integer := 0;
			control_pin_out          : integer := 0;
			recovered_clk_out        : integer := 0;
			pll_locked_out           : integer := 0;
			ref_clk_freq             : string  := "644.53125 MHz";
			pma_mode                 : integer := 40;
			pll_type                 : string  := "AUTO";
			starting_channel_number  : integer := 0;
			reconfig_interfaces      : integer := 1;
			rx_use_coreclk           : integer := 0;
			embedded_reset           : integer := 1;
			latadj                   : integer := 0;
			high_precision_latadj    : integer := 1;
			tx_termination           : string  := "OCT_100_OHMS";
			tx_vod_selection         : integer := 7;
			tx_preemp_pretap         : integer := 0;
			tx_preemp_pretap_inv     : integer := 0;
			tx_preemp_tap_1          : integer := 15;
			tx_preemp_tap_2          : integer := 0;
			tx_preemp_tap_2_inv      : integer := 0;
			rx_common_mode           : string  := "0.82v";
			rx_termination           : string  := "OCT_100_OHMS";
			rx_eq_dc_gain            : integer := 0;
			rx_eq_ctrl               : integer := 0;
			mgmt_clk_in_mhz          : integer := 150
		);
		port (
			pll_ref_clk          : in  std_logic                      := 'X';             -- clk
			xgmii_rx_clk         : out std_logic;                                         -- clk
			rx_block_lock        : out std_logic_vector(3 downto 0);                      -- export
			rx_hi_ber            : out std_logic_vector(3 downto 0);                      -- export
			tx_ready             : out std_logic;                                         -- export
			xgmii_tx_clk         : in  std_logic                      := 'X';             -- clk
			rx_ready             : out std_logic;                                         -- export
			rx_data_ready        : out std_logic_vector(3 downto 0);                      -- export
			xgmii_rx_dc          : out std_logic_vector(287 downto 0);                    -- data
			rx_serial_data       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			xgmii_tx_dc          : in  std_logic_vector(287 downto 0) := (others => 'X'); -- data
			tx_serial_data       : out std_logic_vector(3 downto 0);                      -- export
			reconfig_from_xcvr   : out std_logic_vector(367 downto 0);                    -- reconfig_from_xcvr
			reconfig_to_xcvr     : in  std_logic_vector(559 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			phy_mgmt_clk         : in  std_logic                      := 'X';             -- clk
			phy_mgmt_clk_reset   : in  std_logic                      := 'X';             -- reset
			phy_mgmt_address     : in  std_logic_vector(8 downto 0)   := (others => 'X'); -- address
			phy_mgmt_read        : in  std_logic                      := 'X';             -- read
			phy_mgmt_readdata    : out std_logic_vector(31 downto 0);                     -- readdata
			phy_mgmt_write       : in  std_logic                      := 'X';             -- write
			phy_mgmt_writedata   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			phy_mgmt_waitrequest : out std_logic;                                         -- waitrequest
			rx_recovered_clk     : out std_logic_vector(3 downto 0);                      -- export
			rx_coreclkin         : in  std_logic                      := 'X';             -- export
			pll_locked           : out std_logic;                                         -- export
			gxb_pdn              : in  std_logic                      := 'X';             -- export
			pll_pdn              : in  std_logic                      := 'X';             -- export
			cal_blk_pdn          : in  std_logic                      := 'X';             -- export
			cal_blk_clk          : in  std_logic                      := 'X';             -- export
			tx_digitalreset      : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			tx_analogreset       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			tx_cal_busy          : out std_logic_vector(3 downto 0);                      -- export
			pll_powerdown        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			rx_digitalreset      : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			rx_analogreset       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			rx_cal_busy          : out std_logic_vector(3 downto 0);                      -- export
			rx_is_lockedtodata   : out std_logic_vector(3 downto 0);                      -- export
			rx_latency_adj       : out std_logic_vector(63 downto 0);                     -- export
			tx_latency_adj       : out std_logic_vector(63 downto 0)                      -- export
		);
	end component altera_xcvr_10gbaser;

	signal phy_10gbaser_inst_tx_serial_data : std_logic_vector(3 downto 0);   -- port fragment
	signal phy_10gbaser_inst_xgmii_rx_dc    : std_logic_vector(287 downto 0); -- port fragment

begin

	phy_10gbaser_inst : component altera_xcvr_10gbaser
		generic map (
			device_family            => "Stratix V",
			num_channels             => 4,
			operation_mode           => "duplex",
			external_pma_ctrl_config => 0,
			control_pin_out          => 1,
			recovered_clk_out        => 0,
			pll_locked_out           => 0,
			ref_clk_freq             => "322.265625 MHz",
			pma_mode                 => 40,
			pll_type                 => "CMU",
			starting_channel_number  => 0,
			reconfig_interfaces      => 8,
			rx_use_coreclk           => 0,
			embedded_reset           => 1,
			latadj                   => 0,
			high_precision_latadj    => 1,
			tx_termination           => "OCT_100_OHMS",
			tx_vod_selection         => 7,
			tx_preemp_pretap         => 0,
			tx_preemp_pretap_inv     => 0,
			tx_preemp_tap_1          => 15,
			tx_preemp_tap_2          => 0,
			tx_preemp_tap_2_inv      => 0,
			rx_common_mode           => "0.82v",
			rx_termination           => "OCT_100_OHMS",
			rx_eq_dc_gain            => 0,
			rx_eq_ctrl               => 0,
			mgmt_clk_in_mhz          => 150
		)
		port map (
			pll_ref_clk                 => pll_ref_clk,                                   --        pll_ref_clk.clk
			xgmii_rx_clk                => xgmii_rx_clk,                                  --       xgmii_rx_clk.clk
			rx_block_lock               => rx_block_lock,                                 --      rx_block_lock.export
			rx_hi_ber                   => rx_hi_ber,                                     --          rx_hi_ber.export
			tx_ready                    => tx_ready,                                      --           tx_ready.export
			xgmii_tx_clk                => xgmii_tx_clk,                                  --       xgmii_tx_clk.clk
			rx_ready                    => rx_ready,                                      --           rx_ready.export
			rx_data_ready               => rx_data_ready,                                 --      rx_data_ready.export
			xgmii_rx_dc(71 downto 0)    => phy_10gbaser_inst_xgmii_rx_dc(71 downto 0),    --      xgmii_rx_dc_0.data
			xgmii_rx_dc(143 downto 72)  => phy_10gbaser_inst_xgmii_rx_dc(143 downto 72),  --                   .data
			xgmii_rx_dc(215 downto 144) => phy_10gbaser_inst_xgmii_rx_dc(215 downto 144), --                   .data
			xgmii_rx_dc(287 downto 216) => phy_10gbaser_inst_xgmii_rx_dc(287 downto 216), --                   .data
			rx_serial_data(0)           => rx_serial_data_0,                              --   rx_serial_data_0.export
			rx_serial_data(1)           => rx_serial_data_1,                              --                   .export
			rx_serial_data(2)           => rx_serial_data_2,                              --                   .export
			rx_serial_data(3)           => rx_serial_data_3,                              --                   .export
			xgmii_tx_dc(71 downto 0)    => xgmii_tx_dc_0(71 downto 0),                    --      xgmii_tx_dc_0.data
			xgmii_tx_dc(143 downto 72)  => xgmii_tx_dc_1(71 downto 0),                    --                   .data
			xgmii_tx_dc(215 downto 144) => xgmii_tx_dc_2(71 downto 0),                    --                   .data
			xgmii_tx_dc(287 downto 216) => xgmii_tx_dc_3(71 downto 0),                    --                   .data
			tx_serial_data(0)           => phy_10gbaser_inst_tx_serial_data(0),           --   tx_serial_data_0.export
			tx_serial_data(1)           => phy_10gbaser_inst_tx_serial_data(1),           --                   .export
			tx_serial_data(2)           => phy_10gbaser_inst_tx_serial_data(2),           --                   .export
			tx_serial_data(3)           => phy_10gbaser_inst_tx_serial_data(3),           --                   .export
			reconfig_from_xcvr          => reconfig_from_xcvr,                            -- reconfig_from_xcvr.reconfig_from_xcvr
			reconfig_to_xcvr            => reconfig_to_xcvr,                              --   reconfig_to_xcvr.reconfig_to_xcvr
			phy_mgmt_clk                => phy_mgmt_clk,                                  --       phy_mgmt_clk.clk
			phy_mgmt_clk_reset          => phy_mgmt_clk_reset,                            -- phy_mgmt_clk_reset.reset
			phy_mgmt_address            => phy_mgmt_address,                              --           phy_mgmt.address
			phy_mgmt_read               => phy_mgmt_read,                                 --                   .read
			phy_mgmt_readdata           => phy_mgmt_readdata,                             --                   .readdata
			phy_mgmt_write              => phy_mgmt_write,                                --                   .write
			phy_mgmt_writedata          => phy_mgmt_writedata,                            --                   .writedata
			phy_mgmt_waitrequest        => phy_mgmt_waitrequest,                          --                   .waitrequest
			rx_recovered_clk            => open,                                          --        (terminated)
			rx_coreclkin                => '0',                                           --        (terminated)
			pll_locked                  => open,                                          --        (terminated)
			gxb_pdn                     => '0',                                           --        (terminated)
			pll_pdn                     => '0',                                           --        (terminated)
			cal_blk_pdn                 => '0',                                           --        (terminated)
			cal_blk_clk                 => '0',                                           --        (terminated)
			tx_digitalreset             => "0000",                                        --        (terminated)
			tx_analogreset              => "0000",                                        --        (terminated)
			tx_cal_busy                 => open,                                          --        (terminated)
			pll_powerdown               => "0000",                                        --        (terminated)
			rx_digitalreset             => "0000",                                        --        (terminated)
			rx_analogreset              => "0000",                                        --        (terminated)
			rx_cal_busy                 => open,                                          --        (terminated)
			rx_is_lockedtodata          => open,                                          --        (terminated)
			rx_latency_adj              => open,                                          --        (terminated)
			tx_latency_adj              => open                                           --        (terminated)
		);

	xgmii_rx_dc_0 <= phy_10gbaser_inst_xgmii_rx_dc(71 downto 0);

	xgmii_rx_dc_1 <= phy_10gbaser_inst_xgmii_rx_dc(143 downto 72);

	tx_serial_data_3 <= phy_10gbaser_inst_tx_serial_data(3 downto 3);

	xgmii_rx_dc_2 <= phy_10gbaser_inst_xgmii_rx_dc(215 downto 144);

	tx_serial_data_2 <= phy_10gbaser_inst_tx_serial_data(2 downto 2);

	tx_serial_data_0 <= phy_10gbaser_inst_tx_serial_data(0 downto 0);

	xgmii_rx_dc_3 <= phy_10gbaser_inst_xgmii_rx_dc(287 downto 216);

	tx_serial_data_1 <= phy_10gbaser_inst_tx_serial_data(1 downto 1);

end architecture rtl; -- of phy_10gbaser
