// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b9oa3kr1Ib6NL4w+QUs6vUVX60NX1zvMcDBDHo29MUb+vTAAo31gi0ClYmq/1wWX
EzwykAg7zDdgWuPe9JWnyUeGt/B6jXSVjDKhR+qSQh9WTFQHksvFT8RqbbHtRgZs
ra+QWXrY2BIcutIsMskio8b75AWU4Wv2lr9oy2SFHdM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 50800)
6wzDNlFBYnj3TWzWfkE6UkCFKIfdPwE/pYLz3a/i6qltzImYG+SgHT/hozyEvYO3
MdPpJl2Uhg5NmuXDr780dmPlOtR8RUjaZKq97nx6a+9ue02uBEumqLZjhADcsqmN
U454pJTlI3KiiDL5YgE168QfsqR1ygZGVN+2jT0LZKojlmNaUJ1c+9KFAbz3xqlI
nhNyz7BZAui700lqSNjWWx81yUKqtUHzLeUFFHQUPjb5Gl5hlOQ3nknyy041FLT1
qTHAunUoTxwwDRkk0HVe7Fr+axNzGQKi+VI7Aulqa2H2RenR1L31M531Id8wp3hi
caX9iLTV9b/xNYbC5M+GSf4GNvjrmOsYPzEmrXEMQe0zs7AnyBaYvQHbhPjH+y9o
6pADeDy9IXj5AHlXrK5UQNYM81cS0ASfRwmWVtTixNLLU78sUp/mWc/jbg1pFuF2
amC8lum5OQoV9pf+lE7Pv9TuZt2gV0GywyoluyjRNQJlv+E+npYtqdN5EXnE7dn9
zKzVat3OGDJ+2RsXUTPrpONOQe4AA9Jk2N7pfrGDEwfGeGDamBjndG9FAgNLCgbx
2BV+6ufowN0O3ZQupAVnVlKiLbKHThI6o8kvg9IMO42xImuKblLf890DdU3m9Dqo
zdh07R537O5QKDWHuh9+kwIYalefY8Re6gPtLGf2CzXATNrashUtlGaeuPy4Gczw
9kOVOngSt293NFdqCV1q4vYCYCBNpY+SnUvvMQzc1/dqcSvlpTfrbMbBoSqRvEC0
/tdqZkblny0DahTYb/7FU2VU7vbt8s7HvhWpoQ+A2XJV1PJVuuXNW2jfKaLunE8y
Kv4uaVgHxas9tN3Y6xpwI57MIYBDRd30uuIPYyVAS/qZkKXjx7zcEu5y4Q5GkezU
UG80+tbRA/g2r2mNiKtpBliDo28aD3pw/KGFsCa05nkz/z9DuFrvkOjvIFn4cs8H
OU5sBx8H4wOm2v/nIw5HWppbsUV83fhniOIDUe42a9KzRhesASeMvFCd57OEoAxS
lcHtElhZD0K9iJoleMILijM66syOHyhdNHmjYf08eB4E1LCepjIynvnl0TnQhFU4
tnW522eCGk3XAfHKy5roN4HUI2SoXdDtimjSHpJkt74XjvKEFCMwso7r87b1pl/Y
z7IvAi/86PK+vlXBAswdoUqiKEBBm6bfmJdTW1we/NHxgaRsIt8pKSibXv0xrehk
mhGWS4uOCXjBwI344hcksp0iXrgOA5wB6+hC2mE3n0oc/5yj9QWJDhpWs3Ytpmt6
S1Zciy6ttQ087ybVZylvL5a2IxsegHDez2QG0mWosBEr0hPRI2u9rhX7VDQC15rz
jSrP/K2ffdb6XJPUy7umdn+U53+qfC+rQC28CRWrnMYG2u+LvQUC5nN/m1Aff7+f
Mp2j3PnRhM+6NK9Xaoc79LYpiyL5Y/NR0rXFXBc/p9UANxJoNWF2b/ySsiX3pA6a
VMI0j50crtDFuRMXexCsm516NVnFFmKKgmQztOnA7Xw4pTRC23wt5Ub40YQ0rvc7
ZKcRFlRdJuUNC6t914orTZSCGLYgE1JKsVNF/BoJ1DFMZ8UwIX60WO0WF/38AzrN
Mv/cS88zh8pOvzPX9fS1HyqhMNzvh5cd6MgFHJUCelP/cVoVxfxqaMb+stPCK3VG
MPt9xGItD7P04B0xzenCIlOi6aCejS8UGjcDySPR2knQssezY7Cjn/UsuUv3MAC2
L3aGZZrwohmsagLXLuUeoqiV3Olwwn/JM8JvXdkoMxJs1a56Xw1EtAU69e0+RNfS
bPUewSqLCzLPJ6woHre5PB1/8FNUBfN4iNXIkSQe7U2F3BcSRe9LSbgNk+TW7o8x
sQVqTbeh1J/e9vq6Q4Fg7xLFGl9lovcrc0J5Il/3dzfWA2cilNhO3CfIqCqXZyN/
KNQSLq0EkG7pjjzTJFpu0fiYAgY5roadw/YKSXhjcQcbDQJEeDHjMsd8tJDjfn6y
cKmo3/7BhlAnnScTYgTSZap28x7od70rDUeunfh79571RKmoMpsxGxO7FXfCnTm8
AsR/QyThU2Zo/4U/w9TrnPScKi0F8alj94ESzKIYUVvYfjcf1h0rot5zNwvEQT7T
L0SiUCLiKleG5shJdyl8Dww5t7XIwUJx4tV5qqGMl6C3pQ3uP81Gybni4dXrtlJW
ySqkX7B0mrrre4XLrqXX/SHJE9q3P8rlQ29BDEGnpIXCUSJx5fa18QUjGGngc0WZ
J8nMGS3PsxN8E+3BXvL+k4CWr6CN9aD22NZpoDp3kiuPTH4tawfdpIzu792SHorE
As89NH430nYik1CNKemeckwMf9JeDk5Rpdtv/KD3JyWcaW3KzZdF6IqVik3BPrCS
WA62lfuZ7ZqDlVErxLjlg7zmvP/dusi1i0pMdSbNtgwpcorhAtHhQd1omM4j7QKB
K9+aLkrz7/10OBMfom3RXbjiE+Zh4Ex6Ttv+TgX/MiQkDIIDJpDCB46p/t184y59
P+EjoWgiIQ67dmquz+basfkQn3bA2SWLAVLhfRFm1h5CWK5R93v/d2r7ybPwknZx
L9c49wzEnyHrledtDgo8g5AxWMpZaCusjrTlYgJc5Flfphdqdx0cX3U8tatjPmaa
9bAJVt77YMPdplHm1fF/rgi5XuPkp23kDHf4GyIsdxPcFIN04p43gOoiD1q+Q1kb
RJOkoERZigYsrFulhV50qBtmHnG1VaJUJrtFzKO6c8a+JVZMlJTkgg80HMb3W7pu
ceFDLa0tGXtrxTcsFJVjqiDdjw64K+hADHPEyrKvvR7/V5ggUwQMQ+oCAGayWVv/
0BhEzQ8OZqd2HX19WvGqZz4vNUGkyxk7kTFONJ1j6BwaJpJfZ9WZrnJ13qQwb4g8
1jwmkhF/nw9hlCYdD+oFCRegs1TvUCs2N1+0mNstPSrF6txy1i6EmCvEU39vcqCQ
cDvrD5ZHgJRJzNEC/b+s8s1gkIi5rqMNCC6SrmD83saXdhD3thVx5e+Tp9+6/LTA
PWfGQvanwFUxIvWFiz1VuQirVpNzeva92KxOgQhcqoXXOdkJf4HY5h9jDNeJI0T1
OtHbfI4cPw8L6mbdgwuqI9wDjf64qNQqzJWym6eFIAFE/twzm8rzLGMzP8C+dksd
qbtljFyV0u6MyJ3xsURRwWaj+e657ocalarKgbIgTZFG5wzmXTqBGMaOOQJnPJ2U
3OdT3HKvz1aF0saiPmPNE1HLhjrGvNUMQFcTWPG6m5mhngcRZ4wopVR/SE82vo1/
IHxnVzo0/YGJvTTe1+vQ+YpAoMK4/e8IFM70SaRC7A8q7uruD4iLnfMpgmhcUafj
AbZBDiRiPdj55Dn9Dr1hH1tH/IkMjo07mLQUWpObEF21cjnZcw/M+XCMWlN6t+J4
ZieqmWIYZFBLDuRnwBYa65eFLy14e/aBOkcIO6HKx31tJd2MtVEHHJiYw9ZHal+h
zkPRyCZjbqSA1m1bIfGb81kfEjLvOyIsDEh49xRrXJnllsSpfffj2F50QhIUAGpb
nwczWF0a6XdkEDJ5c4uUVAvBrgfl1nYnJZTDIKsEi75vEbGNe3Cv8fk7D3zhhMgx
JNSoFaDd2Dq26k8EPNvUkd98qhpsF6X5mguzCD3n5bzyMyq74Tdd9DRKGwOVRldp
cqWLWeNilPSGSN7v1rBgscDU6RyZ4ysotFTb9DpzowD6CbsrOqBsjDQ2kTEBa3hv
z7OCP679aD9v95t66a6D8QCP3DYazfXr/kYPONb25CTF+q4nnh7oaPLuvIGFWw1k
Or/cJbgTuUHfO2Jiz20zzRto3Lx9g5jeHOhM3Nk/YShc+2cYLiYZEL2xhBWljUCM
RpvieNqpI76YRcBqIXKSobHdhLGWJFsq4vY4eQFHBwSYEnSaixymR/wyGw9H6Cba
9E7452sqDJhplWRXd6ai1YHCUziZb9KlxBxWLF11GFpb/gv0VcfuGP9S7tQgl2yL
D8LVvO1tAqqeN1Et7MYXQqAlvF0axoMktoP/QFym22CeyAAteRQIQiwcDXOR1DaS
tQfnIE6bpjmsaxsuW4500mp4XXE+6XtCy1KuMZWZV0lLxbCsq9kMEVHgc7FjlkgW
s54+qD9lUo3HMtqas6aOtpqEIr0wtHMDCfNf2+HRgqQ0/O4e+pwonDkSNfqWFFNg
B6gt86yeMULJkw6dXQgohPDweA4iMqB9HLG/J7wumIZH88LJXcNtNWNPs9Fat8qF
mUTScVsHhROMoyoWbc35OVCybm0qd+DdprsvBs0iMCoavVuMQ0kTPaW83QfJTIo6
K/6sAUMS0iEPJsbi5j4hCw/4wB7hNCrxZjdVXDxxSichN9OraA7TFWVxulnoaFL5
f84HWNUwTvBwlu+fWyDjOWe/l67Ao5xO+JB4GsD1rlC3hN6q4AgKqxC1Sg6Og5CY
FPZsRIPjbB2VQ7lgk84/R99pZ/gxpo3Iu5OgQPwULkzpjfHRl29bM2mrhCRJuv5B
aXF0k4ClYY0XevoyL7ZsGK4Yz/RZwI+134xn38746R5/nhf/OLVmWMgp7fIYlBU8
lzgHtmdAg0gq9wyFY+mYNbMsymHJOq+hb9X3IFm76pgRW+OflFIl78196uTJQ3mP
rqLrZvX76uufE0k35aKFA9V2CxBs9YmV0R5NGah8hILZBexmL/UILLqOm1N8h7ql
kkPcZ2E7Jwgqw+ohvyPntSFZHJChgCf9vreKJKKPycCc0MpCHx3rWVyZqRZdHv5c
hW6/ZH2snDMsoEhxtSahBPHzov7gH2bejyudi/9vev0a+U5epGEg3GzWE3fzLxtB
3BMQtbPCvpQkdUR8aIeNUXN2ADm8ifStpr4VKjLav6bkSaKkKjHrvBqc+fmadSmu
u+n9NiTff/TVmFC5JhF8x/j7oCLzJN6lH0bEZl3uIMytw6GGpHEp5SBlSDDluCqB
sACrTa2sSK37ScVNPIldZbXGE3StHGljvOa/Ba3CsxCSJ/U1kXv9GQ1jWM5PsDMX
NQx7RF0s+i29eBmmozFshKfs0fnHLZeWV357i9q+YAFOZFfbsuJuNtvVGm18kx/t
rfWP0hALtCGZ57DlusZw0RSON3lBJIptHTGGiH3mqk/ik48EE5LBXRt88NCRpQb7
CiOV4tT46fi2qbIB8+ty6bxBiqoMKkK8iR85KXFnj+U0v98PbJRpGR8wmw3505iD
1KhBHxg6wzpfJL84p/u12eJomxuHYdOMPYc7fwv9pi91Jh+zLryYDwHy5Bt+Z/wQ
Ep7Sxo+7U8BBMgXK2GAp4G9nDrLQ2f7DZe0Fjf5eNO5pfkgS27OSr4T6l3cGHaxh
wenrV326eGP/ZVAFGVHXjBUiWRBnSfbrVbJt7H3DOH0ZicbWTPMfjAp/zL9Rlwzi
wCnB5SN82+vTGqYKpc1XfqiQZysM63XTP+tMMBPBGenOTGLEXuX9+6+KbBVCclEU
E9Jy541MFWpQeEb0fP/HKtT+EhTY9RA1ieSqH4B5zkjCQ0kdGoeKnu33pa4kEwUH
30/AWGlbP8j28NkvaieFTiBMX2nWSlRVYlk5fyWu+SUnTAyORE/ZC7h4LSy6BJ/n
w57pqdXFzOgBMNZzGHJ8+yU1cXfpX73v0RUmo2Gl/ay0Js+NMJYLXDX1MUzx9rL4
N8keI2lub2MHkxGn7BexBV7jBNWxDER5+Ck6wobDVV3OuOmy0rn05x5b/hJr8vrl
+y/xay0PLZgZ9JdNyhcrU7EvH+Jfv15rE3X5s5ilPMXEQPy3tGi85ZIPbvaHw7xT
/5VZUZUtczRZFMGfEW4Khpqp9ftKO5l0ixB9XhG71f6qHcLeblpBAji2dPH+TNIl
vfJXWLlWm9xUwAtGJpN8HkJ/03P1nTRokIZHMOyFCrVcSrjb3+OrphPlt9nUyktG
sgeuoFSoovvI+Rm2J32ki60Co/Bzjyypi2QyHDwcm1iaKkg4oHDVdyuI9bvYt8OL
xEJ/pqadCByPWjE8p9Th6Hkw76oEN8NVpSAMC8cs4Mgmit9GmH8Un8glPVFjySji
dliQpRfnbzjOHvTwhUNCsLXE9bJ+r9Mri/Z4rNW3qWNME1HBL43OGgqkwvFnTLX/
0r/JeW+/gVw+dN0GO71o8zWCPE1KClUkQEDyEgn+R8q0t+zYbYePt3CqycScj2Bn
aaDugjima2u7wHsD6+Nx2f6U+6VjxqP0xhhKEwZuwb7el1aBVfB814u8AxZwv6Bs
Z535Roa7otBMIIkPsqe1Ih5PeYEv43V0bpeGbG9yMMEZ66/eEGBkIDsd3KYjTC5/
DfsOIhokcT+cjBF5FD0mj7V8kr4s1k6cbLjUpXpTHWiEYr+X+ouAcKBsp9OAyh3/
LAq6gDjH6hTFXxRD5ubsWzuiqBNhh2i9P5CzQb8zVItrW0f3ksI5J4mk7KloIsl7
E9FifQG8vNjyvZBPo6iZ72TGnv3UWCp3Y1J5T0Apg15nhInFLu4ksFp2WOQNOZLt
JaF8wNaNTaFRcnjIod2YDDwqLULYkTYJqofCIaLz0FjlkbLFTiMxJarVbrHLfnsC
mqv1stm/adEjulNdbXbN6Fu2bWZO9V0zTY/Ut0cniQCllhd4tmW5W3UwcoeM3/kB
h8qNI+urk9K8SYvqHWD1PHA1fduSX1Gq2NBacRTOjlJO4WhRWYhvjOB6e2hnON4/
Jd355M3HEyDJMmZWIteib9Q36LjgnGCZFxorzLxEYy7hTpnnrjik4BcAxuOOXACg
G7w/xMpJLXzmU3dPM6/OmsvhieoeO1f22cOcMekGD6tNjXh5ufdDxvIueTDuchmI
eEIl/p2As8RL2oJvx1Y9di76WDDCI4L7aWn8f39SXWPdG5hJDmtMalCVAcXx7F0I
8uhowUkfPfxoXElT6C+j6G0pyd3yyMakYBEjPIRRv6tw91WNT46R9gcNbwhbmgGx
HQs4ju+wAols+HUCX+nKZRz4Q+fnAhL5rjCQpK0QnVtupHwgQRWfI21/R9edEQGO
mW5A9fWCHw+yXkON1KWIXWnKlnnMq7WRggVjfHTears284+9eg4xAIxT3NQ/4aMn
ClXWf+CNUgHCP+emaRYUfIusuHYeFd6ejsqSDhvFGqY6FoGUUBFxSWx6WvEpH/FI
YnUBQLNgiNvTG9O+Defi20CI7gw2R41J6fHpaQzYitVlA/1i1Kz8dZc0fKCQeE3P
WE/8SI1o5ZjjGRnIGsVwApcobSzkxESaQLfl+Gp8NOZDLOr9+nMHskRo2Mt4WGhP
YpH8gQ0dhMOm/ANTtShKfrPKbP0NS8EuvAJjhPIIc+pjlAzLBUgGsvJFo+7To6Br
xNqCXIuOXL/6MisH+/zFuEQL1gPfiZ9peqGhP3PZwmN3UFbUW6kgdYtD7CB+lpVc
1Onwsea3paLITorAK0zN3ZYM899EIDKfAB/X2AsOhUpW4hwgXBYrJDeUPnVfWl6T
eOfaaNCszekH8fIGXLYrOrUTOd+T9zTNkrZ6ouIxOcj7+jix7OQuLh3eKTxsTbRq
HzrK49ejUiadEeVWeDIw/80+0lV2l/dw1ckLtVwOm73TqONYJBpAkn1OSxdtPpZF
eTIOuKWM+6SFmZgdcZYGvYcQ9qhAqcHQ5XvNA8B/bh51TOdDrFCzUzomXt6hJr46
pemDF97rUNwnvzUOnUer1tXeStPrd8VcOIaEB3fcDXGJueSpvEDYawW3sD/8zVz9
jFyQnglnPJzhZUZlLFo+m64yxZnbVrdi6+Gg2pFN/ozvaN+zKdYuIws82QGjWNeF
GosIxxTw9XvMmAI5SnQ9MVj5Vi/iKYgzBG0DpmXUoMQaAjZHjsKsaV0m3M2LWkgl
jGlsLu84+SDazGtWXWx+g1iLauXV9oDOhHWDm9FYjN/iChVWlQXEcMEWrqsVCWnC
cylUVy1vuiJp1ZH6+meMQ2uKtgg9RiFVak6ITDtI+bI2S9ARDealCws9/AuDW5Zq
bDPwkWQMyOos1NQ2HsOnEHj5KvSYBMtMCvOKgdUL2eFkeOUOm5Il9nP+sNov3W4W
xP+kN5jU2BFvgWjk3X+FG5OCihHVHrUJ9Q+myNrkbN3G6IZRBpeFFKYRWNVjemBU
nSuHvTpVDGod0oy/Bn+y1s8ytOzPZrd409OOm+8iqzYWIxlA90+B7pZNJA6p5HPY
j2a3kSfHN5PYeUN+nV6DQYxX+atEGuF4LpIRXNR5//ahQ/GJ+Hh5Xz8EZjzwbxBY
d09ds5+IRpATVXlQkRsqA+I+QbxODqkgF+WZbGGvnhpsiw2NybYSZ1bk3UMAOuw+
uKu1uM6SLWSPCa1ijjWQnzArCN+qo/+OmWf5aSlu9N9uqAPyhewedlPAaIVavVUJ
rvHHzIe1pxu/UgX3nGB6UR0VkPdEhE7KIInO5NRrFTJQtdeRDl547kjOb3tu0H8A
ef5PMjW6QZFh3MBa1sydxhg4QJdr6iUE7YTN7maNVhJk+BsDmpcdKIVdUq2NvIZS
4DkN1JB/mM6LXu6hvMBDZPFs1q0dRKPAJCWZnRJ3WTeHdNqs/UqsSqpYEFEnbyre
mB0JLoqnJJOxQ2OA5L6EYU8vwtK7qi9GmCDjXEhXBuP6joJ8lq6tbmIGFyDplKbq
2AGPWaDh1c/JW1M4RosXfuQfKFrYTFzgoTMXLMB28IxyrORGrjAbbISMC/R9xTSe
QfE5aSbdZVIdpKGBINk+qtpY/fTQm0axkPj8kWOgbOZfPfb9FLOhcd6e9MK68u/h
k3xiyeT2buDIQB/FaUSv2J270iIXTDWwPaAYrUvAkOw35Fw3df6MKwgOxKmgWke0
tl44eOlePjuucYsRxWwN204MY3/kd4ChhR28MtCIWQ0lwz0NA4cWr7yFfVZUL0FI
r03DKSqlhDfTpxguoOEj5HFxFFY3MQHWi1Ry9xc7LzI05Vf53EsMTNTW6MF0YyLU
b/LGjuCdvSzPHPpKMNwaYC/zKge8fQGAZQ8toaeCqrWCZEDpC4lDeuxEKoi8AXI9
KvpUy4HZ/+/e/M8OIuO5Tru7Di+4DmMMLc1GIMtK4Wndj3qgij2cnBNo6hqn0R5x
ySDMkUbn9t2zhMZXi9oP3G9RWFFROdYIgRYYLfesdlL/hRyjLQOnxGVC//nMWUma
OtYvCEb20+/az/hy4UoVImdHy+YfXUMX8XV0XzvwuipUYJYn9Xa2NkNEGj5/zpEv
97NFFjc2Dnmqk3UdAMfSlxr4/Er1GmDMmtib+LqFC9njnkfvHbt14/htsNVLDy9q
sGgscvovpB44yIfUYzES1ATWmFSB7Q+KT2lFLPdf3B10mlupS9HF1vD+bhPxwJKy
0e7qioTS3aGdxQEvLhA2I1YVtxynGPY3lrWDP8azcCBwA+ut6lDd7+FtUoLo6uuI
nGvp7nNSnnRBxhpS2p7cXMSA6dBvj3QlVsmrZLMPvQ7xDc3IoUGcIjlnuLTlGiDM
OM66KDVImuKnSNlMkYOQpf2WpUOaSMtMzETfg/iaQCIk5vb2DuUH0FZrvnJFf9W3
I9TOTRH86/y9+ldDbU9skPYLqS2LJfFqiS5hiuRWjl39FWO61aTxRrc++rD14vkj
gcZf9KOTpwwu0uEVQQw2TnP0plxIK8gX1XXeNI4CkULpV7Kvw2YwFXCfD2ipjluI
GECNV9hgSai6jlWfdeERQZs2Pb9C4udpqvtsN0+ByQlPsGZ+467JuJwrWiaHy5SL
4QHssHCuITo+cN4EO01W77hJLiS2c1bQX3opmzjflUz4ZrklDZGKeXjzKnz3bavk
FOwKRnn0uEH8D1jcLMtidEKqW50UZwk30ah1b72j3dQcranKtfg0ZEFOEG2KUA+S
w42ai0efglWPPkwM2UDGeZzQpZfPWMqi0D31UoDKUkKc9lzT1FyeswDpf0vzl+Hk
pEs8EIKNTLQL4Orj0lkzqPBY4yDJMMrqfIxir7tMDGQS1TUItS4QlnF8GdtqxBoI
Ktc8ZSwq0zbCo55sTA0FNOvt2xvSsQlYNa5PEMr1ofdRCiZjRfgmShxur60VRKM+
rSgYOLaMyN0jhSlErXhPitpbiF2JF3FW2wey/0BwrRf7xMlCGofYPJUQEKe10h7p
zH6rhFxzHS7N8FxBY3wzbYDG6kZVa3Qd8lAX0SUoE7EOWw8oALsCiZFOJKPZUost
8M1bMvuHeSM5/XsbDBJ9PK6+uKxupPDKyo6zYyCqUP0Et2KKvzeEyWaRl/42feMr
taUUcjlnhDVrrgx4QmzFxpKraIqtqUje4pBLkjQin3pvbmU+qgoftBcrdT+KqvMj
57JfSe8inbG10GNATM4Uw9UQluz0QzQ6QhWFP+bPhIuvDmPnU1vTEsJ6JLrAxUxF
PAKjrMvM2IQ3F+WOu5/EP6cFEJX+UvD9+mMWq/k/xOEtCXm38FMSu2ABwHi8H1UL
naDpFTMif0BgWlZ8qfMBtBhpC+7I9qGBjjwy4dnJxFC1Ca9EV9byyKhn+IFrMBoZ
YG7qmw2/6KLddu69fYUcI5zJYRez+E9an5iSIO5nTLfeN/yESYBcgxKRT5UQSJFU
a4bmqjzNNn6rKTZ1w58xsbrcYmMo9rbP8WaI2GglGgnVapYY42YgRDIoFDVJint4
CmiGSKu0vE9StfMZnG8mPuqsWyO11DBvS/54hO78DMVPt+7yyP+7PmHSz+l57Wf9
EBV1TvXL0xDk1fqutX7qNInOmsGZh5yZIW+lg5+FTJCSk1GzL4o7GhX6PuBO02pN
+wPoVJ6Cb9IQ+hvmgVef4FhfBl4mHfpvMyQOclLvnYHZE0Zh8NWgnz6ld7gc9gJ4
Y/KV+7OyCqJpelvgV5g73y7vxrSUoc8Njpfh1kD2WSoCstw5YpYN788pMzkloyIy
UYQ03WBXpKf/3CpMyuXZR5JWmdj0BdOk7D5bW/U2mupdmGWKVORotIX5y/+7CxPm
WsGRuHA9G59h5Ggx1EQbyoq2It/mXCaqryzbg81j+uZOzJfAJ1Wr3fusnZXSmwvb
Tj9X1DXlaqFh2WXn0X5UREpBcJoHDRTr3hEIeG+1VmNwhRDBf+D4AAhPlO95AzsG
j+XNzoHPdI6xHF6487XJWWHBiLsC26DZG57cBbficHI5Bsx13+yyhycZKqKsl7J+
haeV9yXFB4X0YHtreRgKypQAL3Vw3PLsGJk8tqljm2gYSu9fPhx5SCdFbKGA6Q56
7tSXQTSy/ny6XbpdW2xfD7eOTh44oELrmtwgQ7Y5eluobInLpAB+bSouFQLRPtW5
Z2W8Wed2f0+6N9KZJByC+7x8XlE1FRwqoSP6n6+NU6E1CUT6y0uPIJnSqEZ+Mc3k
pruwk7fQ2DR05mm9WFIrYK2THj5zfhnkyb2YBx7WoRtpsCkmeUNoGlvQTPAZYavd
kbZf2/aqmSySXvaiKPF5axx8L4v82ZZUDQjvGkogUZXk4zL0nv1pbY4sC7RooH75
LNlPXtrV8mOaGuvgn3dYr62R2rk85b46DXQL/PPpmChsvE/7tI7MZLkUj+7v3S9T
kkxPnPOS9djI+tcANRMrTy8trs4JW8FCHI49DhwXPxUFBgckJwSbPwfnOCxihxSq
KxXkEPSP83cTiKgA+tvSMr/+BkCmtyCJ+GlvJj/2Vf59ZoSKPOeQd9osT+orViEB
J+rARpSB76LfN/siWLKif7mSVBih1yM1Lx5cHbe+5CLxMTbN/O8H2UrarK4WlYPE
oQseGhCzgfjdLml5yKx8haZj2nn1+RlsWiqZI1H6F8ZMxCx1TJF5gSJAnq18Vqrj
GdvY93UF+pcHtVBT0UuU0Vjea5dx4dYWYaNCbsYRiFXzNRvAd7SkwiEdHS0/LUxS
iXOU00ASEgUDiQmQQE+B4sn92gJKQdFcFeKQee1uVttRkLOmyQGCbCnqBrKoOTFW
if0zl4UZksNByCgKpVr3smoYiQCIr+g5qE/5OAD5D2aX/l1NII+0uzl7OtOHEJRL
iwPvytSGHvIwgMHYap/xPJX7A/rVOnrWaa5tiefwO+6kd7GR2/e3IQZFqPjvy9DA
aM58dRijrdrpvezls0Hqp3k8qE9VsxJMvOF/zDfj79uqKZ7tBodl8ku7zLC2z3/6
AobOs/HEVXUb7XKiMESlyt1d/fDJcxjFWGLMzM85rBSK/+NyNZLbEWh9YcgYhq27
8r3RkayYmLYqVwNnFg+q4RmKdK6NWx2HjF9+QE1ranliJgNkw10ZyPT6q14ULTpj
mlYIse7z8GtAydWple8vdiAx8gJsiJuLX2rWOTQ30W8m0a2Zgh41qlFrUtBHaw5y
U+avfcowN7DDL/uPQQ2PFCh9g29jF2/IjK7weZ1jPU46Wy+GdVKUewrDCsm2nDi1
bqTyK3KxUtnedb5e3k9tp9meLIbbeJ9roxhBCnYpaT/pP0GgU18kRG2zL1FiTh0n
kXcPpXgFDAb0x9KmvXqKk3Sw2Y7F1Ki5909xOdwq2GvQY+akVo82u4ZJQaUxv4z8
8zZfnjC/QjztqIEig0sZRt+2yDx6akbxJ6hRu8R1ahR81eRlXZXHx6rVtq9wDBvL
0bZRaGM5RdvzSFiwGCYCk8edaRWfOQAEWpjVvHd3y1+p0sKt5T7Tp/84DdO/NYoz
QZ5dbylj7paDoRW5PAdKh3dFDRKdga13TBb8VYDrBjF4rS1dNzFUL3ko39MRLPli
90lI6VgdQ0+Zr5QELGIz7gAZCB/rr+WMrmOEQckcRzfUPnabMuJ+k3EXATCh1DCd
CudZcp9ZRrAI+U6FwcjyVSxmLHZH3GLtS9/KaN9XHtyDG/aC8aR3GA2JpNUh6WDe
yYxulA6RhvQOjmA0cbODvqYA0mzDNPUz7K9dJzLRNVHx0Vy/NwHJjzj6D9v3q1Hy
I7qo5zxjItMBetSrwb+SpsMiXasYiECzBtRmcTMBPh8338qFXY/U6ujKsxOKJqrg
mc5pyw80WIoNLNbqKasAu3dhd1AMSPyq8IgKsVOoB9Z2xvgjv8YXz29pEuqb/Qnh
Uh683qu0C9GLejYlk+wtD9rgfEr0u5GbaN5okG5BqQzVW8RAv+ssoRC154+IOzKe
0Vmb3tb9A04mdNYuKflxfy5459bHmHPpZMNBonDtcBliy1PcSLgbOS/hX4o14Ym8
OkiCJFwwtD1RDVQ4tkxXmSfd3j+GjcR4HLQIGsKLTNn8yOBkXQRT72YSLreFsX6g
4DX1lhKzyY8sn0UyXYSNOHYryvJKsj57nYB7NFSVtDLtUrItR5fy95q/kI4o7DQL
WKvo9LsoINtF2aTDZDwmOBzc8z3peQ4Yy6EsdRs/rGBlHVXgkLTrIqv0AAE6gQVj
TdKo55TvxS09x0ADzRDhpx2pDNN38moYud6Opl/xHN4ZjDweWA7VVeIxrtq6LQPV
rFFRXLuI4/wYae48s6s5GKcxFU4Y/2pKizZ8cLJ6S0rRXzISrJiEm0kp+3tXBcEq
wlXxscLHU+WE3WTfDU+JEl2xfpWx4bMpQ/0B3CG9SbcBeQnTuAr3S7CTbAWF2/Lz
iawDjbCjuXHxVNj+5h5gx5Cz8DnBuQNBIWYyJayoOpNqoYwHBGrT+ISQX5mW5etw
e+H9KTbSB3B4hF7t5o+NUDkP6R68Cvte88+Zl+I6Ipw9IMP7818+/A6J4uQ8RVaD
BjRknNVRB0sykN6b+m8JLnWLm9jqh2ANVEsMOgXdKhc3RW1Zu15sk4PyNrCzIlQf
W7W4itzhrvjsbNl/XP7/OP+E5kzJjmmyYEaXrNbJZXSi8eS334e9Mb4oZBpyBYBy
ORINgoHgsjIsfcXQLnsjENh963l78/dKQE4gKahAtvnn/ngjtI6R9ewH+RQ5n6RP
FyUTv7f+Shv8xxuCKouUVmQyDkaj+vSB0JVQE2W9VBGgk22CzzQgec6IAO/dJWh+
ioWK3NAA/MaL7N+oeacEcKoY2FOW7dPS87LYe9lUhYbvCLAbmmv0Blp0itbevorW
ObkJykNNyC7wZle0XQm6JlHdRZmCiti8BUuLZj2QjGvIpzruz0JRP51ovSFDv6li
jPzhmL3ONEgvmFdzz5ipv8GyHQPsEthkXZ8/5ppMEbHx9Xz20Td1OQAwmvBmmPBY
vlMlAdw3PLMVA/Lt1485FOHf2R5vmMXjBvorTQ4eUhCGwvpXKixbav0wCH8kb2l1
D5ncVJ1RbmOiAaCq1uO+aOPF0zssEN8QAiO+Fxek81YrUzYlGLwLripMscq2zk84
87mFKOyg5jCemZzMbizAmui0iOPVzD+zcfp3xD0j2vFkBoPkinSqvIT5HNwbTra1
N6amEc+4z1A6nmXAiSdLcAnTzLl5pvfzfGnwtg1omLIYJGO6N8w3OrfX426daKa8
sGz03AbAGV84xBn/L1z+n3T/gnhpF7qzg+wWSOHvEtN1fiMTQOwNZyPeAxJl3ooh
mnQmUfDxRCalxWVFwpM9NXE7HF6wt9PNwNjrgRs8oDUzAejO6VBzmyADUKlNJtbj
v8Wxalj0VUlvgN1mhIznFgEu85/sMSAURiMl0MYdMSQWp0CbQOnDGZ/9szhR8SiC
eCp75S25vUhZFUfOf22Am9O9/Ste9PVIJmiMg4HzX9hMv+8OYa8vc3DKi0L6x4QZ
ZU+BTMLiNhqyz+tfAOKEXkL/PJvSzhNU8WVJkQk/KUMhLiTYE6prjKlLzx733JaC
T7SJ8ZPIryzQvQ98vEmjtYlwz66N8tiG5bB5A4NHIxZB2UMGrLVThtOSWwkqw3Sv
7RLcrsWqLZfgaOh//76dnO2qLw6gwhTfvYdRzGRhpizryg+s2mf+e8iDYxzb0wvD
6vg4h16JTsjLdq6Mc85yIM6I0/RVTM+wajXHCUYs8iMdaFtfbwNFurkScYF51AvK
Aq/ElLWHw3h6W/X/eyI7KPWa32iIM0KIRu4gYuxz3rI/rOSSH/yk1GiOggDhciQs
Po6eHWJYwp7Wh3+qRfRJgBGN3FiljbVVDMSFEZiDdCSlWCE5E362kx9Evs8FEI41
+QTzhXepMYqUGaENo1M2SsJ5iwxJrL9+AYgA187UQO0lgxKyxWv/aoTCVMpwvMz+
j94erltVpsFF7YuxuNP69mbt8qfriLOrjgtFSOic4GFyLt6OJVNlgXwYc3l+6jA9
1eGLM903sNcvZkti7opT5WYJp9Z053rJfsdsIQXrtVotgJOBcxOki+IzqK132JE2
x8wFSukeluhjJUYX0oby6JXfy+SVPyYLHaoXsoGcmAzxNREdGUZXjxIsaWLvE63q
LchtGcAdM35Bnwo1wBAPYPDIfpMmg8ysaxGRejEbCfok3k9JV5Vy2I8GgvPvleLa
vxo/j/t1feWLtB8JD2PinSQ7jLgaigGGspPpwiQYKWBtrAd3VQc9PuV78D4LbMUK
+kZYfXQJ7le3ytohO9wTIKDtA6881krfd+Jp7mjk41oDfbn3zi/gTC0tVb03emYL
anBje61nU1e7lR8En4OhBPix74Ib8TujI57YzljHnq2RDCEtmk4kuGXRyozIlhWD
9BpUS2Fn8PJsCZ6s5EuHNFsGsp7GkEzKWWY9TS6wAn4t/7AkVjVyes+hn1E3VKof
EwlgAFvAtf4ysSppbdifhmxnSNc3XCto0exxxUDcvFORDriONVhK0M54nSunM5st
GjjkI2I+JJPO79XkmDCPOlSTvzQIiq3cfozBRbPq9hwWQ0rN2yj1fcDnBAcB2MVj
RNFOZrTxYDAX1i/1HTp/BssdCI5lwHEUUzY8ewq1ht5drw9YpTybYci9+QyW39hx
W5UeFReT/80Y5IGt7Uff/JEsDdD+PkJ2WqmHGRQWQSOxrpRUMXLPk4MCiH1vR5L2
P4KEmxQl1dZGlqhBitqBtEe6ZaKzCQobHrLB2cJeVsRHtSJBPM9IB+ZD/7B3cfeW
RLrCMLSYi36xLCflmtM5ieU8HYzQH/rUdGZEO2vqVrJr5wBov5/pF+iRCuIcyXrf
LPTah8Nages85ebx1EbcDOmS7TH5N0POQZxvP3bI85hMXov+671oEDkUoFtcyoHh
UXWGHJbUlWNnePo3Di6jS1/LFrRRcCGkTzmnr8TuSygi4ujSDFZ3QPTd5HlMAbYQ
j5aDjPF0yLGUbMCs9qhmtaygGcpfqA0ZgFMz+e6CGA3RC0yLztvN/yytxPSJ3QUO
2CkpBLF6LhJvJxEcSIjOvC396ku5iZST/oo5HK0bdR8S+Z3vjJcRHhxJIvOQLZNf
iOt958w32P/KxuNLEA44uEcCsQISfEc3BlqBV/ZYe4O882ACtezy9/Hmbb1QBc0N
1mCrS/FVs+1ElQtiqdKI2r3s27vBi0jsMVoa/4Zf7EXFElo7li/v4mDiz5BLjTw1
qAXVkJncfuy6xIusHWvMn5Crw/nsHfblDXy4iZ2qZO/GT+cuM2l1qGfboA1wnb+S
CGc+JFJBCJdu/2IJ/CSAu2Fo4gaFVleNzBUnfOEItaU0Tu3i8gslo+t+0d/qKTsM
clWHXpfzklKmf6m2SOt6jBmvnP2pHnhCJEjEv/em8Df7u+eUcyKmP4eRScsWBHyn
i58zMpXd+tIyu0wMwDFivLLa0w/qlvf0glPOFkS9/5JIsGN2Pu6/VyNTXV+GY73T
+d+I7sdpD67EqlHxODY2HsjNo+ItX8JQHOD8lHPnPtdU2e7SHtc3tz0mb7fyeHTM
os2GS09ggxe1zsE8hjUR8KdiwurvaNbS18O4qdgcEvNsmhnfXQs+9lzG9LKa0EY6
xemN4slQSaERXgrD3HCiOXI1odMB3m8Wq/QBsmOzR+ISzaS8mga/aU8ZMiQNTfYO
9Ql6BMiEtPpDwYG2qEcSWcAf35K0H5XjnqjUlabATAduGdYw3ciwSUM8pFL5GyYm
5J6AWUp62YLlg4na0yz9yHMd+3P0OkP6U4Ys5hJpIzGa8QoPmR9S8Ih6HzO5L9zC
AveOCzlR/TOn3CjHXKRjWU8ynMM61SccoKd+BtZCT5tyC6mtah0rEUtJvY0uNqTu
F42hxN+E3FLJg3KLyAKK0LKH8MH2HycPYKLUfFSg1UZ9BQQYJuUjHg847WQcdy8W
NQesFThxYA7jJ0WDbf8Ljxz3JsQ9GpoqEpIDcXIFMhDTUhJXhdo/rYZwkLrLdHXw
o6/30CLkHtDNpBn5+GQm3+up7+RJCbJo6Q05QWS4BfKEK111U7Js/ABQbWf6wvku
m5wg3SjXz+c+yvDt2gIViGHhTTpIkcQ1jjRwoRZSp9oGio3WjLzpZVsqizYdeZWv
pS5iZHbTFAK3Qa30uMHVfHac41XisiKjywRpFg85+04ZwHDVHSe7slvk7Ju0T3Gf
oeAYz/BlV69522WPmJb89Aq0Mzk4zjOfrkuuFOqAg3xE7CmgiKQLQzUw9IYXx6HH
lBr4NQ1JvhgoIT9Ijz5/lIyZpwE9AunfHHgm6kOtF9K8YAAslESTEgiWL63xhtSJ
56Q8wqZaQhQ1rdhIEsmsjzpgcbaBzWvgux5EpXJODcMOZKI89LtJ0uPhz1oNkGR0
lxC3VwWKI/KMtHcDuV48FxZ5y4lD+zh9dRbLmOIdy7nYHhyfqOXBrmj8n50PNHhm
NofnsDEr2PSTA6WS4sfAU/uuql3PChO4QeI3gvNoN2xMRacxTqESgF6o2QFwrNVx
8Gv/AmHYtsPmF9EeKT+5W574IjPHLkUbEKB7ODjPGoluuJaGFjLYcDh8Xc/cy1tB
9FoW8UO1NKIR4ORntiBiPH9p6bmZzimC10h3md7CXUiDs0BqSjTv+GuukHmRR3Yk
F2a4FoT8VLzkYYvbazOjymYrFwT4VCoVaw0jOtAm3TS3/A6YL1nuKpKEAisSQ/wE
MIJmBmA41X5+TbjUikNdQXtUJZ6vjLLXoaOuxenV9MwkNy+uFr7isks6qozT6MoY
Y2ArHIZuUug0MPbaUWvTdrtexO8mFNF+unsgnkpzKmvvxMtDbtyThYdl0WOhAsIK
Rhe09zhOG6mYKlGD5Hqau78/YgLiHU+UKxcRQU4KeU/6gvA8Usxcznwqtir4EG04
3bY1GdRbW/CuIY06MQkz/sdrjvgb/YOIi8V/RwPF29nAampJ0ypCwgYEqbpyk5H9
WcvbVGfXyCWnfaabFGMb80SPvh/dDO0ErKhHjLuXHDP2uvJooRUZmwCEM2wFjRiY
ucfzeKj1tJERWM8QjR1fDU2mh8ko1Btsef82tHoKawTenkoxwD5tURIps84Oinp1
PZnJDt7UEECyFxqo31ksgMIn0OUcPDIa2WgGqH23MfZlMYm95N100WeZ337osIlg
L4Bkjpys9nU2fk0NriNtP7Igmdj3ZKVwnoHbyQ+VAaCrleoozVnZsjG0eDUOvBNh
dT7EnfQdbyxjrzCYfAvsYhslqxOgxkEx0Raya+Sd5OwPnuQ+vHzTr3cYkSrrQ2Lu
2RuX9DMKKtJQ8salQLuOPQDj7DGerSIXvQ55WyyJaR+zyZ47JSopGd0Mzgn4H8+l
nJ+dUoJQm5HkVgXuEgNInhQioiBMFEadeZ+jisQl1A4/A4/IvOgysQPZwC1+N417
/l8MHjIn1qb3DBTLPFhgEbjtAgus87Ow/XTyjs3QnhFjigBrR+JIZqmr4s91Mo8M
8Z8KWmOWGbRee76pTzctbAct9odCPjBUCZt5N+AvtTgMxTg1m2/tlfUoe1kBqnsf
MjcJJ8HWTCrkoJMoXXhmrksHLP3w+RsKI5K7KonLCFPdg6BCbQsyv5R0E49yOfrn
BP3YSk+07neXj0Sd7UQAqTms3ozcSmNEWlhT6U13W4vAAqRAECfnvBRz3pQImoIB
kp5al2KKHWxX7SzhFI1gpPyvvJdHFxf+XSygJ76PVvnV46fiK80aEEDuj9M1PIxM
Cla2dW0IaUTW4OwnQuC90oI009EDXOAXr3gDKjcvQFW1lpdgSnPIu12CPPBxvREN
PHnZiPIOupUBtoCLpVwiN1CneO1j1wtat+0vs31n6hqLC8Y+WK40nZly9YvURa8E
IVzpCWylaRwubiWkQ/kaYxfUS9Z447/9mj65WqRd7Vg7Pn5eCod0ZNrKg+km+8fg
YHKD2IlPx4iR/P/b2CVtQRkytqVzV9CXXSVvT4stGjFqk1LVRSf2r7Bw0OVLwfF0
p9YnOgOUVtLhggyeTeHWlJndD+4sjJFzTRRZOzqQt39Ja89nUSsaeV/MJhs5guIF
0OFMjAGlTRF/HkYSVueper/dbo/tFa5GRJi3wF366vvzNUmVVmwZla4zl7hMFoI+
VS1tPCKzAbdEyHo0ID74g57yhwfYlNyEYlFjji2NJVR1MAM3r0dRC9EJTt1VxceB
8t+AeRvcQJ16NMnYtTQUo3SkrfC/zzajKLBSjLthVLpsZw2NoDNNCH/yCbmnGhWM
rAAGZGxEqfCr65sXXSrt0kOJYpSzyAWiVnT7AlVPWuShgPZ813dyT2wAG/0s8ta9
lPSWynjs83y7/L22lIKz5LobS+mSLD23oOHBQedw13C6NWfEm6NK9FkuQ6TtHt1H
bfbVh/rNqhZv2HkW/1azc9nlohMswFkf++nj11Gm1RUGEg3+vHAcZNss2h+oxoYj
RkHGeDMyuPvuC4Jo6iuqeVhEfm0aWUWTph3tDdzg5vb7jRJoHOdbvxb+pkbCUENH
f9BARfdeg8DO3wbkE9fp35VnX/sSGagOQ5YpSA3zqVANVvgHa1efQrCxr6BoJUb9
WXnCETE3rdRtcPgpCTNvB7x40betQsFse6qu9CJbqMhjKcskf60tvRLkba8/zaVl
oMONSqr5OCOsZOAuCmn9zvgdaWWactx8StUDNERSLeWj+fhpQLPjkxztTT7r/D6q
ru+cDtpkQhU/P0ZdZYYtO/+E6FmqOy6rU5opLpkQzgugzxudr3KfYJFWGPKDLHSy
kwbeNgX1APMaN6Z9U44+2darCR95E++YTBniURXUCb02eAwbv2jBzLkOJ34BHhq/
/9pjXLgZwvW/KgJvPNm2stNvlG0+epT4FttQrQh8TVStiMhE8YNdMzPWVLSqjqRM
iOxA8SZUMjuG4XDCQtuHTSlsqJnUQSowpAaPV4XuDaE9DYukHjYRf3xzfSumFk22
ggjmkgkRN/t9XfyY/Z5f8yAHWrvoS37jKaVkz80TgZG74b6Yfipm7je1Bf1SWfDA
iuNqCZKCDruQeNrafquBJl0H/hI7DFzsE1UZkkSz5H2e+2ebtX8UxBlJAPHpljVc
Ah0iWC2xbmhoSg7QMAVnxa065M6lAYjEMnn/pH4n/Enq1p/ERUZMEJgfelA3DjWw
otmp5pdSskdHf2nlNivKcC1Zbe6CzIows2mZmDewo9fSHib2d1ZVOt4qy4iZD8uw
rtBd7wn/9xY4UwyCLs2dUUO1TCih5Tff4zQz6QTdCv53Dg5WtslWOoUfdwWT1SWj
AULLAziH7m36sUfmFXdPL7yZKKNcPAnG5AeK339XkfHfGmyUTLS5TLZEZsDHPcY8
0jvaCHAcF/Ij+dte3CuMnLKjGAFuL+6Y1PntkILEZuFNXwNT6aa6ayXKNKx1Ci2G
rHw440Qx/CdwuA+aqjpaCIXnVxj12onBQTADgT26gL85HL4bmhGAKzVyqMs6bbmk
FvcCPCHsN8EsZkZM1O0WVAoKPoRwE/vPa5kjprcAj34cXu7voSkfzNHLuwZ/5pWK
qavxi/Uj4HBYPqfnA1YcNWLYjIBNdzu3ZLaAhj/iy58XIbFhpNi5YTKG6DjxbNX1
yUlb7S+6TrFK0GrZpl1wEN96oEx+r3tGuirvffMUEE5p6KUrQPLFriJWWad9Dlz5
lTYoWCMy9E830tVgiL+FfryUBkS4Po9/c4O1D1ihQyux0CIZWBbtmAjqArfT3eiq
LT4kxrFtgTlDilQy3Vb3h7uk5Ua7scFeFduDy+xM8nY/hE6Gyx82IVmWWfG8p++y
hsuxmqMMlKvmGs9YxHxp1Bk3JBfDcptwenp7EuwFdLMc0IXya/QnEkrmPwiWZ4ps
JkvwddLC0hr7ZA2pAr/F0yeP7MioYeVULKDXfDQCHnayszKMv/cx2KQ4KNXz1bYv
NbNi5LCqGOs1MhpuuWYDWPA+xkVRtUkxrquEW6UkblQ9FcZozySQW+jB7MhCJ5pX
UYoj8yLLYJbEuoCHQpHfZY6OU8MqiMmfWAzi/V/pF86QaxDX53nkd1ZM9CrZP00O
9c7CYJy37GxIyHVRmVRe0ziJPHqY14DzXzYiyTbnjybEdDho6OKqqPJSKCyOGaPn
3sen7gz3yReziGYbA9wsulOj5b+/Ofm3mIdJaT7txbQe96auiapYW/0+ADqaTZBk
4MAfAAOceKKMavOz3aKskbK5do5ejjfLrAQDJ0Ra7rXP8VV8Tfqh92Q4J1TK3Z67
2bzKe+7sXCru0iXtMYN/v4lBom5W9nox6ry/vAB/OYGvTeUCSEGPnuBEvILhaEX8
gqdpVfIBDDBE3bcX/5/dX6f9gQZn9pqcwxuK4M+fZoW1Lq7vL3xmVvUG7nYGDUm8
YQHREtilo9XQDkHn+Q05hOAwzpPfHLzgQPXc6x0t/od7+u9ZYK4oGfzySuKBOA2b
TeA0enGy9GQ4gi25VmBS8J3WCU2b0dMjZN55AUqQEag0LkU8asuaMy81WYgVTVBE
B6FoFVDi7uCu47xOILDhS7Y9i4dJy6IO33KhiPbF4M/KiVFg5zqiURQtjhhtTtmh
Ui0K+x6t/oCB3FgJZwuj32QO0xPk8BklumaD6+QjQny3G99EQIWnRJTjDo3Vvpc1
GeKDHyupaCbeKAZUbsrwROOK5/bx6VLVh1HWt9TqS4GNI8P7y8GrgFUQtcLGZVJq
GjUzA/lFnUw59X4lXGhnsC5XLpR2DYi2KPaqbi6r8RsV2SI57R3V7bG9lqEIvu08
fTS5dwcStb/mHZ5MVRSoEjHwijJfgKHY20ia5Li0c6MUN9WD3qM0WBHQ7NOZV911
YreaQ5eDUUPyBL6XulDaoDdZYmASiZBHhNkASB5TDU3epsJp+bBGOUPKE5wz9iC9
UwiMKxy02Lls/p8XYMy/aqR2MK8pkAQhDAhq14JRrUyT0TAhNmZANTGkpm+acgVp
zrY7UfzgAKmoe0n7dzAWfLVuvd+EGvK/y+04eihS+WoZga+U6mLVAvDKvSlHscEP
u4FlcOd743zTz2yTpdBz3+f9i0QShX6mY2mFt9QqKn/4FRgJXlzwduw0+m31PLpO
f2v7wHruHduBxJS6mSOVGM8cdUNsnRp4UMGFbyg6pmdWZnC46Ww50uUyxqC92JvT
6y+swvLLsTMg6Ciw/+IYOSX7Jre0kBSM5dJOj0bCNOZOkDL96Gsfy7odJbOlwQ/9
vPMJEVlVZYH4CMZz5BN2IOsl8Hb/nsq5nPXI8leNQeHMevN9H83ikuTECmRiPj3m
pcxFGETXIyiFzprcgGBsAr61OaIXZwe4mwgpWfL5cPqe3LgyZFwDh1hHCV3HE6DB
c7n/Hum4L8gdQiLEz9ubJQb0Cq6+1MIkmkYbK6LbOw4awJZ6gZNmChDqwkMtJFrf
YYaMFlVwjrX//AwReiDJeLeOwe5icXSEcyxk3ErgFtchHU7RZzC9X7d/sR5gEQz9
n5fSlzbQqKoc8HR0c2VysvTOSoCcrUlnXn7X36e6ThrC2EYWfECodwaLgUEUrI1R
3Ra4PMnzQubdJdwJVobvr4EKudoMrRuiCmHJopO+5xpOaPqwgd9FLW8jUu9T5OW0
+BLP+fvUhF+dGkrj+k55zP1tJvU3DiCh60HpO243xzWsv4Yx6SS1eAICpoF8to/K
MFL2eGM59IJO7WkMdGZ0GSvTddcOErnpT3dCdR6ZZ30kqYq29Lss4l4dDkCgtIxd
sdFouZlXX6SEli6gkZK2bVFoQH39vyi+0pdDhwjqOebOSqvKWC7Z0/POuYbm3nQV
dlsfkzz9a4soLxIPV1EsbRUYpD/RC/Cg1Nxlhra0X+tjguLpP7YJkeqfRYulF4an
Kj6haMHKFTx3z/rXk8AFTXn+8vGYbybgU1mVlC7vSD3uafNFGu1DxBp5XR1om8qC
uVcs0KcEr55P5e/r/jR/oOpt6j7SiHFN+ZJ9gnopsFFuGx9qTzx6ihqPTyhPGbVI
s6Z8jm+Cy+MEUg6g4DWwIP419C0599USueWh1OmW7LykTsCpBwYRj+QF9nmNhpmN
+XnLoO1wahm/74q+YtWTrpVxlppkY4+sFUPrgMzeesiWlc1taT6YvUnhZnT2LhkE
OAkAFso0jlJ/nu/V8E/g2dW0T4bfP1QwTClBQrTJDVl1wgeMa4hIEjmkTK+EOUPj
ZSGOZCgzJFROhj/CiC3u6ENrxagIevuynHLcTb07PMEy4aa/lCdvOAK+av6G2eoZ
rKUOanCgWi3j0FUvHLoM1W5DUtl7z0LmAuAdhoXoxB858bfxzXB2qc/euxJewqOO
TOKL2J+a+cG1b87CPjKnXI/lUqAR8UH9HYo0XdxCD+0zMiUHjgTMNJy+0ZwvVHyC
GjOY2cYzyP3xDFlTCmHe/8kPN/FBiFi8rxcq/f9UNPLCjQ0vZsLFt5Y4I5pP9Vy7
rzQ+wC19gGwjwN0HyOjpcrOdcnQYfYNlHEvHNqvGV2Ys7KcNfezbrKJhXYTR+wtm
GJ0hVrGLyF1Zc/SwG5s9w4SRQvNAZ9/Kp/M0VvIBNHsZ95/B5ies6y1RvtW20QDl
Vb8mSsFuJhgv1Q0MN2PgEPZfdLhJ8ozfWo07DKov5gST7YNzKy0TEiW1ig4MpAo8
qWZsv97eSxNTcbkg9HDTMvaQqclXP/6WVbipqDtvTmnPoeYrYXfSpOUskLiCBRSX
sDOIYS4tp7YpU51k6btwOF7dHIffX94sO2h9E8vbhu3VAbmp7i+mJEHU89ySj1jc
piWFt65EXwKDFgzwEKBfn/Rp/Q6MvBFJE735VaKYMj3IybIKXh10O6e4R9uj1xrN
dN2iL7QnpT2Vd7thmRKUQULcpaHCiqNHu9HaJhanjKWgfQbo7+bFf1pFEFJpNll1
5yG7BAGLsLODWihBcmLO2r/zWsgBT3Lp4YN6lYWBzayAy3z9LXdgYfG7WNClR5XR
/h5/Avjh/apYy71n2PenrFcdd7/SjxpdVPXF0dMgySX5itM7VEPnjNtnqW8p51Ee
miLWoiB1YA8K/ifhtsTo1YoMfdvnhU5DqWn/Wj1aCa9yKL7+t58girb9TR6b1QqS
nERwBDn7icB8k/rQrD6nLLF+9sEwm/0/6gZOzS8gCDcEwjmgodgtUnkc7vhRDtUq
dEsANd27AB1HYkhwXZPrrNCWk+KU154Ok9Q7zKSNl2lECcLD8fsqmNeOEdKCi0rq
rEMrjrhQwGfUXo8ZI3xGKh+jp6ae/ENEJe8YILtznn4TrEUuVGVi6ULhPsnPdNaC
06yBLyOFUgVGK0pfL4mmEvgQ4c1+vajXQ2oayJwOJFkeXvI/OFStxq7mX0XNNdLp
qUqoWb7nGUelbitvJ82z1RmqEEGmYIvNpygb9Oco6j7XyAeY8DDfWRLG/01xHkcl
V1KIcsQhuei0s1lp3sbfmz/ywbaxoKiGgKoJ6WoScn74Yj/of/Ai1rOOtst+7yj8
UP7h1vawoU5EjQJcJ5e9YSA9GxzmjoRQ5RTW/KYL/IUXiQhhsbtQxgT36JCMDw8X
/lrkkQouWdHhzBb2i6qH5Osj8SaQo8DZnmR3zky8xqe6MTiR9g/1/yX3F6LNgku/
qvbbV7FR8QCBg/ZWCoMMKx93DMJ/IAuI4y+9vJgy6Q/uqf0GlSfAKZpyH5QcZcia
OkasHqn/Cf3ujei9tAtAllEGz6ui9AoqBUnW3nfRLHL6uWZyLjxnnUs7fwLLnwW6
8TrQJZ/09Hz+9NKsuIPuro8BAVUrx8zn0T5cG/GgUjf4dbprp41COkWGAc9aKcLV
vTx3BklEwvMfHJzWAUu/CbT6lQZRvzfxc6pUhEpdURqCdA1tDI/74IL1InDKHm6Y
Yv/WKnN06qUNb9KJEDiik2+IfQ6Nbyu+ox902Dbz2RRQ7Y/wftiVhatEa9EL3TLk
81NHnxFcFxPN91u8CMleP+ZQ0LKlw4zoENqW1nbaSRBx6FEO32SlveVRCVOdFaLU
exUHDcSPLSsrVR9icYRKp6gnAznVRxm4El0GDQYVLVaCBUdkHKlzSnkrNmspYNn/
DSRZ9Zbmrppfaw7P7yUNP8Ay9+wQthIoOH3W5tc2KY4EB798t3qw0B1EqxsXa+ov
igzEmffZtA6y5PuOq0DWmwN8uvjQ06n/+Jx1KmLLFKMGo7Y4dXSkH2HbNmvd86wu
vr3BYOS+82slMMTx5SI6kTGFcw6MyqoHOTNilI8I9/618odKuL/At5NjxaHi5fcz
eF91pX9S86niliniT12Qjl+EZvQ7l/ZEr4YtPu9+z1/BjDqeBg1Jj3KkPkqcYcf3
ZAJLqisvtQ6jIWSJw9xVOAph1D0Juq7098WotCMYUKTBGH4JcUGRIBGz+tMXNhZT
GjMGWnNf9USiAcnTsuI+5Ql21gV4uQ+AyNZaHc/UBG8w5r6bklrT0WiE/W50tKaS
UrEE2+6M89qwyavtTyZRg/atMkeLWn4Iat3RFzTtR7TUgAPbLJpjp+F4nNX0OTTU
5Vpmehv5qbacCDyLZ58abEcbAn0NfzJ7gCpoEtFayFKIxAWdKhHESZwuQHSHHTR+
C8/eDjh9BFmCvzJjS5k5rULm5z+sR5go7auRgC9rW0v5EwxkY9tKCHZAf0D4VrDk
gUB3HSt7m8XwpjarRx5L0b4TLl58V9rT1Bi6u7H+hOQ80pT8E9lq8JCiGvs49Yl9
Y0kWzwTyhDHZVD7jM2atVgSmOOtGHw/HO0UcOTJc0TPe4sWTdDvQm/cad37WdYna
Q5X7B9/Eu1IZvmD8S0r8VUhrGkh0/XzDgFfglKIqS49/sQLIVn32TmzFIROUdqDw
cmXQUrowo14KIQLsH3RdCq1MMT9iOp5JZi6/Zz0869mZjbOodbfRbFWBySnYjB4B
zlL6MqG1lSKKWy1nY/w2npYuiPd5D2v+JU0lNxa5oTfM6YNeVber1GEk3+/BxTq9
T6UEFDYOzgTW38EKT59UqASm+Xj5JfAgdn9Og+XjBIU1wxcYz8YgQ/yRFPdjvqtC
rJvJ9yP38ZpSF7G2/c+5GZ3G+MFOTpWE4JDVfsfEa12aGdCHz+Cwf38nkMMn2/v1
fcCqMgnru8vEN9bvcULDhM2BSuUjRC8+4sJSfaDhr6B0Fk0Mg0ZhQ+j5xKKOd9ry
HlaOX8AX7nR14GR1pr1lG1Teqh03eYTj2awZH8LZtu9dX09lUDJSXMqdpBEfd/TD
+vajQIX/g0PviE96sTWgZKpRBvL4Cc0PhGOUPr6o+uIZbwiKMspopN/CCU2goJFT
egjSyQYSVfJaFbZtSNTKu52aud6ofDY++TSpqmd0An1qi7nhgTrAb6dI0uRds/5m
Z+YgbO3LfJ2V+lbtWZn5NTMj/NwKW34kU9IWt6F101VF5aiB8gxWJsp6cDdgr3Tf
hcykS/GHG6nNhUdfv63yTZAvJc7jHb5RWHXihdaNwepF1EfF5b8cqva8TgNlctDP
6wzX0M3IawGvo6A4AZs0ONG8izSRTPjCTSCu3vBtBXFumfeHT5Hk9WHFYlm6alLs
qIcEB8YEnY/ebNjaQV4YdfZR5AC2yW4sOCWElqEtTgks9/WMUfyMBQ56g66hofyK
c3Ojc92p6oFa8nSyTEd4ip3PgUI3tCGTDysiHuqCE69X06Gci/DnW1RGlG6iQfPx
UVWQ5KH9qtoqSZ9zTYRAVsYW9TcxIBByTO2N2yF/+IlaNCUarNk0dC10r/sTeOHw
cgajRZyrJJ+InJwLx4BNMwZ5rPWE3QhWDJZtX77e/lFOGYogyKwzRevsmBLgZVf6
hqjE3Gnr4ki2VGxXhdCL8uNBY/mz8kGSSUswPn4sCVtkYPFwps29gcotLyMhWTHM
OnYCb+zctojFgVHtO5gBWyirysJNhan/yarvWtcwfBz9JnPS5wrVZ1M1XlsXpskM
d6VKDRnZfPP8OGbpF4oxThKJcEN/FUYioAjQIb5FI/m3NZcl5Svr7QH7rtmwgrew
u92eBCNA46TqCtC2eKfccmHyP6K2QqYAp7+/+770itVxRUC89cntIqoS3feCBUgS
gRP4FE+UTlgU53IwZNnQ4HSf0DPorFlSuJ05zSktfZOKdU0gUyDay5JSEogf1dTa
JNikfmnD9epxKos1r5pY4aqlvNOrgMKMexv1mo2Ssa++UQM8DDt1BJ1edC7F5DqZ
TI6B+9817Z1pA4/QKiXRODsMlN0+lEm/Jr/2YUY2Ocr2qvjOjiNS5UNNPEOTy+S1
HpI6m6r1+CHmjKuPDPa6HuaXplrSZTaKTTq6zv5oks+U+Pvx+fWTmz73V8qZDGAz
Fwke/fZaU99hGQHs1RaPm7GHZLsAeC4bhMkhF6tmruYDh9RN7rfObwpEXamcPx6x
wwvIDkMk7/r0EDxt31i+HMVrXJD3cpDB69yaVUTShxbCEd5VJ1f65ligefvnxPTu
pvLgwWuiPHGVzgnnzfcN5sfXMk6a7BAlaxbAaE71RJVy2tD7Kpl8+21WTqiGE+Nb
lharhU88dkEYFDhpyo/hEfWVQq9D6XAdlwOW1Uy+uffDg+4VeyGsoXKjCDU873p6
CZnEmijUkgaJHB6SbqUxx0egskyxuwPKOSAIc4dVYYygDLIul0Jrm17joSi271+h
VEJ6DD2uZRsM2Y5CEu3dfmJRcAOo/3U2AKGRdHBYJsZJhApZUw4Mj0t594ttdux4
R2MAxmj4KiyfNuQpQMRySFu5PATymWldNoI8lMuVtm6IxKNUNNvGpxM6zzy2Uio/
EtOvOa4Q8S01CsEmeT6dSqblQu5udL9ZcZ6YDjDuIJkFX8hh50r3zLnSgIPRO/Wm
PJviOxPjsFDhlO8E60ViGRouLapcJkBuYP9TP20YT+60JcBbU/4FhaLX3cyDbwgI
JF0GbZ1ZdW2XW/z0bTpZJPqyWP2o93YjSdTDPriW0IjqRALb07ZMghI1fHW1gzLG
LM/1JPmc2nBP8YiU5DecQ5D/GhwEbZjTRiD+hzygzfUz5p1RW0lpDH2MCfI6S2Dt
fducThWq/9IJsi1Jhj2DyJ97/nD04fg/S+Bnvmru9G8dUmLiez9mnQbvB+Ta5NTA
uFf1YDC6ARmKYb6vMAh9IsWWxgiDxFVIZiFNB+7aZTcB4tEhJBh2MGF1KpHLCAcS
OfklbACoCKKmoAFC718NXNGpyzibVUWCEGHYALwmI1BYDfm/typQCbyy6S3FQLny
LSrvbJ5TxT3S1H0ZP2PFPJMGvJz4nyTQjfWQvi9Xw+sHoiM3Y89AHOeKsrqVR1Bt
NtvbLOiB3nYILISsillyLZj+YoDHw8Vd1qGsDBqbx+ak4E9fUTdCmRJpX+f+n4Ew
OgzBjUEP1dL6EC33xGKYC0WlxUp3X6iDvm+wRZGSeRHUtwOVZY2mKtV1xoeAD5QK
WvW0pommbVtavwVZKrPdXgsMTBaCVQVBFa5ythzRQDmSMmT7mBd/S7COQuN+5t4t
ONHI92RZ/fd+95KBnCUkPdAPu6qR809/+cpxBB+spTbtzKYgESCnES1QD4Ai3X/Z
QCE9OMZ05I12fOg5AWDeCHOWtZNbf3YSWJFBOYLmKPaeyjSfYeQj79tWHVi96kE6
tmeNQ6ElRZ24jkhO2NzRNrD44mesmXSDizK07WBRaM77cm1xuvppVnYVv5DAQ6nZ
vZetEAbsKoQW33vaH+4pKy0A3O934ITFJGYuZyYKAVTtFyNJ+A2R6kPF5TZ5gg0P
UWKxALvhL/MlOrKT5xb9cOnMz7uL67NXDzEMcIwRYmKSwbap7GVkoaT0YwusP2po
BeWTyOSP/MjvCrxSoMVkLCESqDnqR6bU9nIFYszaUcNp8vxc+3Y7A3JcIX2g3s85
HC3VoISNcGar6aPE+9wm7EUdnWODSchhXhZNChmzrQJ116Ws5fokOEVHLFGxGTGi
mqIau/2myN+y/mRwo7klQvV04TAc8xp7oftZ0Ip9tfFy5Bz0OMrWrQBijM3ZKKUy
cw3UfQRj+uxj4o+o0s/HhGJqQXuNJ+UX/g5pKHvajF146hFXlITPXB81xWsJ+iRD
DbfSNQegSbX9sKUsXlKQx6uBcEpAbzRixV2maZqzIbcHoy+TlmBPifpnDQJrsUtJ
64uZb/vH3NQkt9KhVUUWK/q3PovozJX0+QTkgy63mJWE70d4uBLepMvpOl/2rEgW
8qyBuOrbvd8HcamD8HxnrauSd5Lq12GbavFaIcu80QRF83WBRWyU6KH6fJrM+JB8
tJPMw6SxW0T9ZllvmrT/mU2K5j2CZq6dSiD/WC+fg21B2haVM57mxI2W11jeRLp6
dO6tvmgY9DoU7rFs84CY5Hs2vPBCEHB9YbjAzkbZtfWmOUELDhaTU55uh3OvFlQe
M/PfHi3UMSCeLUlGrYhJs7fz70FuWhscrWTFcf6E0T5KZgeKhcd9WJi3219mku28
xZejv7euXs9oDbN6KQivU3xZGy66oMOdWFtTR5ObbR5IomXEnAiHJ61XolkfGWMO
pmpVb9eRFn/QEYD0SGRGYV2tHPe0DIWiIZHlX7yqHqZSlbMcdz9TyQk+uD7umA1r
0og3ABfcJKitj1KxzDIsSqEOYi48QLcIFdgJCfpITuEBdM6qv+OXIKZ7eSUrGUgJ
tbV1oEJQPDn6l21lACe76BRHsfZ2/eq6uJ28f84yl0uXidxrIeRuBISiOZTkzR1C
eMCsv2llji5O0przxy6IUR7xTxM3qMxnpPxYD0lilfw/bfAh03I+DYoWf591qyhx
rSJX6tsZewm9lzfoErf+L1qD2fbg8dYyd36+vmTtlCy3uyoU0J7DSaw/H+S3CKvG
2WDXzJFP+R1rUZ/qCLmLapwLuEHoT6bfljFYxGyYs9vungSrdmunqStg7TeLCC9b
viysdSvw74k2Z6ZDkfQf+954pFQIsLYw41b/X4I1DDhZEq8T+vWdB3cTCnT2rget
AAdaDDcabgg99qBilfemq0XBbFZOBKIpmAtuhScdWVX0G3ZYtg7D9AhcBHJ3gOMD
iDeGqnNsFK53kMuQ5m5bFLoFvpog/aSmaC92U4dDL3qKjC+IckPQ5z/u0PYOKElO
+XXNcfr5i++HGQYt0ou3mrKM2tMFG66tpVpTmiarElCHHG3zjI1CMVcTjBKDts5G
ZZT+01jVtFc3nPQu1/H5IgRq/o1KuOl6dO2hNFplEo/9CXQ4ostNduYUvatrZpv3
IuiQffBZe3ytw4/yJE4/qzKGAOfX9r6wRasOSjd5HpG6D8/93BECSHOnzlQiSAIJ
g14BY8hy1KfqVH00s93lYMMILCmq2d7xfCekW9F2YGfPUBvm9C5RGFJOgQfdcjgF
45d8nkOjnO7dLhPx25XJbO1yIUcd1vEm8jSblYuLJTBOY+1SCgBeDusHq0l2fPkM
As767kp3B1PlDtDSn7P9KdFOZuYN1Ifb/BlD5OgQ1BS7skfTge80O+v8N88JuTcD
IFwrHzIs4DyukTxlNZqzA+LUqcADsf3X8+Shic4YSENHlkDhslrfQTmVq8D8iH2Z
AHU9iO90Z2JiRAQyTDTH4dydVAfjYbO4QMC11u4pM2YF4EOp8H9+eCh4XEJpk26s
Ou0rCsycVahw/DgSxQyz8DUBjjVSBRBjmPdY4cGdwziMaGe4drdhCGIntBSeD1s6
2p1Wk/n1KWe52MYuQxClCR3t+IlOao9IATALnGfuJjzZ1bqv3j2vAsyUtRjxdc9v
ME9N1bdNz7hRu6AZ6mGMUue4/o7TBegF3G3Dbq8jHBFkLw6W5qZeyeAesmTiITcj
3vSfyrzmjlQSPn7IkdtASHt09RPwyW7qer9I8PSKzYtS4CroTzIBMQYq5pInz74F
7tHaZO4sawrA8v+ez429/WNPTFA8PNY90KNSfPiCgBQlRBNBcDR2u6uQPGTSP6fD
vHalVtYKtegqkPHDa0vRGe8wX6bBtMUsPXGXe/x3HsnOxhhp+LB4tOx3EOnUUhUm
uAFHzADV2tebBFomTL9X6p0BbX4D+0w3K/VHV5jPlESw4j+PedR1bJ+QbcNKOolM
EGTNZDZQj8HH1xWU3F+NzNjd3Uz0p4JdRU8oLTqQ6tLvHlEHp81YfwGeONmG7i+R
p7BezvyiD75LV86PjxdZIFfKkicETM4oU7wtSTZVt/Plrbs33MkRT9UbpAmEm3lB
1WjaB17DCvxIi9ZeP7gbsk+Hh/rSQQaUSdek4/Ln+PeDGV5uh4yHWGSS8A3wDfve
dBk46Sud5QajKNtsdOzbGugvEHjUPN0VVunwFMDRiCe7xVBy6DWYilnlxRHAqdxi
Etvux5q8l9fn6dRXjmEYAD8qqbMpPo3VCmKDP+VnJF1HQMXoIgvDZoNb5vfAO5fU
Ev7B1ScGOV4n9TIbPhvdC0eY4obA/8UwboZOXIkWWGk7/OsrWDIQMDUbsaCIlPQb
lWurJpuCwd5GysOzt19XoDPZaGFmZPCAmcfJ30vgl+M50U931ycB+qIuP0E3kVM7
IyWDYdrq+wmT/CQP6qGz4K17ZeDuMDoUh9/uDaol7dToEyYrxqOUXy/5Z+Xv64F1
InwrXoVIBRQIdf5EV7culPQb1jCBa3DNviHjrhdi6hYNzA/NDOGOCKmkI5MSgsgh
8xJIH/D9Jzxn5lPFU/DcybH85O70R/+bx5QvApnunJwDK1wgIPizRByVq4sWsQaR
RBmbc5OJ+RdO64aM2D0W+nPZ9DBA5eyCmdtfQqydvbUMUvj9DmqNZY/gAA49MjPr
N/Ykb5QwXlvilMq33QWwhDGTpi7avd3jWAkVyHhZX3ylDChkLbV0AUKP1Z0v00aH
JqvDM5niLzkHD2tLqd9LHFb7iG1DtQ3jI2dhGqpy8sVpiZJu2lpMJPNeWTW3SAj2
NZKSpQ76KxKSWCoMAJzfDPHVWM02U2EvcY2jpYKlDgHwnNnCJ80qBIVm2qRRcrpJ
TIkIiDFrDbSyW9fbPOlTQUh4ewIJbOYU7R/3c9YUku3BXfmy+qx8u3jkYkKPmXSV
TC7Tz0hSa/1dTa1MmCKj9y0+OaAOVP6AtbuOjKiJsCfHKTlkv4HjR7yBPSoht/Dk
LKFZAXeXrwAj+R7n2HnGpXtP18rvdtjSeEGhwDCDvSI8MwGZ+VP8cHgiVC8eCqXD
1C8inRErgPt1hNFU5i//EgklGYAdVrUCiASrmWSEId6KNFpvyhLviUTEZysBR0z1
miFis3r188zSLAJ8dULXDCrN9lRJbjE7HWGVadtMyAXOepY2ETq5hnEplAB0BLDY
O7qvoJqdgBJG6V2aWuN54/B7/bdLXZTIeN9PX35qtyKzGI8IqeeTEspGr3hC2K2g
3ivmtG4/H99SfTUXA1fuBiZUabgHaa1whWpGlVh8QnP+26FXlWx5exaF5lecDt/5
DmQWjlCSAzx+EnGHsI+Ko5mtkwW2RbO9leKnWCChBo/zOllh5d2JquvAAogWx89k
j4slICoonuz/7BCYJC554TDChJTNsn+Xt7OUTQBV3c/BRCowSZpvxtiB/9/24fOW
Usw2Bhj/MxJ8qkMgjRUi9rvILm6r2mrPGj6pBHNN/7B3lEMZBF8CMRdjNC8G8vEn
Rb0dqQaKNvj79Xv8t7TQyBGjCOxLyXiFunFD/1UunbkDVGIdE0cSJ7HcKHQ+iREg
GXFsKA4+pwLjhpwR8vWBGif0w4jZVQL6P5eyo1kBXCj/W7AK8f/SOuL3XYGBt6aG
cNDe3Fk7DEh7pJOFAgNWx0maKeoQTxDFXUXGZsjRN6Du9IuS3xWRCXNqi2oIovCt
ugxjF1aQdqQB0bhFqfrjk0JTCBKU57GBnwmO22VZ2lgSs4+jDWd7xlPTi0U4qdYA
lqMCesRcqYiGZuCTsQl+td2/ElekczBuPChq1uFxe+uaAjdHhUeMNqS2OFZru1ru
lsRpOQKUasaPVxrQ81lrFqntb6GK5/ahXtY7kbrj4eeFaR1fwsY9B8y4MCEQdTYZ
wtytR28j++IuKUkEzk7HPjfVFuB/yQFVRZGDWOnwFRhH6nnsXmB2WfEU6ILC+B+j
LYYZFqnKGMxDepEf1L8IOJZ9d9D/ZP/tfFzBD8zPqkbmiqyTj9NwuPvZDKhOyLMS
1yY1rzpv+uvj2Loq3EZ6JrFXSi3auN8gkO2DT0W2bGgEEkS+9m4FT/583GR0/av5
f9XkukbShMdOmHzOqYX3iaddDZ+uk8Acj8Kg420/DThktWXzQg3q5J7V7yw+p3VF
23cHYZIgoDir/vTW8hIkRjc0GclKnNCWzurHnjaywn0/QB6WtI55pgd8EdXzabMX
whDVdd0Lzxd7/yGQdTDW8u4dHarD9kar2M5y3qcP3gIZTQLibxWJCiwggNhKV1kk
O5c5xwl39RwfqhtiqCY+6t8DwbFmlfwx3HXKZhmXr62Y+N0m69+6AXKAd9ifDhJH
RGwLIx/tFYajHH2MUcHF5mauf/S5B+FemT5k9SjhehYyuZnjlPeuxoKqihRU4hJ9
HJnGbgLHXnTDYwZkM+UrY017vcSeFeTxYmFZJeR5zs3K65mfkW4m86MNEnKF5nA6
fXDDEzW60r970/Mzt0/7csFgzkvP47s/cF5I/2/ETNQxdlT8n6kbc5KR7jIyCl59
cI4Jw+sPNl8CufcW76GCu9qU1Lt4z1UuFZGOojzFLJpvvSXvGaROgpjAuA9zrDxt
pK3B+UIz3YAxmo/L88q+YHRjVsmvJX5Fv8HWxyhQqcdeaOtzy2/9pYHW9UFseK3Z
1GQy4Aql7Wz013j2o+9KAR2x043uH6d450CDvoWqgL4ITbkeWjLofxdgK290nsOO
wtB3JR/D4FAt3KHBk/dgHslsyCqDszhrAI+coXR89IxuHxetHWtyjZNJaD8xrngS
Q4Js57ABGOc8hZfzzVZVzbS8fzEunou/C76qN82LfsTe4FldHNzGYAwB2EDbhGzQ
CoxKgnFHyhZs4jpMZHdKrEPxSMJ8Y015W5pIsvv90N+34+nJxSt2x2OcVSH4KJ9K
0iFBkZEG15vEusnQ6iiXp16/l29Pl1MdWGB0jMmdKJB6IUjrB+7kXKkfwPvTHkde
YSJlwnt35YxYex08Ify+p380aosDEJvIDKLRwKQ13kmWwk9F0V7tNVfXcOMR4QNE
CsAcTdv6aC8Acruzj/hUZODATnMHPYN6X/UQbDrVspiZOnjzmX8PmDAIZP8LWlbk
a3HSas5NVpu6wSU2yB/zAvMfUyR8iBAT4pCC2i1KzcXYA/JR3xDeYx6SXACzwNWQ
/huTn8MMt2KhrqFyVA/Dr1hk1UIIWpvfvi0ZIO9FrHj+Ax90b0oTq23pgH7Vb0bX
E8s86kltmWQuhp5Dn8AwIxRfvbbtP8H4oTvn6XgyJtnnYNdBMwmo0pARPY70mPvn
X7aHlGdDcGZV9vmAyBdTi/MdQmebCZs+dEVewVk4+eBU8gfgYzeoNrW7Yxuwmpl7
a2R0L76l/fd/XoPZRJ9A/wi8gT8pCFeIUu62YiuIlVMMulnHNB92vifWV2CpGgag
yejkr1uv9hxrf7w2oVwDAd4bmGRAVa++b7tVNoTcexkpO6/8P+lEImmjpKCqivkV
r4TCYtCMjgh5iHF7Pm8CymxCP71hXA1iyJnz76hC3q3iljoh0ofKb7h8VmgfWHg+
Ln9rBH+Mbzi1FQAlS8Dya46+tLm+mdJqrjPrmg50Oq60guUO+yrNVREbD8cYde84
GJK5MN68QemGDyqUyxmcHWriay1d4wxjr51p7fAXbk8ihXJcSL5Ap/iRlOxnR7wX
A4EomgE6PhDhF2VIySIWuVN+2VABOifWH6h/YjnurRSlCSLJWN6xBljPcrzVM7cQ
E6OcNUZ90+DsRxzKiXu31Ys2U2liQNmxK8FvGwTAEkb2GOO1He11fPMK8nBobKvw
Ms9URpeuJd8GUKrNRa2gmPlC0Z2YHF8x8Filam8xciNK/p9ePOtP9AEf95f5fVtk
xErYBlyNicr/glD5Dp/tk3YCgac2OHRqi1zUdXMHE3lxXl2lNE8iMkuVXD6SXF5/
l8fRF8Hwsdw27LxO8p8av9GrrAan9N2UkBmX+SwYz493oMbL+72Q5W/jQkGEVFCw
EM7Yjng+KnMxj5l0WKa1QNByrrBX4On0ejDrSPvHj3EfWZjYQlkN4RBHTL34awlA
t5NqzPCTsc7+l6NcjjSJUCZPE3pxzImAiTnNYY/Zun58OWqaI9lLZe+mobnHGsvf
diU3Y2ZXjRGiYiQwkkM0GycRuUo77RdKvqiKDe52jqj/7pyaQlARh7Oij6CZgZXF
zeTHU8UUqB1cn/3lW80HDll95D1DdHYTmQHiKDcR+l/KJXjTocXsFjFZcSe7o2VA
xPgo0GCFqCfQ2oE2FNleHdSWiDLi5VpR96JsvYL04C/bcrsskUQlBEFnxieipY3A
fTCquCdEH5/qOkhi9oocA3qZyO1JT8sFHjUkJHT9NhY61TB7QN77KmMCHoD1bbdr
ViDaf2TpHLdje21lahIyHMAORGQj4Qt/9XIYJ7/TIC4vDnKhqvq+EzUnp01FxG0a
4dnylsU59G6euLFkI85Zh2agSw8c4JFsM9Ey5dk7ieC03d0EHryLKNN+M5dOa6GT
b0cHkVOqxGI0npp0/3WqmEYeUaQVcjy1uL4n9HpmfOkKsOM3Od107GUmGVfvj/lk
1mW/uIe3WsIcJS7FzBkLZsoXyUXX1iH2ajZreI7374sG2GR9SgwqpiSvPtx6Lal9
RfsXhXsXlbI11j1ARps77ks28nmTSwgYKatRqPuvVCVON9NTY7aJOP9A/RsqW4CB
InGlQCMGND41cHPXB5r3OtrSD++6YrrH8UqLZIhe7TKld+dFHNFBMKfoF0h7ISkF
z4aFqxbKdM8dTcJLmHm7oCOl5tsFPVXPTxiQYmik0ZxB4L5COGASTO7J/3iEphaA
ceH5MDKH8FPeGS3SrcCjRYsQqp+MqyFr8kPhwK5JkKNhwzztdnFa5kCCL///8ivd
D19qcYPrCvL2ZbfJI/H6Q4GrWOsSpFcwXSMZW36yEayp0D1Y3OnodPcVV6oUzByj
goOU7X3Ca207dD1XagyzORzTWq1ItOVtNuII6zxZxtRfIwCM14hcHvaCE6Y+lAth
Q+0XEDb7TH7f8oi1f9pwnUgH05ymf1jHVN22lL6Sr8fYnF2Kvlnts3bExg1au9Pw
oSaZ9D+ztIrZ0hL998R80zx23prJ6yzArAVcBN5chRW0ET6XVjVDskAta5KZSQhU
V8ej1Dib4J+qDJ5tBCYGqrv4pR1slCpJ1nFcyLT9L++Lg07Kor3Ur9BGf/rOU2QP
DlqLQWJQtwaGW6FSk9haZqcSg5U3CCmzT4V7OiGJ6u0OD7y8+aUtkz8tzJt01CZp
baMIoqu8bJrJaEaqmCmdZtO47xzJG+Pyj6zv4TaN0SK2XexnNYmMnibE7a1swHTx
XDLluBlIlG60bOzvG0JM/R+Fh/jtj4uU+dvoCxeMhwGAMcTtfg5XaxEQZhKF21d5
9w/bUALuePgFsT1+4HI2t1IcST+OWZlnEYbbDxQQ502R9K/6yXnylpdaY+03iO6T
OHQLT8P8zKTU9DnvvdNTmjnh/S5z+0iBXdlztQ7n+Fs4KJdOVq/SYXUcxHc0/gwT
BQlAjHrTt/tt7js0VLLkwobZI/eiVDh6qtysV86zFhw+C4+zBl05zaU4hQ4sbCi+
pGXIfQvl8Lm8WWEY9BeJxPEK71SNkmviTa8mnhpElp3rX2JuFlCpLjDRK0yb9CQV
jr0fHE+NOI+HMCCFqG6dMPjQoNd7hYo6AvVqUeZY+24+EYYXfIH2venvgjR4k7U8
C8F5zUEApGh9PynYqLc2xAaaQ1/cQVbN9XWnir+yMZ502AFYS7jEUHmVLg7CJ/rJ
Xe2Yf80jYofhilQ7W9tJ1EIKfg2XDKgFBhi2ZIuPiEF5T5Wg/FMx1+z1GvQrPIxB
CQIFylyKAevaJCdN+lWOiKLNDUq4xqKjZGsxAaY8jP/pR7yHYLLX3PAZ1v0aLnoi
elIhEND0Unsi8BUvPt8ViqFhLnNlIWquhI7QljlCYa/AILdNPbsuohv9aNhO6ie8
ecCfkbSRlJPZS6oYNJ2gR3vk59amMrz7uy8SGGsv+4opK6rU+wARIGR0MqxeB5iB
7ZlXjMeCteD7jbElKxsgkhx6Ipf2jfZRhnOtFSmFWVC2cwfPAYWieVhXcStcg4Gw
dWdKMKqTFNl+nvUnxtUp4pGEIPeavP6LU3g1u813/6r58ZkSrkBu7pY3TZRpWrnE
q9pklvbzjJdSssQ65WJyqZKqDlA1eT+s+45iIYn+Uhpeu31CwZnuAlcVOZBWj0+o
nBVaFpZVPFja/iUy1G0vRo7Qyvfp6Qj2kDelIHMxFkYkRaKKQnnukXX23tZjnzWb
77xjWdQGOvMoegbnlmyiQq7e0WQ3fQkVrpu3nvn49jtt+7YOMDFXJpZWB1aV2PIb
gFS1M1/ufrZt+AqOcyqwGDZyUI3f4++HLq3ZxrfEsbsr+OAFnnerho7qtt7R9gQb
YQtLzh2THk/mjDikiqoK6616uSDJjQw4Q9vnq222+IcK7z6pTtB4HvJVxuJmr/X2
bn2ZTk3TcEa/IbTldZAWiEkOC0I+ii+KNNQGCkyRAPPaVjGjgug4TweM/Zl7q7CO
AxEVTvGh4Oag2X5iEsH/0slEnCdfQjEGD8biVtJOLcOkov6b55H1o2c+c3wSoX1s
07ZzfB7Sb2YBkjjHdmCgtvnpbVNIlOTMAisv1q1sF4MmRSARxWJb5IBXMAwbcAtK
oYiXKFWysyzMxi53lAwTLRC5EbyLFSZ5o5sZxQnygunPcNhzZinjmvwMPnhqMNm2
K/5ngOf+LDcEvwq8Pg2zcuQ5uymxV5iBOQS+aqJGnOdqp2PUWAXUTd1jcAuc98De
G8nuLjU7d65VmEZNWbV7xh02taQEaJCI+nUXEtRzy+C5d/BrcRoXvJcDFzV1sgFy
PVBOowZ7By9EvxP4q0I9uvWtNdWAM7vpXRY8Asv0uJ2pA8HvrPUJXyOSgbDSXCkW
zNypiMWvY45+XL4vmvWnwc6lVytcDUzzcl2OzND7As9bQFKywHLy2WUgAWfL9k+2
MVgKkhyqkIbzCkLII0H4anCO/Baz0XeNXt3POa0IJtbd3E3LPQiz5iW484r5bKrQ
0OODnIWViOy+Tx8fxTh90zucbPxtC5KpnlWQNj5+f/Vnaco6IK/XAreJ0BB49mZf
LOG02aGdGOoKQOAoEb8ChCr4rMpmkouJv8sMnodo3pM3zbquTNcwLTPTpa59Q7s/
kqkyNtnreeOKlAYaPwPUKwL4K2zMdvAj9Ubxbd5Udvr1tCYeguXZfpv7q4o69P8F
qfR49jwncxgdxxg5vJbnT653hTZZeGNXsx3a5Ksj1xclbzfWF1z/cVn74Q6iivSv
JM0JWfptTG4EXERDYeMhrrZwkSggFBK+/r6zQdVh5ThhYUC+JWF5h/zDKHoQBUhR
aDaDIKeftn6QV0kmqk0nF8BMYFkzaOqy/qW/jsHvAJ7BxSASKSfbk43FrWQ9J0N4
UmRVK6eQiQQ05MQI4oo94Ii+3tUccStCDHiqBRDhB5p9Z1wPoV0C39yBK2REqWKE
wGwKztCPLLfoduCYN3wUCwaLb5IU3jMIAZdZ+CFcbcYWX3Ev+EZ1cGiXyJkw7/Ua
vwy+f6qEc4N7U8lo8tLCd51FXX/YmQc4Vp8Jhdg7VbSrVZZZ0J80Vo7NsJQLhDi4
8fkcE5pQt701H8w3/7mX1KEl9laFy5pBYy5rcvUVtqQqQKDw7+/AoP0hHFAJhlxG
EbXpM4lx6wgzMkio8uRSeghNym1n+klsh4+uNb9ihrqYP1Te3DPdHwxtE8yDsIrn
47RJodwNfla9hk712Wqjo6MAjrLq7hep8t8vfO3QKJyScT96gm5XAbu1Bsh9oprC
+PMKFs3Q0HXK2jvOR0lQiuvniFfTwhLeO8e86eC2tvMFWAvIRkmrds+/eIamGrdX
fLqfvsQ4MhCuH3wEF0kxSNlzhU8z/m/i4v0A7eRZSlGnCPna1v8m35iaB4dw8QRo
62aFh37WWUFYOWZCObcyNgAonksi1O2P+jK9Yjk22Qsfbc6N4fJRV1wRsQial/nC
EWAycB40Eokd9FzybmZpyIYLIHwYDBeO92y+fMyzu3X5Z9B8JnD05ow3VDUVtfLF
Z1doDyTMWC0r7TyzLAf5iKEKctuwljA2i9vL3jjn9hUEGeuYoaEdQR0kQ1luLh5z
G2NJEX4Xy5fmfgOXfncMbl+xt4K8bFSVu5P/xsNsz2EhN7GgWeqZlO7cBYZ9ZBZc
t82fdpVtgJiDHQBmX5OTGYw/WNzr10wWsNXgVKWBSTOrP9OC+S/V7fQXiti9uMgi
QDTcwooVUZ/VAxewk67Iw7N5Y8gqVInfcefK0GZKZjIA1Dny0CkhnQRlxu6Qv3Qz
LH7t4yzaZEOGhhjo0ShAi3iMdhdsnqqQMGqchaFJ01HQtaLRk+uRGnLaFjMvJXn+
LF1UMWhUnWa+0KPQ0WtYdbDHStnvVoORGw4fBD5CMUdubeqJHvpbf1n8zDla2snR
DNLG0jXPegyLX3oiVlSfySQTd+/6oXqtn8l8ZnkUQrxVI0rQVBMBBWsCoks81CHw
3pFobBVCNsYBVLX2QDweio3pm0EcK3zQqlJR2Eg21XGi240Y2r8aXHs/8tIA52uq
1HtOCDB0oDo7DRaR1ZNIzVCiRVI4TQMe/rfm3ybxjvBbOBscCleeDqFTex19WKc1
lW07p70Xt/6+KmRKeSR0iWb505d2GlxflJx7FiNA+01S7n9O9PeJVRWsaf44IIl+
KmkyGVdnyJwa/9JTYGpuhcGbGuAPQNJ70adi+PEsJJYDhQS5LvdC5BaUirasaRPS
ASuHMxXxOKhAVcuG/mn3M/T4ECl6elVCIOq6qvvLLMqD/qg8YRIidx8Hf+An7/KG
tLDOgb6+hitb5wd920NcwPfv6+TLhIBL5T07jF+ks7SNutiOPYx5m0a4OKgIynlW
mH1OSdJY8hA423RCg0rC9CjNCOGO+Zw3ECKdZXPSBoGe2e8Qbi1dnzDaQM1GTZMs
i/asQqkz7O7WwaRgYFaPXinrEITen3R7TLUMxB7Q5kALLL3phALikTr+XPKoB6yG
Kw9ELc8KXbUfb8rH1Gof2oHEOxphyQRqyO/mJhJDNFMkF4a5iUL6NcNIqyx1Kn8R
Zc7MtL3EjEpk2IVl2EoXzGqemPHZh/Y8DsOQ9I9lBucGeZEnuz4Uwh4FTMD5jdUl
k8yY4lbSAMk16qFteWmOykgd/hbOamL4cMv4OGx5uiJCJSVzTTq96UaA4s4ctpmH
m/ZsNvGZZdgq+gC5FsGZbC6XTryqCfP6aO93tZHQ4v/glLn3yIid9jly/Yj4GuL+
8xkDweZsIQmEDqfOL98lgDqIgukjsQORL0+3m1Leh+Vba2g4oJTby+VZdc/agKPI
BWRJSqiG+hTFOXr9Llm/7VsuF12TPSpzH1vypzBFiXymssht6RQgzRlweFFjHsma
1mcrBFuNw8EW7IRrcNA5awnPoGUIfa2UB0fbI75Pw7+Gsewjnqc1u772uitar2Mg
JTHefih8nqgkP3EBkn45IR9wYeX9lGasAtShvoP9KrHLkPmwR4/oAacOYT+stTAE
bKqfOBOn/VlH7nimwcpr5if8adB4th7+cplw1zdSOXzzoZMH10nsuo244WZxT7fG
QkQZRwXBgyakP12SEcKw/4UbV/SHJ7h14wKurhWBN2hpMLJ775KVJ5CG9/uBd2D9
UuAWvrFfO6sVRSHIPz9r/DRmsELJm456qsRWqda1UQPMaU/qYkLfeePC+JJcrVl8
5LAEto8pOnc/sBa1HRXsQIoPvG337gb6ijFN+z+krP1+miDPbAA6odx3qKBmkiW/
Mf3oYf60ptYi0vBNvga4eUWDvZcnf68V99o7CdwgypQ92yKnWs3Uy1q1PDwlsJ3k
xFTxGjmS/hz2oyzdlfg2F5kv6H3Gr3P/B2vftYspgf4h8+XILA2Ygkq89roRpQyL
vzNSnaQFsOj3hoRA3jE0JAGDEbTm9u557dA92SgRlikTvq2FQKQHr3x1ArEAGOcl
cpYguc/QY+xmS/0/XS2foyrH+pTtLRW9r4U+penA/a6aqjPRxFwawOUZ1peuBYWY
neHHs+0DGSFKxrmqaYHTPDRMpoPLMkJGV4+M39b9cmVlJ/jZKHAtMqnMfBicnTtO
r8vU4oPeMyEi7lWVRSyT0mc7wdZl8L0cs14W1uwMEsgcsdREB4RBQxqdbyQ2OQ9t
GATSfMjMRLOqc/acPy0zWsUUCfBxHABEzC7WfwVj2CKBm7k354tdzgoynXXdjCxd
3UF0BuJ3uVfkfJtZBTdAp1iS/8RRrVbA9NF4+GNm7dig+4nBQikf2TxHZDQxQvoF
Pdwol97NlIQKa2yZqHfy/ZN4xj+vVEZN30AtCVSCUoU9xwlO/Kdh/N6k8k1aO8j2
UKk2CmMDDIGWOOJ09+a7gAmp2YHnYKfPDVQodhPOgPGWDUQ4WOYq+E1w3UT2bNxB
ztGtzvx9IEmlxMyAFoDEBlAuZ4NWWMsZNmucZouMaFTtL6jNxck14kWJ14khqbpl
IYxnPIZZw7m9GaKVSMiTTQSjNSB+iaWhfiA9FIcdnkBcdYZQyLKuSP6XS9JRShui
L3YkTt7gKz7z7Da5petj5NXEeZVYJH+/gw7NCGIs5ItI8LF0rVHn5YLg45YCn1P1
OoGPuj/qXsb8lLSO3/7vm4iO/41KWfmR5WCZL2firF1jATwaEIVDuAcFAFgSB7Dt
px1W6rfA+agtbAAlGWYUacX/vUkJTTmK9HWxoc/LjFerVPLcvEcmiu99nGSgQnBl
Wr1VyIfIpHc5cNTY4xHZBJ71L/U2VTRN/7MGR9RIjd/LNzii8DCLOgZqrKbidvSP
XAtwpp3vA4rnuMAcmJduy03rcr6Cb5mDvoZZakdA+yMQp9hw2edbxSTwIVSLdG5e
8MVkRoHQnHEsXrxBLXqg5AqKWB78qvaL39An+a0a5JyNkXkLsUGTkKB3UIJIFFLe
2pcOJe/cRo5px3rA+ncJxnFrgNCuJTCyQqgjo0L/RmL9qmSF8UfSACqBP3sYfcEU
KPJvby5FyakD47801+l9ZnOv4DPXqUjN6hv1XAboPoRs2oK2EEMLLlbbBZNF8Y3U
+iR2c3Kvgf2NqEDzhPR9tZuNQievUAlFi3mua57i8kjrCHhaExejRbsBzRLQ7ihJ
s+dqfHnUjI148ISq23IYk9nMESSxLq/YrfhjWfLYsPziJSNH9J4bcv6OEHC1DsK6
GTK7byOG5HCvZZyI7zMjcO+adr6+moFrnm09BF/yZn+55VW9IcIVkA928/RXBwdF
Rco6mAnDg+jYi2aG67rHD8+Hf1e1L3G23NH/GfHmPkil8qRjFWWPcLZl5DsVO5N9
PmTE1qGE4Riv+MFGhOdwAZ8kZXx9wDB2sBcUGBSQ6bUmXO8n4GeovYMCdr0KBKJc
z5kAGC9QzcyA/n/878qOg7klvFoYoDdM4fGjaULGfiogS0XTH8ArgR4RDFMzNilZ
Z4Ea9qwrCJAcZrG1AC52qJqHNAAhaenoTOpBSLhFIpMea+BIsvun4mya8yes42e/
D+8RipX58zFVievY3biZi4lQyZLitkFy0G+ufV4+N3CIV3NI8MN7pewkeNcUQ3L3
1jjdeCIVR+UIkgONfhKj8BvKUtkfBXREkj9Ii8Np5nJ8Llt45vePnd6pzrKP+6KI
fGRBPr3cpMfZs1rTigZT2Ub4oOW/wfouMMQ5zbI5bEOWv75Q4tLWOvf1b4kzXB3C
Cgvciq7FD56dhYD9AFWYqqX9shVYhxtBWRyCWpqx8RcA1Aj5psX3yKS3XfZIWbTT
tFHt/J0lQaJZqjAxPm/cnNYicr5H6isv3hz7ORz4Mc3XLlGHgjcfXlN+ncaZmCAj
jeTQgwQl5zHRE8FIiFFOr7H/BhWv2tcN3EmIOlpHCTi++lL9UVkxWL2KFc7RNRbb
A2tnMQGnrB1cUUNzaUaZtyHD3bHatouDmwbcRLh9hXqYDNS2tTakQHmVYRZ2hiQT
GydRwoYiJElVIm3u05LnzZio5bhqWtrZXN6oQKFViWFqAGB+6WNGey/1Wk6YIUEd
hoKp5wLmBM/FGtiZF+JwHSyB0qZltQgoEvfh7nlB+/iGsvBRxA+DQSnB3wL3l+I4
No7jtyVaSMuF+kuncZAOIdOsm/UfPnG2OJw0IOvNVBkVnoQqTkopNYa8gfgvIHdt
UQvoBLxWrMbfyjhJSmMQZKdX++GtK5Z/bmvuG9BUtOLBYdKwt/9zvGZGR9wvJAdA
bL0dKamYciQb9ObRskI9lRjg0ZjglfYsIVdNgAJYaQb91xbmvFnYa2uxNz0jXFCy
0RPxo27jk+B8OyCcGuoIzanEv8M79hGoxcL4obRZbEIUQFIz5LT0qUebdcaHJLmu
wLMKD8hYptNLRP4m5qJ8+4HXiyJdxmgnLUzXlorQWM+lbQZcAfSmkizvZgTEJEE0
xfVY9iqko73Sb0zgySzyVYlpYd3RltynlyMwciwHoXwTK/sDRFXtntBsyeNBYoPB
YP7H6FoBgoJmzBmkP/jlOcNZ7gGueCgNRP6JMGXaj03d/LFpxl1uLXc+NQfJgz1U
yLFCOl8h4mL7n9HYIcEmYvHo9Q/eeu8/JZ0yKgQ0GwCuZWBhnRR6yuOQ4a6VByHZ
wPxxmfD0l8Vx8uOeYV4/VXeSBUmthhTOQerg8P6sxgIW/Tmc0toHLElm4BetNeai
s3O/Ws5rY7Wsd24cPZA2YrikULzFNAQQuZAzyp2EuP5hf8mFUlWv/AM2FfDzWYHg
j1lY9X4edP4ftkSre4Q+FfdULbgSZOKKeILRjtxcT60Z9JdLlPjFRGvttIQ08Mdn
vydWt7PstZC28Pq1jx6iaG63JsvY1Mc2cCu/GPz/wS6FCxOFIQupKhZV0jIEtOUI
E1g+AZcnxi/v87QtGVdbh21JVzWpri20UfDtTswrRpU38xuGBsJncSS1U6f4J5ll
ld6FKTzcr9ifDm9vMqiPwkbB5K3cZViTdGN6cCvjrPhvrZDHFzSUkdg0ALw3dLLi
nh1whYJqbLD8nIhvF9lvS4U+srtHN+Gf8o3G2RDxJKMPL12Q+GvTXu5bEtpEqY1F
FQZP269QErfOJJkPnUdgdwF1GeCIwFonMq4qcaku3I0YDzkrHu00ffqmj7jbSSIn
TIlJf5KDF8D24bZM+aHig7hn2D02IZPd+hb9sBLArbVB6QFiyPEJVGHd9N9WNLPR
rjVQODDCif4gZTYAq7uRE+kOfd53DscsNEI+vrg82PoN5haUKRR2I/9vQnI6WEgE
ttR6Hwa26KjO+D4mRJ1YbP/BwzY+kg2CGynoujI64E67s6eENoqxXxmOLSwxNHCD
aXHfXv0nDSbAN2nfJjTMRwHCl1A3KHtHrwXs9tLPGyAgQFtg/meENo48gEL5NbjJ
e3Sr+XAyqgcvbcMGZTIWn4OR63hjTHxY4i4dFmKGQc5+lk0DPqwtyBTSul44l2DD
4xOZp96Tgrkf8MeV3VZZ0vwgv4w6CNygZWQPW1Pf45P+uAeIHpbll0CkQSnWHtfL
FpW8zSS6Jgle57pmwc9GcjRUkCQOOcy4ONR5aELhFBhmncSXhs0UMTrtzldhh2GM
Yvd1tcqXrPpGhYN5DXViF6dfeHfFOGS8U4d6t14LmQiJkCkF0Oh8uiKgyOnhsl5a
PWY95wrc2czntRCSdhZ78f7it7sGS43OFFg4HOAt0Ep5/Pszb7uKUef/Qpq2JqO+
59IV+Qjcbj0DzAKeqLmnym6g2IahiEdwWEBDyT+TndSiy2HegxjK+zEqvcY00iam
+RmBzSsyLl8rekNPt7NmAk0tF3A2+Rqq1ROsZdb5cgTVAMgfzFpdPSyGRIVdxQ7i
TMQxN1DLbSWU2Tz0tcydl/1zprsvSm3iQ1f1YWMvVoMuq6/8onKrTaX+9TDdmFSt
SPFs0oTCXnJirRXiHoUSOsBXGGuCBv1/KcpbvqMSxvMavcm9E77zYhxHTC9LlY8H
oFUgachagCLHQU/L8eA/X+H/pwh1QtmNN8+uihY1nvpVQvj0mC0FizdexMjdQBlg
lCDbBTPZvqrpjJIvX/5KnDRMiAZYw9F7GqEDQWwrTIEee4q6ysSDLbvYtV+Wt7we
qyMLUf1ry53m0O5lgVX3OE/4GCK5DquZw0gzd62lhlL0Wlzzp4UKrfx0uelttej2
ZRdD0TKorNgH76CG+Dr+80Qhcm+e/1oGaTWsGsu/wfWFMAzUlGcx67VDEGysPhIr
hPUtX5ad1kWUtvGd8rkUGQ5yJhG4iNNjg5yyTvylWCrH9/1fdBFYlFusnk4ebQv3
Sw1DoLrZeOCXh0dOGnryr0BAeqcrAaHraMP9yZsNyGC6Sn4jTHTbbU478H8MR5RG
exyD00B+jUZKRyqku0ySSww5/JkQiZQLdp9+QybRFIJPU3wJjvQye/KQcjW1B8tT
JPo+Odj1pelJXTCwmnBAzrPtJy/tI/eEMd9syr0ADS2vEcDfErpTsAZiHSE1i8kv
vyDcjLvzGucArAEDk+5HInoVnAagzNlDKF9oUS5gXsocp8+BSfdfzthNWBk8nLX+
q+vzm/TJo/aqxQHfU9sp7vwUy+8i6jduo7yQF96DJOQ+McpOsjQa2mRwZK6iLx03
4aa4GH4pDYBWrOeutZbfvqFhThIaQSiKV9nTrbyLTgyKm+W6mk3ydXL1dZx0Ei2p
b2nHrBg7vm1UtqMWRIFT+dpsfYcFcTTHzma89LjZYxS0vxKiF7YXgv3wyxxtkbYd
z7QJmFwiawl99UM5DJaO0Wx0FuZ5GMB0mkZ6WGURxWDp7c3/B0vhbykqNm+pD9Ww
may7uyJvOj8v/fuFWmmJAP7YgrYZArg16fDYloFqSeLiJUagB03SZKXqeRWfZ7Uy
+gHCTG8AYiE23DUH8WdiM9wKJmh6uPbegU770S4gimLKKLCA9MDcWRzOjrYAF3Vv
UIDzmYegf8W3/cakIIsKshP+togfzH7NDnQKG8grrPubnwFcbEcthcsufDgmRSbK
EcLBRigyfgUVjiZJoF2YQccdCpvrTRANHIv7uTrgVSHrDNtpAR9IyXyHbguXiWgf
VLDEbRRLliZbVFeKr94y/nrlo0rE+HErol4xSqes4zrRoCgCpZL6BGIhmo3VEfSV
sx+I1zblQ2N4+yBxu5NPiOyYFG8UIRWJVEthirF87q80FQ3mW0Jt+IXT+ctsOF4T
wTovc0yTJ/ZSuPtWvHMnoD3Utp0uJZ/+H56Gz6Kgh59mIMs8ixh0SO/g6APEprPm
Gqg9pSNRe/0HJYcnnn2kDJcylJ8oQy+oxv81GGZd2Ca/7nrzTB8p2ikFF80CCOiM
I3coOwtRPW6vlVPTwvxGmROv352ye278xSHsYFaZxxm7s9t0SS/ixrKn3QTZlU1W
Kq+lJgJOZxwj0VL98M1xjI2spfrjTtCToqEV7z6qdq6cilf+3RLOdjZtyQVSy2Zu
yz32W0sNTJwLPpREwpy5pwuTE8yUiN9AcBuoI8tBBZFhxHZ0TwL1Ea/WkphSe2eT
bvQaupFb8HemP2HIVK3cHKCgxrRz0ZSuUUu9BwovdQMFZCaiCY0v0TSsTuHfmr/V
8KvOivBVdztI3U1TdKgO4jTfj1XrgbU20EEe/jtQ7y9LItb6u1VvK+hisn7cS2Rq
JkhyZjqdyAjmQIU2f4LV8XRT6aAS4iMBZqIrttfO3fcvUFqZJyTMXABzVHHb3pZe
wjBkx/fo2/1WE+pQPWK29fBifhatXsLawUUHA5XAmTqJMNNaxA2ghw4YkT1Zh48Q
SN55GFWTd+xFpUe0q9C92/D1sckG24HSQFN+IrvzPSA22ZEUfefqeVqPrU9GY3M+
WJrtHdzbYautsi5VyzmRHKmJho8ya6TO8BS/VnwG0NZp3SaPjS2ol67rNz1fylZK
mvxNe2UoaaDsgMdCycySlQ7YQrE3TIijYb1Zsptk/SBIWwQ503svXgBAB99O05aC
vg/PZ64hkVXwVXcNIQnq+rmSJJge/S2eZyqIxjiKRbcl62B4KmqIQckrWG25Yub0
noOL6VKqIuLUDq9O1kbgqbkfa+KnsWAxTFBco0D8qsD+vrsNCtP6LYliCOKpTSti
Yo7lPdAnkHaDDzNgzy2R6EHE2VeDQfPESsZAjBRwdr9Cia1bVdDLnYqqTAwpss7f
6US9zrw3uLgn2t5QPgH+j/p2Rn+rrheXZOj02pXGKam4ZIdsqLaxyGva8TKrv6ms
xiIm5e0jiZjUHJc34uyEm/WYoiHo0zwVd+XlGeQpD/ou9/tuMU9fzkm9NvE+8U7V
dXPJHOsFAaJAz6A7eSvgZVODh+eCgfy+AYHzgc4QZVRgRZIFjUZwUOpc27Eo4fX3
5Gvn/Xu+fpW0ZhkuwiSji5fUKbVDIkFFmiapPnqCtTaOgbLgfpEnGgfrWXUbPE/A
cKzhWkfXE4udYAUaq/FauyYory84hQmmTByDHGsgZ43IhBcJ9WHoR6fm5WaWoqbI
2wcQfSnB55AO2EMkGguhLJnLny/RbNWMxy30XuntnKbx5saAW0R+SMrqz2yf8jb/
bZuHS6Y9kStXyzN0cUg9Kw2OQsSMKXLYB2fMGTe1BzNV+Z/MlFOxzIA15wfn5n+r
Qy/iGu/pmcC95c4z3CUIxhw0PIq8N5rrkjuFrIoy2C9BMhWSZ36kTXrgeaU+j08K
u/6GP7JcRk73tT+ml1ucyjGgsx9aiy/xRk9KKzev57dYMaeIzR66pfEvy4E7zkj0
yjqPDuZ85WC8iziukxrHq+pbslEVJwHYOADTs2tPHNOoM6JsLV4tJC60DZE288fV
AdR2zhoDochnTEqhHRnTeyoA7K+HhnZzTXLORke9gTxwaB3aKFQZ3ZmZIm5Y28Sr
fGjtMD3kY1lchNnau9kHi/3S8PxKG4FO+/V7B5L4yPvvwiWKckutIauNO5Jdv/A4
yI79PNsprXNdV7a/Ta/fHCzUs894l4jOXaLtTuw8rS/ItrVBco44wO1+J+95zj1t
RTEPRXKAufVTSOdk3FyVURQf0h+zS2Bk7hz5JzYenCqrh88ECnF86KG4bZCX4S6d
O2VYnxExAk1zjSdJal3lEoJQBd6szvLZ+8dkMbJCExlbPbqTzGgDm8EwWuNxYYfZ
n6E3WUh3MP/LiLuFQ3s6i09W8/czaDK8SxCEqhz0RihUV4kZ6bK2bPiUQVhcfjdi
NYB3UZ+Sy4ym3UG2w9nrNCFtGLYPIHtSGNXI3LL3GmNwGCNojUApRPDacddcMEaR
y75MCf+HSk3f/e4x5Rnp/y7216DLGG3fRVn9ghGp/6+aSJK7Wsl2NWXEp4w+TMO+
dVjkZf4B7UOxFqNhtqqR8nLQet5azhWlxXa+k/yInT92iPitD/H6mgAw3FZw29+C
oczEX+xzXWktI+dOobcdV2PMhnNkIVOvpZEmiqSt+vF9nzQocy8qG0l3tKIWx40f
cx3jBhW1B3hp4yb5xpxZEw+NFTIgZuyLZDnymSCt7h4jYk4+neOaHKj1Asc8RLIp
sUDkUJlCz5hFfo7tecnVwHMR6plz5HJ23uE9k2WeC2o/AvPiUzPToC9Xgrw/4Imn
bAqV/GEmWfO8aW/UAhuJYqRcTBxRlS0pL/rzAAk27ok+h/C1TiwOxMFKB1QtZhU4
9UONMoYR55MaeAOMSRz5fBf5lguHRu76qZIGvl778F+f8vX3SUdMsoA3qsL2+dk9
1+Mq8x/ssuhPNa+1qX8tqT8oyCrBSkQMcwGc4asaemVw64kOBkRzFw6ap/FevFFx
/I7rd8jmoIJOBPG6AS1+0W1PQm5ag2RB8ikrwO52B5x6gWqSR/Onv5Y5JaB7og6f
H0W8WHmapin5vmox7CFxQhb6HZvt9vKjKJDzSik3bdY5oxBR1T98JRpJ7p0E6/EE
73lhUoFDwxnIgWR+uYu/iwulCDyIh5pABHWqbUsQTWLt7KbRYR0OXkM2+uHj97PA
+SPPkISb3ySio8TNn5vUC4aGJgWbXgCkYju1pgDMm1ANj+L4IM1ihsOettEblEJZ
q61WNtPfArXO4PSGt7Uxtnw8SAyrdzJWwQpzWvo5NX01FG1tF+aEXaos8uNVX6ng
kTeho6QTb8S7G3h4SfOd/f8rDp18+XbdyM7/WuXD7gRiW9yRdbk3EqcqrYuZKieW
UAtXnGi9KmSF6nOh7J26sy4JYuKWVec1mNye+MhtcKKW80outkH2M7rV8Lak0IIo
tK3xKACgV77zME5io1VtdldohT98/D1g0O+c9WKngFCrKripHhgINZqVMJDgPGGU
GxaKsFFIp7EwixDMraP2hZ1TyaNBxDNB7jZ9QBoM8DWg9UtemcQqLLqfegB/FE0u
7ydlQKIWt7PugnXdAZCT57f93toGk7LMCFu8pm6OBEh2HrfIhmcbCGti7IJtUq84
y/lTxrcJcZfkPeNcPnbp5AITpnQLWHWcA0gWjVE3IoqwhxcvBEsDLKmQxOxdOaAQ
FWQsR10OoOssdGdco1Mi4jW+fPG06B38Jsksv+fEAFSFVtFWtT7jFDH+eZ534Iq6
1SFh/yO7nDfZoooxWkwuts2uG784E37yeukO3ACx+YGrzSvRJshd8KCnTlEuf03g
qggl6aVvIH5H/7oy3ZpYq4xc1E3JYJIisS6w6wTk0b8wAURuZZd20l6UvZFpaopP
fcdz9ypMEz0Jgvk6n2bud6jIlZUut5Bz7DqhI9i21AMLQC9e1m0Jm07fnOvcO30/
H5Gko4NXVjjRj7XTLKERrl08ItqLelgAORvWjCWsBpFHd8cIWX874qVsiFMwZgTB
BTTRBrK9W4KCc2zefTnh3uDVwD+5Ak6lsfitxAyGZGNpwhuvtznU+XB/xGlCbPX9
gRQIIdbXs0mYM1bgulLNzYB0FwoyKllLaCj7O96a8PEYxQDW1XJOmBnfjjIMCWC2
ue2TUNifzXbZKex251pHB4CHluBumA8/M3ZREjYwd5d7JxHv8eR/oMNDWHu5JX4v
MgGX4OTXgbKaauCGXcJFGFdpUpNDluUPR/2iEXbGTfFOfGNduAqaNg8nHBogSdb2
pNh5NMH4bkevTd5+zwBHBvE9bK9H90TkHphDJrD+LofV4WKgmSYGC0OA3E9sK8du
Bpb8vaEPsuyrHZGlxG+1GoKHXNqKa52G8aS5KPPbEYvURVPMJxC0T8i4r8uh0Ywf
dpIHdCd9PKERVuUvENZ94motqdKa5Ta+2fPo8TnpLGfk0Mse9EXD5mZP6tE5UlY/
pClA2AUHJTiOooJQkMKPGBEqzBa9RKn7UBdn0mXxN9EJ7SDx9of0Fk2gZbKvsgPj
XhTMWZ/inIGSCRkgWEDXa52EoUcw7PnrMtspxeu3ueHB9/MybY4EM8ZaIkYA5iM1
SwkRC9MYxx8aBKaRFmyHJLmnn0KI8BHF1nDWG1VOEQC8SM4jmT8+n31KJXo/izBS
F89nZsx4zVFbSwQZcwDdVJvSLGW9fJRdkIJvQmgCbfikvqA5ibpKHvgLGZ+jsHnM
GSnoGEaK0F7lM2+1Q6o0LNOCPdl0Vzty0mcBXA5Ound/40rfoMuvymCi1NbXFA+S
pm6bGaH8gnm8BhOilkxSrIXtLhMQR6/nKvS19HgpqsXKYRaRVAgBaq0E0IhAic7A
u4VqVM0zCsz8AuPkqcu2aUD5mnfcnLDKhY3H+ZEw9xiAeMqt15xtZBW6VJoshRoN
3RSWtychLq0tSyTF5N2PH+zn8Zpei/r3fXATIdEpdbnv6FBTVnlg71ASFgFUSXIF
V79lUHFjJxLmwTlmXn9DYa3z9iDuIqlnAf43Wqd2XdAGUrwfEEJx+oFU4F/pjIzO
iQOiwU7grEzNKqDqqeDC44rpvlepqAqquPCpIPsVX1NxQ3aoeC806imyRmem7C3Y
BnEgeNIjEk3KZJjHtDpzl7EdfugULIB/3yLV622RUZ3sPzBSsej/FQ1BEOc2USzW
UDLFfYUeAwNY6dFu2FjnUC7iZleYFqXAPz0dpij8RzTSQzmQXwum1GLfItwEAVB+
9/T8lg/jm+9kJJfarNhmO8fZwrfVWs7XkoZiw1caVwhJwlL3m7G1VaQ+1exdFsfq
rmabU4tzjVYljN8MuJIJPwF8xurT+GVtE5/aBxBRs76GZAyXatgIX2Dew+Efw14O
kDoAUXdT5y8rF6DpV77Imj/3qHVhVhe+LVbWhejlsYFhh6lMjBT2kwjUOL6A+jmm
V5D1++GzrwfxeMsODaCeubhS76FExa3gg3YCSIxYosjAfCuBKlB8yV1JZwMSGWnD
DBlcP802P551tiISqX9WUdSzZdotTEbwf1rR6maShJs/XgbbKdeV2oIHhccs6oQB
z+t/0ltch6Ks4O+3ZVd2iWUilA8CPVJglSE/eOLGuu+TOc2PRE13PVhCrxkoFxqq
fnM23R6dijuTLMTNX1EdijGI6nDRuvRMk04D/cTdsMGWGc3pGL+IAQATh4qQTE2W
9J4nH/bYqVofJa7X1jTFcLF3G/J3vH6xuGN7El1UQtYga4E03yzvvtcj3k681EgD
YfxaUDbjVS8FEQ6pg97W1Z3O+HgLtsctev9HvAH9eAdwYqE//7fL7/A0DfdHF0TR
dq+5LEzcyf/mz2E5hRgIXgPUSWO1FRPIJbppIFYrBWZRFT7K5lWgaer3n2lVLpcs
jf0/xrxGDdA+N00i73Z1cSlKwmw1tgg/Y/eHGmq6AVeRLpd28MBJOJDYU6z/FdEC
L2VgsB51axQAcWozTJ1IBQBchILaY1p1w8oxMVIN57yc1KTYoKFh218r4UAvFfhf
yyyzwf8L0hCkL43Rdwhi1nm5Y3tgvENv7SLRqSLNu/w29boxqthen7j2Rt468cov
IlTalK/wdgGxB/f4UzBLPX4/gse/Cz7C5A44wtPdkuoUydIp1yoQmy2MvPAakgQg
SSeA+K8XVOZGNeFcaoSIQ7N3FYV+IruqRSinCPnKkuWM+FEHgV+YC3kI1SvvhTks
3PguXjfgzWNLFtK1kbB/zKMCpdU11n3at/amHbrC53oWmVccBYgHGvN5gc8sFUc1
TIq7y710a47vrQ6SF5taHMCLzwCLLxWC+J0lRi7G9jbeYM3pGI5MR1DMmkxA5M7Q
t2awulAIiSk8OCP9fq4O+hj60TeocEvKH+gpf+RqiS4cKXOn5IORsdwPIJLNrx3M
yPSBKRFpHkjybXaBqw4LzhOcN+ZVAZTFBRMCuaiCkkubGpcrDx1lHXzbSbqEkk+3
PmNObgWv9/3v8o0oxRXOAJ1fQs9P+U2VkYtwQqag24obavX/14awvIyqzDxX3gAN
KXs1do7abwqeRePmWllll/Umo/rSUOahSC/KLVVfnuIYxaUS0mH0d8gARea1kEMn
apTUp9tco51kokaK0JLUVtvr9JVJj9m3odNKiqDHjPeo5UBn66tXwFSo9yDm3Wmx
avjYp6N8Wg7hZ812ec3xSvQiEMHwdJfXs8HuTgKe9XlGWh0FMRnkKj9fYpx1x2w8
CA+57bzUGXqXn+6q+mIMtDYhOB5EdoS/8TzsXKhcy+YcvggD8rPHifK0EyWDt7Rg
lyQpa9wNUSDQ2zAV+S/rdXulu1tUAuu+WvjSqAnzdXp0fom7D+4rk6m/0Jv2VwXA
22mszy1m99N0Z85m9s2x33SjJrxNf+XGqFl7Xq+RXdFtfgJ/w6T8vpI0aRPg2JZa
XckaYML+D5XEq39hDNCYTujUrpkbZ373BUrGq4F3PBMMDlkWfugnFYzJWeo+cP3s
AM07yiFW7BBHwWCbPtd1SLXxfIXZ7XTWO+hBaYg0QTcE6dF646VLxJkmCVSyhvGC
26CkkaG691jCt6OKdYJOQM5rs0cU7SuQnBMya8wFnrY8vt0wxvn/gWlN75D+91Da
nTCaOvxTnEr3rawQ+rwFP81afmohz7pDa5WzZaotK5VNsTo0mXEVUb60DNUGkg2Y
pFgqkOtbZH84dDv0KCgy3/rkED4m4DWjs0VlrqKk0oEURYN9If2nz4pHGmuHdox6
lebGH22eP42c6t90TipI3dtSS6uP2uCVKJDUSqZRYdz9GHKDq0io989tfDZ3zuwz
QP7m+LuT85xeIeZwdM7yEOHg+pPTFyq0gSXVitiHKCOh1s9tQw/BrgU0nbOWiXD9
SXHvsdhu5ba3YztYyv28VjrCfAuWtVlvo7xIbgL5R/yLXuMW0caA4LgtVQ3680Tr
IlN9kxjm4ZrODqLenM+dXFDNQgPMPHI2MRE+yi5qDKEiKtalcHmAuv0h8MTm7N2D
6oAP9LBNAuFABxGDMobRqBFCYwdwEcym7wScE+k4diPepr+vbJtASdjJs8qsG3uK
Q/jp0e8bOH8W2C5hLpKV/1Ljed0en1IKMvTTf45oZfIBoQK3XPLeKHLKn6LQNdap
WEe8qpda1AH3C/CfPHBMCxI1sHNts93IuJNy+6iEfnlcgDNZ32mpesKcXKya/yFA
tu0Ov2rxuvq1vEbrBY7WaBXIA/McZlud4jEOR/hdjWVljzzymMn4n/uTcLT31MYL
V3s3XBBhFD8FnoJ0OrdUaEGQFBpvVfz+6DcHW2bUzFNPq66e31QGI8CMFlhJvijO
BjPlVVqpt6adFjR+tG4daiBE9zExnSjLPfgz+K5aauMctRcUlJ3CH50asBhxp6OZ
5FfXvtj/u37U74vox2JYuLPt85vfuu2XBH3Oc9yQ5WTqxk3SqNwEiWRfsDzOgZ5v
JBiC0yUYZlenF4qWi4v9w8bpgOqzp3XWhZKXmdQvEv76+4dZqFMdFjtTJxqcVAfz
4hVZOWpdUIithJlxvAiH4TLJY3dxifQ1y5//CuMM7Y5Vvkvs6fl3atInR6S2AB8h
B0fScE3yDkoOvJ4QJ9+ZAwHiWcKUICrFjUJ8xv+z3f9zX3HngludPA1VvB5jrq0q
hI6bbi774EN/3Znxq5m7nrdLONveiUw6y33CpJ6CCfzSHW08hD1HKCCSNG4buPSa
kPe1S2ZKYcUEWywEzVgh7DDcNGJesdLLQtUv6IocbmeJWUMHqIgTFGA2cmqcEKTN
LKCtzdjQAPpA6sOjuFt/ktrcd+bCegOL/VLcJXQk8W5kXLCZ2/eW2qqZC2m27Iw+
JTDshNu+mzDnDB3Pg00uKkibjVddZPf6aeDRF4Rqk8hKdUyW1T+eeeIiisaamyIo
OgN+VPZHFw3GETAVK+nzYLuqKuCRS/jNylKHSOcrS17BLI1EAY2NG6CMSszE3Mz6
6txsYnevrvft4U+jLw5pwnZXC3X85kUH3QrTy7bJdvwR7ygkWpjCQP/tAJDZvOLe
Pqsg3T1L14qLm6QLxni21tCqWdIfqXFBYihDhdOThf0XlRLGlTJxlxYOOk93qHvV
G79rb2+j0wS8A8CAZygNIJxUxL5PiaQtCXTVWOGEJWkXOWtrUSzyQj5kza6MXfjG
M3Ws+PnKpw8G0amFDzc3yftWeIq7TfKyiAsImBJg5+iU7ECyUrKjaJ2Zb3gXrqEm
fF0igsjeJhezEU6NShA10WZ/CojQDCZol6lvHJlXqnYH5PYW678Y15x+EPjco5wz
P3BF4FRAEuW9jjFo0PwzifFfsuQ0QOo85UIMlDnajP3LM0EjCImYqqrmRkp1ywU9
vo3dIplpvUZElQVWVa6/kldodX1kx185UTGjN3JIO9DydN2A3GzxgVCv6QokZiQ9
b5c+SJiIQodM7uFaylm0aWtTlwA4X4DH49P+yR7f/5CMqqiwk6uucU+pnXowU4Fq
AowgSrXYi3rIFSqZHtqRJaJ29CBGwO0mtcoV8xYfKlBTvizQ2RnlISlZjmu8qCvd
d8SZAhT4mJJSksju/uFcWKzP1JgPVkIjz5q1kRPwfEYgXxCqyyQCMzor6ovD5hFP
BlJM/G0wJK3smdawq/lrljTJqWgW+v/jZqnkOYrVjc10va4iXRZg1G+TMcvCnacA
YzOz3Alf3AOLJ/HHTJiJNd3Zg6yzHqKRUIpfArPHaw1jtzw+21oVwugL0ZwZXuQ2
7hi7NKNGME6vOcBEg+OlcDK4AGk39U0jjYRkvpgCv8rBfwnnlPYbL4pTrLHl7AZD
xiPeyQMSLB1nRA/wJk+caGTvEVsbsC9CpVrTnioUWS5qbInFgdCPGQe8UIJKrYpu
Hu/85wGlVkjOHTGAYg8S+/jhib4hyY/Ia+PXcYEz3IcwY2k3LP7t/Kb0FUyI12sk
OzaRE4SpnbibQ4rp/FbKVhiWFwyw8vCRezAAEUa9S34La48GOFNdKBIg6s8QBzTZ
JVhQL1XNHWdUQCeOLSKn4+g5MOM1to0nPm4j3+T3pkQ6G8yNXNYBrnvmBy8Gebp8
iri0dDD4s79aqPPH30peTGIYsXGUbM0sbo8wJ5Dwiebhk4jKwuH76HZdhfm0PwVL
wWiYJu5QPJeDmblFdmUvOw43VmV4jxDhDn5jiY9t4+jLI5kRaC45EZt1g8ZtszeT
BiqVniG0/QRnvJeof2uQT8hk/wvBoyOmO9vnJZln09mQE9TRaJjauo7jKnQmHug5
UE3td5kDDj/CdStb9kmmMIzfddLcdPj3eY53KUogTRGWMme3Nwj/md7r5C65VPEK
Ny6mmsMewG+Mpy8bx/3pPjU1IjUjvbmjnCqp2kEIVByRudE7WDGTxrs+388C9LUd
JhFfjnSMHGQlE019AQ1pZ4FyIduHXs+0Wsbuy1E+Z2CE69MGWB2ceLzJcGvLZlXx
MWOae57hvAl1X1fxhggY1QGK8CQofI/1gxp95QO46sL+BbXSNYZuICyF0NMnhlAe
eXhVQseAr+vVGqcTgR9WlysElWZKjFOhRcJj/kgC0ocBleOpEjx9RnUWHD/dDbqB
mu8ksVjXx8LRSMuOxzQAWVnfOYJJnv/FSr2/Ccpi8Oh2q40fqY7w3bTfs8FNhufD
fuL/0drUfkMwhvDjrDY+HJc1VtJ8hmt6e2Rf8D2b5agfHCC35FGRDBGdxawY772S
gLx6MQHaZi34erk86Rgv4WPel1+zROM4yH5zdh5YMpjEA5djC5EJytzYn3v9Z+O7
oeVGb1pHWUcQysS5xeE2mJe10eCTKQsJSBUtnc7BNqiXCVQDLuC5Fa5JX6LvfFdy
OQejhwldtjZSfB/3yH45PdBbyLRk2vfCv3RzjYtuzlTnVCpfZIKf5XE/2UvgJXtd
w3hQEnjRUSZB4AzzaXRY+zHVOcdWIWwzoqgItmsOWrq9ePrZF9xSwjz2bnw4lNjg
2HLpN+zHr265JH1ZDAddqKEqJUrXZV6javpxpwd3bchP2rTyTdkPUDW5jdPOXc9P
KywHq4TaitIhy9MxP2kkPqvTZlaD3UM77Q1mef/tljS7tFmYKpuT2vdt8HIF4qJi
ZbJlDxn5YG5nIc5vQ77Uof9RnytTQ4QRH8IC6A6vDRkqBguQrC8qq0o8BLcDeq8f
vjIfORbMBa/pgVetV699Y4JinrNoch58L2hoRZIs6980Z3s7P4j+WV8h1orFbgEV
+e+eFCeEAxDlv9xd6r+5+ZNT2XFmf1u4fd20M/PkWtgUDEUz8LznZgQpm754g37v
4io4w+BdiayGIatNm5XT7rJK2CLa4NLqnnz7+ywl+HRh1IFhjeOG3RpjWC/d59MV
1OHXEG8AyfWvwU5tNmpBW5XAUoKOu29N4YwyDeNmm5GgvNwenZelRIIyCG5pIqKa
oWxGB7vdL1mJKOFSdgf5RXTyuU7vB85CcwwGPjmTJpLOsnBl8yjPZOz91y54Qad8
yKQCXY/zIYn47tBZ0GlYZw2UHmaejBPv7udvpGcVRrZSGaFoUkibileBjM3cbQqp
LmxHx6jMRIMhYq9UKyAPK6HMtpdL3REp56f8p22uG5rzY6YAEUDnnVx/zBixWm0f
j/HbJz9vuKmfZ5EFeCrf5g9Bo9wNysgG0zK5knYRerthFz6hqVPd/MLrKaJobcmy
QKpgE0ET8P2pnyBBkaTZ5Yvzxz2ZssAVj5SGJ+/0t2ZhDOvk0EHZPVX8MaBJlb7R
HyQfalSeH57U6Z5Gv/ALKXJDAgDA6LbgJLdeakv6uFmmFPSWOtPp/mFx/G9WkZLf
nx3pv56ID5KudS+kRho/qqIO2jZr9vYt/4rH+dHRiBKvuY0Yba8Z9HlAvg9GsTCB
2jke77WgXCGmqwvXsZN7wlr9R0N22Lvz1aRWcRM+bfr0ITZF+FT02MXjI7SHr7Jb
SszqqQpnB0WUfq7qWlz+t6XM/ysj4BxocK2gzyvGTv4jf+qvyWntacUXo60XZtkp
LycfR+ZbhMbLg4d3nkA1ZwngUqtbQoM7sZaUTGejMKLV/Vtn9PjzpOI8T9B+kXSJ
nMzHqVWJdc6JmyoU3uKy1URmfikcLGru9KKNXFJfOt72VV9tsB/iq7sK/4TqB9JA
Cij1Or/kO9VvxSR64p9TfzmQwQ2EaGSxQixrromEDhsCcdMfwjDSnadX1EnqDb2S
+XXSv7m4WGTUA8fLikDvwqUUuBgWh8WMheOOBVIlVtSB4tENRE0xzumtSqYo5rPr
x+zNWabJHbSO0gmiN/3xRdOZCaTHUUw62mjMsUVKAhowI/72qYIbx2Tl0Dv6GNk4
31HmwDHa1VLK5BJMepYmrB3Xjyn0QMM/2Vlq2OjIcCkdfnW7jXF7L8krN32NN4uH
jtakA/sdqKTigd1axpKSdmUWoAzjldn+ARUmQEtcul334VKuJuZG/+M9nF5TtU7Z
NLgKwC3w8NZj4pkEcZsf+2PWOMOXKmv0/rHusY2if9N3idM2t4llfbGvY8n03xwu
m8kKAyIxksXOlhziGLvFO2aLzCJ30+Fx8Xhjjb8UqTnEEXOimB8SOZbaRfw2b4hR
NEzrfS1Qx9AKDvWPHHar09q5LtlJuKgIhqqOv06Mjnofy/gjxHMuGskoBoxpvn0Y
g5AHo/+KHV8QTxKjjhe7NLuBppSA6EpxYpTIHvx4+Q+k/e3pl2dDac4gIJ/MITbI
Mb2fZI71y/kC9OiMYQhlsCuuSkltLBeVHpJBvGVsOn9TItHwf2nSsldtjI5wzgbY
rpdyw5FWSO0AFp4tV4yEPpIgXIVQWkcbie3fuzDW46ysxQLRa9sY94VtB+0YMKKG
HVBG/u4KKiYVuezYoPxttO64bp4oaz2zfXQ0yvpcjdFpdge7SGRbubKzfvcXkulW
v0a+590RHr8XPJzELC+6BwW6yXPKGwF31GPpapp1zLnxH2DHIwHgY6aF6AMDFOrO
Or69YS2x3teanU/XbbC1+PIvnlhAFZpd9n6lNHWID5tyP000SFIDe921PG7CupdX
cqIRvpvneHyBKZM9fOOu9p+9TudblkVgpW+zqtl80moHlXQSawt1Cj1n9xnjcJNp
olUT1EulLd7nvtgfXSMx8djw5hXxxl3LgZICeE3SsqugribsIKv0Balpmw+zXkr7
3gjKed2xf5htCgPamKUm5Y0Eec/V/OdD2mog0xNfretDmdCcQ8mnJD9lNcnlhMJt
TamGUSMH+gn5LMdu1YvvMzQlQ6H+W3GsP+HZz4rJJehCnJ/s3gZGCjZfXYbN7l9B
9cPutvnhaYlf+7GJMa4I+cuU3OR0jqWr2lKsWU1XVBC7msiqEsFgoKlOUy9pqQ5O
a7pmM8nbC96DiaKbCcGCs7PWlbE+z7ClUszc1/5sOG1B0LdwZmcJqPgpTV9EEfFO
KAPPJzL3OqgWreVstrRAfU6PvOb1Z3OQ+P8sCQV4h476HLCCmTKOja7Vy9gXNYlp
2dHZUljjm0tR8BrbiGxJFpKuuYLV8lC+jF92Hx46ZpJyb5ZmSy3206AGXQym1TsJ
A9j/uoUzVC9Cl6GeJvyGtlMX6aARGcZ9BvOBYlC1PD7kjbZl9HPaJgyZxqoMNiba
ea/uRlrPAsgvLRv11ewL6XgYrwRlcmqOEAR0I7e5BCIuGLpJ7WuFX7K13YSQh7CF
bNpnY45/ZrZh+W+KEybni+jIqDz+oL3ohdQ5yAn04YQ7sZvOPWTq6Zpw6eXstzMs
tmQUt0R1Cqc3dKM0e6HyPBjK8DILxOIE8gAvP4pyjPIsulYjY6mKyOn2IQiSSkDq
HIXXVEjlrwbp/DETpiFjfFqiAYaJlQdQulYYd7olV2Xn3dUzJG83SgrUIkgyGkx7
98HnyylBB6XglpkeaiJsFkMfQo75t0LuS5GDwKwlUU5rL3Jpxu0YwaoUi75nCagY
sYQPcLJRmnujckstSadcCrOr1Q8ail+UYRhF4/W8SGH1+NyMQH4Kc8YAn1D7k2mx
0+A5nUOgpOzzZ7P1ow6C81DnzH1/9CENPj88p89SHNB5X6zQzZzcCEQowYeLQ+iv
4Q48UTnbwKFzcz+GyhlxelHB2KIxuiISFzqD1//ictn6zl7n5E3zyEhh0y03zPQL
4jgWGQioyHwHx5uvjJePzAMSueCbYGnwgTsIaYHh1zX6p6MCD3EC7pnuYsPnoVf4
HEEpfR4TB1i0hcqtUVxUiI4Aucb8QpYO7vhWawmaDcxf5Pu5iQhcuiA/L8YCQNmu
gUv46vLEZpriWZS5SN+B8icFSEe/GfE0DGkhLnZdRjAgDoPoCgEAxRqcHk3VkkVG
ZrNTkQ8QIKmS5THmKR6O0SIwZLowRTVW270t4w9gPG+UepCqecaR/O/lt5R75mTy
qExznvoJvSbFU8Rx9R5ZTOZ3KoHfWf7XRCV5HmwPfTUFVjZX3OzmtaainGYmppmP
eS/zzVpiA2cPDk5E6UYQkXZOh3IbKrEPCZD1qhJ28Q4oyB5TSrfYhECJ7BxnoYBq
wF9D6rflTuLMSdOK/16QTW2bTgRr4zo8aAkLGrqbXc6FnWKZrKv0q1pN9wWJhKD7
UOoymLHOtuGR183DxKHJ07i5ZiuQhdIPFr9YAHrXdS9xSbIbATJizh6mZMRSncCO
z1HWSg7GEL59/q6JWD9JGrav62GJRoZArTgp++fCG0AxDpJfC5Z7wIcxb9iCBKKc
oN1YrvJJKWTnWsksZ7lB3l5EkFtLuX4jXiUYWUcxt18q5TvDVC6etyjzMfiVqbr2
w37AOUrKehFQLRGCWJWBZe4wP45vdD8Vbg/TJUUOJs9DJdmg59xkVCSoRrxQx3AD
K2dZN585BJ4YIso293i5f1SKgJyLWTy+fJ7G3MGEQxafPgRuQZL6FogJyV8IBmcJ
KKKcRL7dDihx/sSVVmjSyLlyEQXfv4g48URWA11QdcODjUsWJQXDRx50tyn3joET
20sFP5R2wNZuprJ1KhK1+phNmdbA+TmDWgtCUfpmRLAymzW30qkFCVMB2P1+fSkP
ZfyukqOF8djnksHp3aHrUhLHidHDkxGShgJEsA41gu7NPaU5KLdW7SAhcrx2FCZV
KxQQ1gM/6tgXjran+bbQmHaTXFvIXjECDHmp5L1UWc2l93BZBh4Dg9yr7bTiGy98
NeqZXVu3pOVX2PTj02JqwVaA+ZH/SS8DkiYu6djWlIVASG2n47zNaUuz4AmkDz0j
SobdRRCbWDIY0+nU24Wyetr97UTPj4maeBdwLfgpMnSlRNYaf1+ov5xfOYSYJHio
033bpPU3Z5dzJjMYYrcBcFI2TpGIAo5GeHmxM+tlZtXwCmgRNywDusGpYgny4NPa
GtjTNZtPtXZ8cQofLzKIIsLn3GiBlui5mCPNaCr2iFGcQ/VDf9bD5xupeLETabTu
O2RWng4bznSbXH9fqrnrq0sodfxeTyi6xrwA2KYOODu5Q/Uo20wI+ARiFrGjigZG
VtJArw7EflpPmbu7U7ym6Pa83I0/mh4J9oJUTGEPpY1wcBz+zcgkgu59iQv8WYuD
rqGcRo73AL1WRiQe0fmZY2lnAsCNYEoj6RHlk4NTLf7+FHxblszkDkvAjXKLn8kc
pVh1cyJCcB9KxFFy7n/EHrcQ7k0k5J/3Xbz2CjpkfW4lEbrqOgP17/5bHFPylyBe
XSuReEZFjBm1hmfD8d78apa4IHOaCw54SDroviZMaCdDyFMb7aRY5YKWReTZnj4m
jlMHENTo0xZ/P+jpSQiNreHObnlTQ9KjC5HjpZvtOdU2hd6fre7OqTCXM7HBBSbp
aG4alNVQ4FCITj1p5rYPol0fHe08qX+z0PQYDGwst9tLinckoAzQ2Ifm4bzYM+nq
WS1gYF16NTuksUAWoR8xsEo3z3146Z2PX2cRGtg3WX/89CN0UV5V+qTiI9+6PkFZ
4tgrACFmNNchhC+StNFMNmJeL5nQPzOw7UVJlFEt4IdsdQNoVai3QunWcZN4jMYa
2qLBPIaf2VdQeCE5nV1RvPEUE7tnrOTxG+KNZdMyStzmCXjG/HR9uW7+g3VCEVVR
wA7MtRpmB+K2BXDKNcF5tqcTAO1hBmfHqYSq3saWAX1LGccUTQi+pIqZzd1WEGxq
IYYO+pp2579FzjoEEgGpFF8o9yWF0SZjvaoWMLqptp2Sg4b5Gb36CLBsPOxJm3I2
a7LZLUh49fB4F5coCvgvS1/pQsdUCSf7d0587qVv0o3jD6pIiwitg74qEQdYE75H
4XCmkOGa/+AlNMHEfE7fRs/4l3rQZMUTu1C3+g/YigRV+FphQLiTz1kItpTDbVe5
LAcCgs7paDV8CAWc5dibVVs2ykzoBhCf1sd2z9/b9aRYm7451+vO80Jh98Caucyh
I+4tUqRyaRj3f6th+VfEji4ybU7CfXVfjlgV51frdDI94DDcQYuZ+UT3fr2cQDIN
3b3rSR4IzECaySPv6N4CdmlmY0qlfziLK5kfUXRMoG/ZnK23gV30KeBWgyxVoASJ
pNYE2tmhOXFHohBRmMMx+A0SqCmkxL4H0pnsaOHHyze1UkspY8/ScC30e6oeG9BH
ZBnNvWoSJ6FSw4ufP8D0aWxB8D07A8DNmCdt6dfysbOQgHM6qXqLscjcea5zJciU
ktuX1u5A4wIHD5W6KI+ORkXgSz+XsHmOomHmRlZu6e+5Z9OzBoo/Tppk/eePPgPA
NJP3MseD/wr7r5mlHauXpCk497BIqPSpX5GqeqdspKQhli2VvoT3Qnyd53TxhwWn
CydbQ4T/DekU1lsT1n2Ul9x5v5PYfOp3+/ZQjuE9smhbuU7i6oqaKE35ZOJqGTcn
oYRwoghdn/uHimUw95jxJPxnLEEoSHmtBIbuhuJGO9HnYgM5nEBuTnDosW9CV2dv
z8XDfvXBvv2W1X+rD5fP/vksKna/UeTYImYbhlZKPZ+iGUUUiFkIf8yPOOPNhKXD
O7OynqImCCQM3AEBfnxzxF1JsmBve4fOJB4reQPGUyZd7zFo+qlUbpWSIUCZY+86
1Ja+Zdzr/IHY940aHcPcXL1/SJyYbojnnoFwJobam52T5aFGxea+Ku1AnzuA2Nud
6lCMUB2BjujCUgxwofmN96pRFkzYrsldGYbdRRnRGOKejkWVtAPGppU33M9+7nlO
iWxJf9ggOdtIcPOMUMkbhc5CJKBF9AhGwshcNa/fjgUts+O2VHWgGzU5TUC1BipZ
6CoCOxCiVwq7z/B8NhKW7nE+WixNWw4a6fumprWEMncNBxTD5rLWYZmvsfrcE/T2
2D8TJ5as44ZMCyyyuLvEFtXs4ombbMa2MGKpK/SUzWIAqEVMSMGu9FrZuRxX5c7+
vLWwlilG53Slln6sa7BsBj2/rCAuDeawWCsQyLLjxqJ9h/+KuVkFJJ9j5zjz90xX
yOwHknHL95Yh65isuqtA/GPhRld+bD5s4+jrechxmt1mEJ0P10t5DTX2yudR7FgA
1eA1mcpIbem/ljdjmrm5C9JOHZY+c3vZb1AnmGWqY2V01/stVrNm3L/EEjMlhUc0
fpLpgobLgUu8GWjG1GHZ4cYigVChlrFgHV/hkS2yHgIer38zVe3zxX9L57ApKd5s
rD4NQABJu0TlOc362swmxrToVWseXtrdCc0M6MkWKpb1LvLHzL76ecg7aqnU4Mq9
cY5oPAXKyAq/34MSMrbLThd7+I4bg+Mdnm95tUgeewOFdb3bf+5WF4xhds8ciXVz
I4cKlm+mreTmAciu3oV+KqRMN9fSfEf92yA6+ZwFw1qRMIIDW6xykHnWUxw32P80
FvqBXk+BwHeBTjf64IsXA/OExLtUdwWl9L+ZQ/W9i3sO3jg1y0TFAJkY+xnHduI9
2FVh5K511XSt9poEuwcWHGk43kwbhVmyzXY9Yg3flwgrgmGXGNro8N8CzLyQwZTw
Khmp71WBGJC8TlHqAz6FNb2Nl/6RXLXIoYaHeERStabVx3r5WzCRpt5ZTPY3if5+
1dhSSf15ceEeYmRJpC3cv8J6Ce+PPvuiSfUneKYQVs5WO/0rBUGzASH89jtyn/NU
g3fdPUl+oPlOQNIMIIGdZgACMv2C8ZKCnCotljrKbxQYJZbUXLsYIaiB887RXRbC
qLLP1q9DkdJPU7Rl9Oomh1s5fPgl9kLoXAfBnpHRuJAyD6oMlby9SZvvTKU9usUv
DgHCd498T+k9nJTqrNeKKkpU7W440EVsbLSUmx/JfzXz3Sn+GqmdW7ffwl4KUH6/
7924zQlMMkF+fFrFaijcIKHS0D4EQvI0B9k839rg3FYNQzfg4w/AgkLcxJK/cKtc
/QIC6kqcineSvI+OkKhGyB5Of2zP7u2WGxXQZJODFo/q/VFEyAKAxUGRrBW/akVn
rs+CKTDM9ogtQl2QBY89llLLAMh0yDEedG7JjlfdIIyQ603bY4kaH5kUgTHo2SjP
6qaByH43RIVpckCZBEI6oN+K0XiNl1YVYaD1UCQwYGsNKlN6IXUfAvTO6xAFiwSb
iNhrFE9NGAo7/CSusaFonE2hWyFXQ2/cBb8pGB2AexbgC4idSHGKv2SpDHZXu8Sd
1JYtnGzk2SsGBS451pI9U6Zr3tzDUIfV2fZSf3KaqFB0XmPGIpZxYgxNI0wtKtKd
93V1f1iREeR+iVCjxI+BYgusaM28UImp3QD4cl/LcfiLEepheYg7gr4QtqJggxe+
UTxCx8DKeXOVjZVPQIB7SB0KihKXemqKqJcPETdLi+PHmFcmxQ7fo5FCgw7Awo3K
emhCyO21177hD4rNXqU+vU5YOwYw28NZl4SMKIuSxuCE3Fsiq4bEmE5BPgp6+Krv
I0Szvf79SEh1mKBouWLt3jbSU2BYEw78meVduL5HEN8eIiWQCcRFcmLoqf9TCwna
h+dqKxND+JPtcu5vi+HGqEZauZk/5gAVRCdpl6CsC9fat1KRA3dmeR1MZMLek/F9
fbo3T9FwNIfAH82UrReuvvduAReAnzshjmIpjT7FMixhbVaT1CFLBV6NYoDOe/bw
Jlxenoo+M2gqamzY5cZ0LU9XIds+vxprWsHn85UT+uxc1Wx0LqLjOWwfXZ10F38b
JkvxAo4w6cXo9yqpt9DGv+FmBbBUBQ8ay/bCaX1VINtLHx5vS7YTf64DBui0K+Z6
GDSHhEFr6rZ3ikVFy6akfDAcU70gH5VhJYb6pm60686Cbz2njzj4Sf5Ad4pjfjoS
fYairMcs1lFXAsneH9c1eOrI6Y7TG2Z1fVKCmAl6fSvyrEOt15fYwbjK4O/8fuaC
JWgZuIKNeNTOqww53y0fj2xBxxnJBmPwoQnYvhc8H+zH4pgMS6rNLXKTg2yizN2h
5EBv1DCkHTqAnA2IkH5cttPLUjm8xe46d2qmQ0X1BOjpYJKEVRzO/VrFullF2xIK
ZP4zGTE/RGpL1U25zK6t4YVgpvmwi5eSnNZ46fBUHaYN8YZwG+rQRRFOyX8bjZHf
Sn3vBXDJqKFIsaxyfiJdr4IQfjljDGjX45FxUTDpTCFTkKM0aDVFr6O/2NtxctqU
THbr+mQEo7qNPk7N8zASuOK5DrRTGF5BKl48tO+1QrZV7a+r/4ZY8qFlE+62iTTw
JTMFC9murTwAuA4T0L5Jwwc9PN4DfB475WA7Ta2vt1jgp4iwc9vPk8vx0PVVPnML
0a7RHfwjTmTklPKUcdzVG+GPVL27HJIpi0YY7bRCp9os+L7m3xpK/c5d5gcdH9Md
YwkK/D1p6ESTLiFq+uyPgjCslIwIIIxblL9yK/StOvp+SzloiN/TCNLq1p5yM5kt
oODW2/u5UydtDNOjA8nr1VxlmhpRv3evIYl/xRqhiG0NUHjOkg8P+2PLVSiVkF12
DZ866qT+mBIdNFP9N9sNEfbrsETYT2YjnDCqNmcskFo6xpAitwt7CE5ZRacwtkxU
QvEmWyKdBpx+cflvBGsUnEkFy2DIjyKzpKI/aK+vRLv9oxS/C9qWv5XhUq5HekLY
esv9GFuzCkbPr+zvAOtviHHz+fSLdxhVloqNRLFTUHqPmv0pcgkU51p8+k2lOoQl
Vxqa+vdVW1ADik7+7xtiY47sJY+2QrDYlO0N6CGnU9RlJWh9pEOkxDAFdnDlKjL3
a1RN8gQg05i/V4ByXmOSzRWdwRgR/5ZJVhN7bKDGnSTjUsFxvnQr7JGNd4xe1/12
tEDALPiXlqDLPiC+HFdyIHp2QzN0ePUL44l3KQsKCvbhMJ+rOWSzWnPSSSYZFdAq
284w9s3R+bRKMzyaUDPpP1yv4bV3Pjxnze9V49COP9AbgIpT7jopriruNq8joE+w
Spm8JFYy+d4AjKl5ZIZBwPtYjeefp9TBsanDF7po0dGf80U0HJYG7eIvDcHibT68
R8joGtv6iNH/+JbIacJC9rERxFhzLPXVuthTDLf5ocZ+nENMqlJx2j3xPiFZlvbu
hyViIlKj3diQg0iLhgq1RM5IkC/DzfqcEpNak+0KdmfVTwSiz5D6K/2KWw9+NKf4
92ddJy68yWQl8cb5GX+QvegExyHvQpsRJaWKmrXUiOH693Fh9ZnYaw0Ry6eSL3n4
skEJUo5q6zZMn2M1+FZM5Kohj796eG1FiQPopBcPS55MkVopziU+RaaD/v6drlr5
pd2eaGJ43cFIiUAUAHmHPxnFFMaOu8IE3xIq4ZN7nr3Z/lrTT5oh02GtqO15ZIME
eGqqE6bDlnNCxdPyUODkUBGeixyUrwUgKYvyDvA4efOSHocPcUBU/kQNFIVn9f5f
hjREoWi/iNmW3luvIDtoBb7Wp+rMUpYVew8eQAn5tFhqRV+zHchA4+bwug0q4t6w
3munsbOYjuJ6WtVpT7zrjU5oIY14uxA9jxWNzG60igM1KHAkhz7MjoGnvqOzket4
ITlo0p9Hy5fBHtMlCCjSwKwQyXhmMBzRGos6asDND8A4+VIofSQ5ACIIZq/v4nFh
GUhxSJe6NJyBcAShvdLyoIpOq374kaRoLUrX00RaO6YoFK6swpUTl6GmuwOWNJpN
7Wh9O1p9BttwDtAKT9+rYDd4hvUaamNnCY2YaHrbfL+k+RwoUZxlSoxfwvPWrBNf
uvLLix+sLQKKXvfuGjqYT7+NuvXM84VjQRvfJdaWjyU966abDvd/kkNw5w7Egipr
dDP7JszsHJTPKzQLlP1WXJ4NOgzE8MqW5lDFoftgYqJmHaf70Y+Al6CDmdlsfz7D
8Tg9gAWQXhcX9qvB+ERjljN7uNurZgz2fKUXHlMSInvDi3UMMLHNHddlToeRgo5L
WjGR6ceM44NKZkndfPMER9nXLWNDw7agyWRzN+toZjNK4g2C4xUefaNFJiYvfo5Q
Rre/CvKswnShR4flYBsOoJBmrDuKLF38iHiqtTgoYObSPdWGP/r9M4I57mnzFJpb
y0dH9pTUp8M7GKB0LKv1TliCZysrCpzYeXtKOf16jOvm7eyj7wBq8SIf60otbd6L
8NiRoxW/PCMsw6tDbRbGdDa6xXL9ViChIyXv2sEqmfHXzn5IdlP7w+/FblzDRS7z
1vsaCWPKXDxROqcSDczOd9zuszNiHeakFwNyeMAbEig6OKoRQi2jBgU/5Gh28500
ZnTR5LMJxjYNCwqE5zjF3StOmrciCtYbeULKFQ5UgSSVcJwjkfTuHT3poH1UWIcx
2Q4dt6jV49lmoVXPmAGqknyJVD4jDDYggatfweHFDDsmHMnHAigbsp6TWtyyCuXG
w5umDxdZyuLw3zdU8HOPrq7WSvFfeBBffZAVdmy11kAYUlluFcSj+gnkPxI4o4P+
UUy7OYs5srQwmJzFioZmoGV+aB2EEjlEUExAuNTgiWEHNf1Qf1ogSYWovBCJty4F
OMJbnAHQBxFXO488OjZfoa3wY2i3B35Heqy3oQuE3JIQURWcGahNECuCpOl2HQgT
mDztzrIs9He96xfBBhAb8/sAZxmK7XXVmM9Gx8JYs+1AvI/iUGIcyo+D5S+aANtX
doP0LnFVIUP9r/zDudk82gmQvXZdViWIeeKJs/6mpAj6a8w/UPzIRNQDcrxv3WY0
2dSb5gl/Ga1mC7fjGHJlI+rqX+x0mGhP9/iUC/ZjQSUMRQ5l9WU1AytZC5CWdCmg
Mr7Hf0ryUZIwBKKuMeVrBZj1PvNr8cMLVzTbc6A1bXvMIdVGS9ii1OXbeRDa/Tys
qIAFj1CbHI8fTy+H7Bf9ZwrO9MRqjgejZGbxwVWt2eFWcLNgMsxFW09U5bCjjzmB
/MHBMV8hUPvBfZCqtVpdJq/cTgXPT35GcILkeRb9KSviZrwnXq7LBcknKYnNQJ1T
XTfjU2BXCBW8Z16uBlCaMnWAaTfenaKUDYMIwpbszkByChg2rd+lUcPwxaOfoWi/
XMXVrj2efMHFaUjfstN+VsMHCdVfWwpcFx+eiRUh6Bh7QQ/KL6HxUc9gZX31KhEH
fOlx9dgD9jv3lZjJ4/jz8j14PVR0++2fKBbRxb6VP1WoMreScj0p3eZiKXRs5AqK
Aamx4FedKXiBMkXpgVP3pgwEB9cuK0a8bY1M4oA7v5sDuo1pdL/RF9xtpGQjhm0k
buSXFtAeGLzAVTBKKxxLpg==
`pragma protect end_protected
