// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WRsI1/ski6gaKmoxha4CNnwTJAH1eH9gO0+7grGixm7Te0eNaJp6KBANG4r3Ao7q
+UNDbUMD/rQj9T/uguN2J094DrWct4BhNaCYQsyHAw4UJj8Sh5FuZ0pQMdwZyibV
ZQ6nvwh8rtjkhheqMKq8rXX9e8AO+t48L9rKUJtxMm4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46656)
K5IpVt7XY7fMB67Iu0WPcEgufa9qoRmyJ4vYZ74uhMBCkAIMuU0tH7MPZeHbfX2n
MxCmg8TK0b3omFa9T2gUciijqwHIXYhwdFJmdIu1rXAod2UFr1i6EbkyfeSGrdFr
nTbn5/8bQDy00qnYqg9GqkynBSGgNKzVjvUNZszuiRMAHSXpOl5didm3v9YjRtwE
UbUkm2vih505EVziZHmqwLy39a4nmBEzGXEoYT6cjzBXT3bs0yvV4lJJUX2AS2TT
xjfeOYZjt0yMGhTS2F5YjwJ8LW99PKNq0yeRERqSyfCFEW98ldLwAVl2WIqiQ2F/
jVZL8dU1m55np6qXiFg+G/OyhrthpxP4kJBp2kJpGuwsbY2D2PX6ccqiRYfSzHvQ
+mPI1O9rZ7/xL/5G2fYIrM2DplqC/+3UkUD1famP7vPyZRyEFJmjl/WHuRCA1cgu
pzUoRfK+nAza+9lm1k0lJb6H0nvbrcTrJdWa9PWYevLMWnuNTosO8/92kymGLTIk
cXawFUnaMLggtJRqJVDhC8eeUk4KItved59P9EtbYvX01Ib4vk6IbK8WskDZ7re7
P59oYqpuuPwUnDu9fn0oyas6jTb81Zyq38iKsQq1p1AeWa1iTY9sWzhEf/gRyF91
JJjiGnoJSMeT8UgtYsQwHmIceKjcBUUZiJewh2JhzvzgtMnqi7ZzEONRHJ85njlt
f0RjpTXCHkI1yxSFYZbaqSdZj6Dfq1lIa/QqSRrKOLZbvvv+I+O3Bd/ENAAcmcvy
/cvu32QavgXYD38Lbpv/FOykfbTxyIwj0hw5gkz3NyXpVoIL9pp+R1xKFWNoQLHE
4tQfGTSxLjXozdS9vAbt16rVUPWpSeujfo98CE/RxIaHkXXDy3bG3Mj7AN/uYvkp
l7DtzbtM+VdZRVJOl7YBMSk+7yNGBupDGrhX6ib9F9weiq00X+9c67cK1hCfqwX0
WBzO1VqA9vj9UerkkXUU4qAuApHsDB6QZDa+4naEEnH2Dg6rWtshQxNRxATtITbc
FgpYPps3L+WygfrsdJctrlCQbZYeCm00UOBy/mbtJdRyeXvBuy2uOUCwyATuJ8cW
Oak5h1oMg+ged0B7qNtnPCYQBdPR5soQ8GsAulNlWKWU3g24bpt/0U6aZoddPTGz
k66a3oe6OHDF1dTUlFb7n8LMoAzEL4q+N2tk3lQXAgNp66YeyyDuM+iR2Q+K4Kj/
yF7FoYtHEdPzQGqOJNBaUSv2soPymXfuxl3cG/ZIO5WNlKGMk7gYIMobhUSe/iRx
/LJLiIZvigyQk7C2Re0aIhw8AqKWp0ErY503aG0aSqabM4nVM8AyO80PbiHixBll
Yq8Py7Wy/fD0AXtI5mEQfb5MIJLuUc2v828BrHrxhtzIgAw7k3+UvTWqCbQZ5Ylu
ZbLHaZV8R0tYe7m/VFTp683iCLKDUiIQqjU/K1OM9uGeu/kyYWPruRDbKsvhAidX
5TLX3GZcmMbqNjNCbf/HEAzjr8mugPstCFdHHMs3qnOFpaEfSQf0wdm66Je21Nin
PEgbEkeI3NbqgpY1DvVVNZjoEl4GV5mcmg7/eyYOL5vGzUYC0i6dr3GrCrx85Ad5
CblqrnTwgaQyxXw4QWlpCMd1G8ZHClCUWDmT5W9xHnAFzSSqaFwCTuYv8kbVX0jU
KI5m7BrJuyaiqLXun5h/oXEbzJ4Eo+A/ia65nrtgdQLAG+G/8E06McauzZNMXCb3
XGM9ZtX9qeYEqas9isXJDhUzM7hsdC+PxKhZpCMOi/2Q7fcXJX2/TerrhUgPjOOl
AbXJ17L1jkl5Xr8FenFIPzept1y3ZaroleBRTSyBy9YpMmnpXWWiA7uYmnAGpd3a
06A6rK70YvYI4lEV3I1srCb7xMGijJzLxdVc0HOHwSRXQwLhafWhMdEdlQW1frL8
pTYP5bCricrPLEh/rGLRi75f90O1Sik9vvAWGj/WxOcRDxVn2PhqgJM/QQmFj+Sm
8ZF0HEIdeaUHk8IGwT8rCnReDAlYNRy57UhEDzZAM/uTdigOC0f1HUAZPyr3AYaA
2oP5Ck4IXDR5u2GR8SirNC4yWUEaRx91ruNwi8Uz0vNjQsnpPQlPpg4f8kLot5mR
C3juoBP/TPM/RqEuUAAnARnR5AZIF+gJRYUBqpgQLDz6B+dMK5uluShm2suHV4xN
wtjTcxfLALPhivdpX49oDusaMaKBE6nbSWiPD4rSqxSEkKRjWerEEiUVRbRHkX/c
E910EdVP4+gctRyA90/dqWyE5bUoiheUdbydFvdGrrsuMV5EaoUy4D7ieAwL7q+A
5syuvZMaCxkEQnXs0P8mO4zZJyyLzCoVN4JAqWB5J09WKAQMAGGUe3QFiyRI9Nbj
wONICRJVV3LKcJWnDMixdk4yinqvhwSLUxICPR+yiK249ifu40k0VZVi4E8F+R8G
JlJ6gOIx/akJX0WoEbK+wsU0lQcTT8tpEFg1VOPbh5ql+chOw0zEKTq/QQl5T/xH
5qPSCdN5Q6/RVF1k8FqluEREvFXXIYW6QO4Bb5w4RBXAePq1gUvazWzhijbGoAHK
c7OuB+bfvWUck9Y7qSHrEkQ+tVR95K9DdcNR50PSIzV/Gvjf6NYDHBZ6ZOCwiOHy
pileIj24VnbKOzSdXpyd5nPwr/E8jUtHK0t8TxgKVaPPTwwjUWP6sz4XpMnJBp3j
DYT4uiqpPUcneJWMzZwf86EB0V6OMClhikHEe9tG6YsZu89srxiJCrCPBIEOF8Sn
POjkL98kudlxzkf6J7AdwzBrsrh9RfRvZHNunZ40+Ys1Iip5OvTkUUqL5NWxhIMp
0DLtA0oYJNhwlHQiu7Dio+5gMPSI4L8xrVGi/HR46CTJWytDjzjjbPY7qnBFIQ4P
pcDBzG+kvTznOhrdrXxxYZY+9JbPoheYbRK6xS1GAeophxNfHsFWhcNPVa51RwLb
tma9Y/jBylaZRHdqcNHfCIYpHX3OD9DGh+9bOqrNBpd31JyUW4mi6JKRdnhLm5GJ
Y47Cr/XphF3gBKgRwZMH4IZAWHme+R/SqZ71+xl8dcbR/5UKLfZJ66HDOy9p2L9C
qPxl56tCWBzX7gh4m7KskA1MRnl8/EbqL3xz2Z0T12hvqX/2Na4I2t4CwCdT1wwp
9ddpIv2ZjWbOECOGM9ZJCjXvusBiAeFhqdmMz65YLMtQoIKOGUCFHyLSsmYFuD3i
MwOM5d/Jlb6HRyUrSTx/NOWDhgKjFrLyAPtD/KERowdeNrK5X9o8i4Uq26BEgiwN
nlDNK0ZTXYQ+H2KW7HptIYE75AGhNfQEZ9dR6iPb+V9AGAq0FaLI4T/tAz4Zixy6
MHV8UZozwgLHJMACiXl5lGfloBFHiqtfO0ZCSKa3gVNB907esJcG41hqPnTglW0D
yDMl+/WA8cs0MdRPMZhU9n4ncpGYhi6bRW1648CkuP7J7Pur6mEk3PHPSYfN6vu9
xpoMEzH+4+VmJ+JXkOw/ygPv+BrPkPEnkSy2mu/+LyEqJujGN3r9yQYFi2t40T2e
amdcPccg03UXOvsrd/AMo1+AXolpJz4IWGGp0z7/qy9Fee08rWx6G+3ApC9tDy/U
XKLZ+7T0cJZ3bAj4kxGfNT07+fch5Glay2Tg4Lik53spEy4jxQtaNV9m+1CUQuEL
OWHjSai3KE0QNXkcOiGGkP991hcDKaougfMo71kRfqg8gsRUREPK5N3uKJgXntE2
AWza/Xa4NI3cyfdsRsa7qzcdm/HAAAr5Gx3UKLxEzgmvYeiCHZ6OonhbSz7etYh7
4bEcwQfc+4R0DP5/9cjWLaBQysqRGva3NJsJq5gwaxOXTmJI8sPx8tdoiVENE8bl
HkyVroDxMdb2tiVTR0yE5sbdQc7P1wKYV6KzfRT0czqaCrSHk3R3j55ZaFWA/o/y
RvpHNAhZp+8key8rtipbCaXZAGXTbYCTiDJmU4+xXT3V8aKc5mBTGiolOhUCepWB
hu+BG402SH9VWaXnVxO0MOCjNTBB7gPGXoEn6VB0+zLZfXdyXkHyBfFz6QYmV9xo
2HYUE7QZbvUkL2IPPMmrOLg/zkadt4rKj3FK7R2oMWZWTcLpYMSn1eEILHzzE9tj
baJHeWLiLPpm/Kee7xPTJ4bBeurZ6qWwIS4QpsHQHflOr2jryPxMXOovKABzFytw
N1BxGWj33TZAKw8YOX/pVX20xji0vxE1q9Mm7hqwVBvkv92LrCnf+m+uI0Ylu9vj
Y7HnHHejc8MBkRJqi5f+pU7m9CTDXarsbB41FdX59GvBK3e9X2aq8/UygrxmtxnT
1M2u6F5Thxs6TflBLNzpRffVekgRRdRgQUKFeuiX4O2ycOSUewR5ZhQGeQqfFyM2
IIHzzjtSry5Yok68BOdX6cTSNmioZPVFZ0aN5SeGDLnWq9VBlJfwmLNnqmgqoPKW
yzUpkr1p12T3vYi9FWQFE2qe45TWuRa7db22qdJZjomzmFmuM8AHTEzBjGlmpuLY
yezK8tR0COuTjeIHT8AlEGl5NZXjc5vi79QopKFN++/gQlS/eifbh/xdbQgGRvJu
sAk6R5Rom0g4e/UTc2HEHHJJDnBjhjr0L5vKMaqnvg8ok5VZerS+J4cVSk3mCWPX
KsLdGXBYaMIO3jDZaDwLmhJ/mWk0J0gOenHjzsP/BdR/G4GOzss1Jz4LkeCk14Pd
wWS14P2t+5gIQjqGvD/nVQr4wq5E6wz5mkouLCgg0WOIo8avDzlHuSaMMXSfF5pW
1C2a5pCsqzRVLOif1RTEzh64CIYLrr/7YMsafedxN2V7en8rBPgnTl+T8mNK7p55
18VW5X/JJqN1cv/7aexMRRrvBVkizIZmQGRRV2rK3cspHerlX30r6LTg13HXI3d0
GF0cbZIyg7a+7oMBxL2nq+0dhw9K54sRnwbagNjSKsJoAZVIOYKcSfUscm1/c2hR
oKQTyLliTBfIspgIdqmgrW8/RNKEzMw9cBVmcBMDrhGIaq82Lek5PIXtzH21v/MR
IkDhqTcvYvJ2iESMVfJIWSTDbXv16x8fTvev40Koq0GiaEZ5rUaCz/cKoaSJJ2jC
leMEDkJlbVPUKMdABjPBKE+ANg/A73fnQqLiduy3HsmSAqMq3tlvG3QorQp29/Fy
FixTkXfXnTMxppHruficmwSHYKptmtDSDlzT8OdHqFdAH22NQtfOBsFXu+zX7+L4
EBsHh5YBTkKw+1YSVHD/HRotoQym2Qb6oeWx5ATMYdEZcssBQCqPkeX92wgXgSYQ
AJLD1JWezI3XHY424TKBsJO8B+YsPsPTf5NVsb2P10Pwsl/MY7SxFefBhWHaagQN
mpS3fC1btHdHHnWaF8nEgitR0xyumiqIFO/p3KMllD97ovjkceuiVfjKE8jEbWjn
NEPi0XB+iL67fZ8esJWOhj1OH3UoomYNkaEcRxOGdnWP+QYodWXUKqIosWTg3We5
Oyn87ReAi3VTkmGQ3rFfveA8WaolCGKbmZmHJ99n/3DT7RyP/b8tox6AU48BNr6J
8WL8tydGt3ijW6Np/bify4fMukqMpMH/wgJaJqM6BAEIfYvnr3YxF7mBtx5AcRfV
rpoIVI9d7dM+43Y2+/wNQbGAj8/7BeJqegBlhUVurEI5bFzOfqfEFhMUy4Oim+7r
fp5AtcTrg/8cfIpYwrfBq+F/R7e/t6ViNKRkfPOlq77g/G6N51JwnzgkauD658bl
48gcDXTQzjiSc3SK0SfKbyvCCpNKXsZLOjds2r0WnIHW3i8hRO641QeasWdWofvn
5Vig1xhOGWzDiUi/i9U0eV8mqjxRxVpsQSh7nDrlNYGRxXRMuNnsdY8rXXEcUMfH
2rhKYJdJPucz6cbGUJBtdLlbf9kZG5bQZVfkqaSLW/Psemt5Sfg8W6st7Y47Ny/i
/muUHDbZd5er7yZ28+YnO01htvuIylQT/9OEH2gD7+TKLFZHHFf5Ru0diVfraYiU
PgRhJsimG4lrZ7vr030VKmP9zByUoUbFndcMhakg8Sh+PgQMK6/OVoNiWvkRrW+u
lj23On5mVz7FUNxu6lvQjeLxpOvq6VIU5Y9j5Yihc92LmgFRwXB2Lli/jXg86KFY
/jzYXts3Kn6eJD3/j3FwqPGjxGMJKyDO8E81AyALmdwurnffebByrBMl2iL/iK5M
gbkixiSY5bY/KmjyzvISlpXsEJXVX9YTTgnW/GhdJsflKEO6BXChtV7qavwNU+rs
X/YNuZdCOjPKcsg1PGE0KrGh9zv773rTPT31qBOsp/eX9lFaeM57DuZQtFV68S0l
dCYh15ehKmIb6FbOsmH7WWhRQfO2v/o+iviMX4KMXulHSqTgd3wGdlON4PY4fCTM
OhVnUd6S594JhOTU5py9+GxBV+SJmVXOAQvIHrJuqgpY+SIX269Pvb9+FfLL6mgC
PwiKFpwglcmBDXpEBnUvNqrJp0wbDk72k1s5QTIPtD1rseI32cHVUJxOCk2u9qre
5ZBwLqIDP6PW9RRvuo6+hYyd3GfmwqW4ThPKUbIW8/eZcsQLjfpUoUkHBhQTyVVd
m2dWF4wILPAYI/UIo0Gc4qmTdBhLsOkAytgDOH5yCOOfC5tiSRcf54I8bU2OEzji
zajyFuG8E6ngluT4OvB7vJSrnvH7ijTdcGzAw1aC2MMVh2kzKtJrLrXYW/g8MD94
BiL7pjyYzCWC6GW3v+K6tIG9JiesuwxFnUpadM7NVbVGrmsfMe5tPJ00aOpY0wUT
8SqL2cJseATymBE+Cw0a5F67/wcnixT6hiFnSzENkmgxMgkobWN0l0zoMiUvp0Xt
gakXj1I8q1UOT3XVPiwpER707DhPwqgxyusMgzOmnybKMBxC2Z4sjwxNYMEeCK1f
Q41+YW5XLZHRattsUPeWiPHsBMDr/rOnKYAcWSzL+zTGLtvErbDFz8/EfBSYF/4n
Ud2AwiWtxIeI2a8QOFdpZUjLefDfkSOx5KukyFQmQj6dYWXe5I9TGqoWwgw8ZZDs
K20Waa7xPeWpS2gI9UvoaFXLJlPQ8lnzwr2rypNndX/JcU9smzHCOYgtYaRERX77
Y0s5I3jQTcBnLaMYSJsK8DcdPgKe62Jcdx75v5u71i2RBgYxU+0PGA2se5qLIRH0
hrVqwlxbNGKgTQQQJyr8FVagkv+jQkfogno/uKCTC8ZDvQ5Cf8iKJTJrwFWMiHcE
zlrATfhTDRZ/h/kLi2ISR+H07MsxGBr/8eALASPCKwGuqs0/DLMPXyB9tk1+ryLc
lkstZ3wnWHbPAOmG0Nkxexbnp2srE/LJimaOzrYq8JuK/Cax4rbJgCZUQ1F1rorp
M2q4gUEzdakT8MEo2UeuPS2h+EN4QQ8l1u0bNE7noTzO/pazNk7uGGnKy6edzN5G
RViN2ckCyHCGnBFth9+N79gWOeRj/6MryG0S4qSZ7NGwDQXF0XGxIjjXsAlSpDoo
AzOlGAe7152OuLXTpdK78aHEG7tzbMyV/Im3Y5UbanvAmdt38gDklQZkA1Oi2Ftu
hmYITwCGhbl+gjhXBLaDXoy8aR5bejG8P33jtKcknVpTiWhshQv67FQwldMIOG8M
ztboTJ6sryIA5GK/Uh9UbZfXqw/AR4GpNSJZey/Ry96YmuFyki3lNaTNB/PG/PSM
XFkxAC9tuv8/2gcJTUn5lraiAko84Vm91Hw0p5P2wP6K+zhggtalIT7yE/6tHZsF
cKF51WzzgpYuU4C82jxCLg4Hz/M0R4MBrxqgVXR7tI2KTommn8pWLItUSp770nGz
cxg8cnFCgXyjVI+71j+6PZgtFSTdFGNZHAomaMz4LA+CZq0bZi+hERruJW4MbLy5
NJte87kUG8Jr6Bjq85kB/EBzYc3EtVD7LRbz2rRaJyM2TAb95HJTStdWWrtF6Qdb
MwIe0pNPLx5aHgECagD/JOIHeC2u0AMkQdDjMNvvpFwZGOf3cV79P2oAfl4L61XI
JFcAoE1lDFrbrPlkDK/daXxNSndhWXfsN/bmGn73I4QfLBK19Yd39e5XBya8fvME
9ESalumXfuqVEzwPoOlxm5p9PtNRaHZGmdsqtsSnQFF9/A+jw6AXaFbQm7tQVPm6
hm/LpG2mqVSqujvmm6xLSjFDFTf39rUPYNP9sMwhi3Ef268aVrnnFmeEmdKpg+bQ
k5LS6mRGyd5eQZbbU2qkjBM/hjm/r8WzD56HTUGi2+PXjCpcGAMGZyl1/zBfH66z
fLwAKFuXLkT3NfLLatuFGtmlgTUeuTcwgjr3x9pLa2eTSbAJqF+UR6Dwl1NCjWTp
ji0XoA/i/0rvJx7qdlf+zq0G2nbEKCw9+pvj3vNQtWVkldSyUfmtd71LLqPHPJ6J
4UVskZgL1Aj4eaxOyxwmekU32TOO8b8BfYMKVRYZXSlActyXpS2uVUZyXr9BRtBb
Gylw/GbrGq4tvajAzt5vxBCmB8Po5+soRIcrg9tWTl2WDdM+2slIfgskoQxVN625
bDiKPnskpE8SLQFIMyCUiOyFtGpQCrn9MIy726UgGSkv43sL8lQxP8G0f10XPBzM
RKgnwYYskDgLVuZcOU0dLR6ajdrS9ieHk71/9FO/NVRWCstxdamvihXNdz2TLT7P
vGnzqHJVdtxD2QcoGATHfLZ5xcTjp8Xp6DthcVx07UH6f5oiHXn0JFe01/4zt2Ap
K0IBhuKLu3MSpBI9SEKNYoJwT4dsJ7HoQqDv5h7u4zuvHQtCEDQvSD0ATZRNrzRi
6C0X798zcxEzQrfKs6JXZKTyKiudQ31ErIhpnIVcZz5iXf5AWlc6yt36wVabRVSk
MhpnuySBeaY2ErqO9k9y6osI5EtAS7lXbWTpV6Pm39ckac+I7gafvJuW8JTvLpTT
pk7kY/Zui4TYJNFwN8EzLfKXHOd1QBZF+lP6H8jWqpi4S99q+L/YlIJt8DB9aSbV
8Ch7OweapNC82A1SyTf089NeSAilEBr8VCnZy62KQWAGmlqxrQdz/LFtZCTqaRFa
o8ZuoczAoev6L7rIK6hnnlRl9OeC1m60rwVNQQU/KGIafp4U7AK6qzRl2QBfgUlQ
uycnpoeDmmPOgUVp1Y7tqbMRqSY5WKefJkIs9+yZ04ko4NnjVjT1UpwcxxuYQ1q5
oGN9iQYI/zYQc368TGPDLpfZgAn2pmi8f56LX2pNWOqMOaruEl1DxmBqOeJJxoJA
/NgGDNmFq92PAd5tveTziS9fbdQT0m/T24WPpvbJvIhAp6w1yFiM8dxyB/vTvOU0
SWm2eAaQrZXIuGHjgykTXozNYbbjgKtGqVn7vKXzkxktGFkWxbfQiQT1PABUQXlY
iw6c/71esEOCHb0VQZ1Iv2eBLznXhCsX5/iXcSmebHVomMru4+o72V6Cppoqyo20
b62vJrtmQvUiZ1pHvE3xwKAqSO2kuaG92LyARNiUzP9vrGobGvT+qGmlCAZjGe07
apU1UZBogiQ62sRhuAY7nYQbV7M4TSaaS/7r+s5sya7p8exTujvZ5uPPgqmO3zPd
xUa7dnnqauP8WUcZUmV4NPl/5QAjTq0ftgiFNP4uD+SS4jgqCOHKGMvEQAeKeEdp
Sns6NdyH9oJWowXAYIA18v5lShAikCZlxlprbbKgW3xQA7lytJh1+lSMnCIIYG+n
vC5eCg4DKq18qJBrL4WwxBwDT1AeA7DQmP2iBeh/wbiMB79FjC6NLY76Ue8kFJ80
L++ZUHr1P0Xz4q+W1SZfSbmSBQjII2Mas/FfNZiQSf6iM0q0USv7dYkOXNY9GvZh
qO05h0aQcvvYODJmCYy+xgSfRcbsRFxcZvtBvWZpNtPOWFbHWvd2imOAk6+VyLDg
oihznEGqC1sj2iTZC50W18jTfvscRAusMVpFre8EfAt0r2BUsnJDnxzPQ1ko1Jt0
uYBjnQ6NpM4ZLDG1qNxO4bVvNqlHGg7pjb2TeypjaWsynspGAW3b8ZsQd9nBgWks
86e/JInLaQmRvw6UG15gWk5PkY6RmibW7a77KToAw9cfGVOV05njAlsIqbGkZW9f
UMPlg3ntYEABBcWCsONhhBAa9ebuEbJrBGZtTAichpaZDEf9ttKTtO/83zFj9dVS
tY7XBgi3w7GumCX3gDIKrjBNCz8SALb49cvH00hhNWoBgSWWKRi4RCtovJtY8vCl
pY4w2reIVb2loqz9F/WiNaobloPWBhfJd+DMewdJrx+9XG7z4aRgfhKeB4tkl7ed
3un+Vxzh93cRR/zfXGX9f0wQ4hymJrdL8xznWUBuQuNuH2Ty/oHJvzGTriKVb9Xs
bgW1rEi0VfWegBz3/eIyv+YlSnUxO1MUY9i25jEXEgAOMWz3tWPuCBLui1v5i7r8
m27kO2zmXtiM1Izoto03nHkksXvbe6QJC7C7Cqu7fruo2qUt/5VGVLfhygEwAc38
t1xIuRGPwigLunYQ5pqcbLb+TyxUJcLMsBBdf1u+iYVfm21c1yUgs6vJj8aho6na
/iZumf+CfopJ2LgCOXhNEiPwJcV/NwmTrN9wPj9t+3uM7k3nIMdcQvTRzUfy4bJl
e98FC8DiYPvbYNESmufoY2kyQlJfEGSwml4KW51giGEVWKUC1pADsloDkoDL1T9T
IkepO2gFtUCogejSqeWzuJs5wsPzSnguM3/4IxVFPs3SqoI0uU5e7CybX8yCN6z+
bQ2SlMS8tb0XXJZrzsD5qJ8pxVS+4qL2AIh2G8KIv83CM7i4g4MjqaBYGpuotGsk
txHWxYgR2Vk7owWMcCnOe0i9NqmXZRehD+XGU9QRjBa/BR76Ihx0SvDIER6sDlNs
9Zw6Cheddg1JXeVSShZO+0duWx6PZD/tJpUK0OLsfksoBEhg0IL7PKuSfA2cdmc1
UB7EB/wa7AEf0YgmALOU1XLdNKxaGOMNusFNU0au9s9CGT9fQXwCMEK22D9a6F6X
Zghz+Di2RQMb7HqbBeEhXeYHiCQ1GF6cxl176k1sevISWR1+PLqGYILhsPbUbZMy
H5FHWau0SX7EjxxuYAWz1Mdf2jqPGWwqsY26k+LON9vj4s8yZQNaFMI1C7V3VNvv
7w6aKkiQ0ThUgnitYZXlHULtbljQhMG1bL+v0Zbn50DUYgBCaJHrjSaOLwNcNJtm
nYtZkmv2wt7Eta4OqBHHxD15WG+TynhzPztodbTmkBGmXU7QosOoc9uOa7s3K+5E
wJu7BAqjy5Op1UkieOY4dun3tfYA5kx/HspPxhz/pQLDEV4RyK6+fcLo9qFBVd4T
DSEvajgu0cuh2CPqU/haCou7JNUGVe7syBmMiNTVZ78MjrAiru2OaguOPSanSBrG
J/0PQ8swPUflfqybkYs8X2YJziC2fpdcR+nN1zIgJ6AubDjUbUGu4A6SmWFXCFP/
fc2cnVbNJ7jHVCALxXcCi9wSBu5MiAbhwGMwFllub4winFPEyM6qfJan+e5VopEK
6Y3Ff9xhVdS7wyeo9XsM8obwaePGDp7+a/sEm812v2VywV+/7pRdbcJhVJ43GeoO
3Z8LuYCjn6fsYh90onUVH4EuxB34DbLBWSQ7olefqF3OuI4d/HvNBEMIEb6btg+9
sqlSEos+4DSPxy7fKr6nSHMHPnF0y+ucsKqTin0GvplwprVYu4F+8KBhVzL5/YmL
ACR04eWu6wTkzXzKANEbYfjauaoMiKIgsuUP5yaVkcBYj3nWoovVVKsOChvShmLK
KquZBNMEIaCJklMAvtIIpeinTnf11M7I6uHP1mN5ouHSOFFs3254kRvAzSzyiMmD
Hk4jhQFSoYxK8L0YsuQO7a2Y0COFhRt4y959gUoYQGcJf1dXmTNrVV0iic+iUWi5
yiFWoVQgviKxVzPGukdSTHoEZGBJT7WBGTQXndGkqzualJpNr8SH5SmJdrSSsicK
kIpOZ9QsSgeCkKOdAn/0i8cAiBAQ2cHwkNdaCPESSeI3sq6RQr0FCpdowOiuHp3K
Iq7/4GSlS/49ylvcSUwOmT4q5PGINwtAOep5HUPi5SHWxRLK5eHac2467pLk2DU6
XIV+Rl7WQf/q6P8w92WwRoFibsM6ot6Tin2Woi2ViB9B4rQJuaHGqsNtyJIocrk/
l+x0IqSjgryE11vNUYR/dNlv90uQQ8KVKj0Ird/UY4ZRsmVcVCToi8UPFiB0Afsv
fCLjKPPr4fomUBP6tOocNWKZfdcsl7I0n/AC8HgURD/Y0LC3ARfJjKJime47BCvI
1TC9cCUSW2mcarB6ClrwIm4vULahzE6BLuDAell3V0huYoNhNtSvvTerNzslUOUq
We8ZZvvmws9l43x+UxdeciGai7u70TyKrv7aIcBNl6QikXMdkWRYPiNCqENy0fMD
ufcIZagDiKGnwgu7aNQ1Kg85ruZ0kAPP3wi3IZagDaA7cOXGLv01VJUPRn/58nd7
GBIhlVnpKastj7Sfl2r02PxJSFIx83a1y/by7CZ/W3IqZlzm+vlq//X/lzVkowA9
UKj/bOctzX3f/clZaOXTZeFT8T+4vMViTbIT74omw0hhdNvziL/iqSOPTrwOa40Y
n+6qx2lY33E83pSd6a8EzqeIsGRxX7aHWqyS1Ab6lDixTfmQK4wHv0X/oO6lHR9o
3ZcQjUJk/5G+ZFcpQa+khikgfl/r2tdNzX7Neyk0LL1p9ZrGo9NoZcj9HRobOywr
Q5kwgHYGlqLXxJsHylEkNZu5hkVbyxEpHuzRW5vmVcfvCzFnv0meS2ntqMuSkk1N
jI90sClRxE7THe+js49HrIosLL4WjAMo2Gzev7DomztGhZoeqnUTCXAbCE+fB52L
Mk0djELiHYCKrpUn0u67k5eXls3Qw7ucq9GMBdITGDFV+wBZHipgNzqL+fNMF89W
Dw9WmZhkDg+6FNkb1igKAW6A55wlL2kZ5cK+zTPcbKD4ZjogJHSSsD19cPbxZKer
SJApOsmoDYzlP6iuMPrcbEAnZ5ZtSIgLdV2q0G3hj1Fp8o/IefIX9UOqSdDcDVq1
lSTsrtYzIb8Uq22Th+rKVOXo71xNU5INId8T+He6tqFCuU1ek/Y8xyEsf1C5SpDX
Do3suSJLRH9ykd76F5y7H+BWE3hTC7OB10o0p0VQf53diZhZtdvizieRWvvUCbqm
qbfxR8oZaMY4TPT17BBiamVm7DxokdMfsczznGatPgMpIBOwy31v/bOhXTc9gdAK
TV11bVIfjCV8b3lUEH4IynZ/mn2FVYU8Rx09/CJbypqJkgD5gRrQfRs6TwpUtbqt
Ur+Uoqf09u0As79i2hNtbfIsD/4d8U/9rwXBRv6002FJ+OAevSZNLG0OsLdUTVvP
C6a1MiiqgWOtl7hij01b/kSdeLXQEbQX/g5Fjv8Uyzm48z5r0e8ydIEc8AY7IAjQ
KsA+lnX0y9KYWDAL/x+PpNusrvngzsfSHf7vERUp/o2c+VsQAC1Xeb3JujigPf5Z
8KHuZk9gjsxWYK0JT+UxYdrdRnzmnSc8xyayB/qqjUGkpdYpgl7r7Ah1FWFDM++M
cfZxb1wmTTNXxapwC9N5tYVd/KrEDew1KqdWZwRZ14geHhL3+FDw37VsdQtLpK+V
VjY1iKPPejgSOMe+pu0JmE7GZ8jyH2BVL35E2yff8FXtadaTSfoED3OdzYrqhL3/
JC9FBe9Pf9YdMvGa6fVqrrxwy+yxmQPDgmRvtdflypNz5sN+AStp3iAQwKtoenkb
x5JzYQ+qkrVO9pRINx0zvGhF/SqMPLSbdcNYTAH3dknzNhdi6KYZrbDwPpGBGNmM
xMx9x/D/TvEpMH9BfmzwCOU1XP6Jjkf4B+MxA278G3P/ED74/DuZ6RZ9QiJTauqt
flDaV5VmVGdvbB7CbwxK3X1zqBsNSTOpyBaaVsYwQ9UAC+e+U9/eYDpbthspUUpt
Evufya+RiPrcNOY5yRt5d2IwnpEKvEOH2ylEGrK0X8wDoCPFk1+2DwU+DS+HYXB8
OUU0huvze7Pm4Oci1FfBtlF29Q0k5kuMcwVqYnYfZp7U5EWptbWuq8VDkalNXN1b
9Ui/pAemsz+uZTqybAtTjLdkqyb3ok7CB7CN+zAMwtJDIilbt9jny3XDi9Hj5O4H
6hGWbjYMLBm/MGuYLM0nImybnO52KWPY72oEUkAyaBur3oTmF22+oWV1oXfbun4y
Tv5tf6lCtxCHyKJ91zrAhHXe5xm2pkiqMTPx5sizJdo9RNnp1ab9i326Tk10MFBK
uvcDQbORxlgpW6Hi86xtFSIFNI6V/laD7gbA4ph/PTv7piFBf1f/VDQhUALOsYA0
sU+64/8mYlKzue5WbZK+bOrYve5zeTFaNPusYOgNfcqRfZ+dKAreAqFkYlssd8tK
W+do29IuDTshO4ePXtGKTix9TfIOCKoLx4eAXGrYNf9z9RTEytEzsr58r9qmpTtg
AVLoKLgLaQV4CqTgW6dB9XCZaa/ZjTF4+zTHzMkdWOHk8Fuu6I40hAlkCwothyvq
7g0cT20JJtTqlEZnKANRoo+oiRvg7k438E8g7YQaTx4rWZt+aw0i0sH7CYVuXCDn
98LpYCVEXAexn5VqA9adb4H9C6ON7w3EBY0eR4poQ2lVpIN0ukbXTHN/gSUgGUPk
FVo6v4pvZc9pkg9Bg5yOI0+MjVRSknRZsUkKvlzEZ4yLApD+pUAUMMnlRGnczr7F
0IBANxZrx+MxGjv9/eTIRBc+B4cYqMgOvOksXVPrQctvFDY/8RodBVSbQqpWhMXp
GvuZkyRFr7RGuWD8ZEgUziPLRJvIQK+CdlhHeX4I2cPUXh8iO/mJQoNCuy5jg9Wq
/webB+IT5lbitQeyKX27aFbbV7Q4EppBE5Vyy1T34O/urcKGJGuWVlE6isb9UZhZ
DrE+sQmE5ORAU8iDlBJ8ShsCxBs1YO3x1c1nXBB4O5FmXFrXFgV4LYJGdbqtDQ8v
A7HWUfmHLkahFFS59hukKn0isEXmqbbqVUkyC3A3/G4o5XeOYoehivEmsN0Llz0k
y4X9GtP+twXH0rfmvKT8bNVGJsr+loEsboCDspHJUcwVSCQp74ir2RsU6cjocYEF
rm9kH/p7nv3rwSJYcskZdkrQoaes2nfZuEMUS44mY9p4Vds9x4yqU3IXV/090Py4
SDygoajDrujbFV1S+tfI7kgQOjY2E/h8YFL4Z1d3Ps62k9wCNhZRKVW5Xhl3dqVU
URx/Pk37ocHPbBaaH70LSO222ybMkinCHPUGNqe4GFZ16Kq7Ytu3CFJyOtxkc2J1
fAQufX6IkHcVlzlYYZRh8glvim5wfw/fDJ/PmgxO1LO5kfujQFyHBWhj582nRYJw
IaTC9zk5ZE2Mh3zjmj4wZwq5RSGKB0jKNATmRZyjE6rRO7TRognS6TZuhXOa4n+b
cchxVZ98duRu43aYd1ABig1GsfJHGT8G6o25hrl1cLIZUcUfXyWALy++tSH0wFGi
RTnqdu71WqIcBiM7X0Grq7I14DJNgGmYoVxPOxaey5ZyNGNAnyWL320xZFTFY5ee
2eAelOHwDJpXIt+nnnFASwnARyztf3bDOpkfJJTgHCywvbMoOOeAcz7GrgIJfIPX
GK/X2AmSTHdBmA4YT7ZsKfXqPSj0Bb8CL0WT71lrf3UCrmS3Wtu2ozUcQgg0B7cH
rqhq1mC+2Hc1bk6FAykYaBAFTjfNRwULq4SAK1k+MKWSDWuSyyY8kL3iTgC6tvwc
NQ8NTziQI4EMsmTbnHI2c0+iDupbpnG3mYBxZh/mJ+xB+vWX0l4OTaJulXFPG82a
YJm+vrlpPddAD1jMxVYqNgMDDkmDMBiCQQ4aWIhvhpwJkTDD3mEiww07qTuGQRGN
b4TFjksdnRKRTwtqD9tXcaJukGVJK5ZOMCnhTEX5X9WgTBiQrQSOgqn4zXgewia/
jGQ0ajigGxniDCUWk0AzvymEuepIrLC0nzT/noc/Ut/kfQlhKvw2aBDenX4y31LS
BYWSnQC3jAi+kwJDjTdnKMh6lQ1gRr4R6X5pXomxTSJW2IzO+kDTfwSDOm0h62jK
djJFA9QfNTyUU4kV/E53ek/viDWBJgJSqAYiki1PqebUGMRB0oA0JPmdMHj9NP9m
aOSyAU/hAk7769apbStYxNlZ/jakkGOzAFLDtbwNSyDdff5XNHIEyYJL7HqopUoR
Yw/FG6sUpkPTkCWYks2PVzz6fk8yDxKzRLgBB85qsl4PbV9uIzwuIKHdwm/cOBxX
oq+C2MGRWjFjgnYZclrKCvZc7+Dds1HbAoxvS0JTi6uS/EyMgSyTl+t3ghaqMrR2
tzeZfKfDU4miF9311gHBfX+TfOKCYsgN8uDMrWwFJ+lhGmunIY7VkmB3bQD409o+
6wI03urpPkNPeWUFqnY1MV4NkV0A9Kg1sqNz3I5uzNOurjnpZbButnXwOSI2tssL
NTR4iHWtMx/Nbk6XvPTa1nB8Jawqn3e/i6b9jCCqX1Pocnzn70FCUocvs1849nID
CKmjCIWrk3GDzKIcjgZYK/lo6t2Iz/uEdslXF1AOAYnTiG2HUPSF/jRl2DyBtBJ4
4icOcsR3grbWBtt32n1xuygzfqdq+g+K+nJAYxdZ1ZnuyiMEFUrJhEtBE1AIqmMF
9e2GrpnG6dfBesWL/iM7fPhIjDmm6XAzw+7ChAD+uQ1iE5VT7cY5quqzgWJFlWJ9
DvgFcbduCywnheBnE3/iTl1CVFZsqSrg71qGVOGOEed9wSoneD1hyhmunwYEmR2x
/Db51Awn1hdXAMWx69M7OIgXe9km6L07zkNUlTKzOlM+j+mr5EHekSUQW7wDbOtp
cUUcDHbTawQIyymWQbhIgT5UtuanWJQsS3+Ce28RBcA1929KSeOkBt7Ztt02N51A
wuq9kTGBU9tijicIWRacu4J5CvNPf89A6DMco7N2MHQA8dIU8QNgQlNgZ6/K9l5s
gh8WqQxlbiCWl9oBxg2PyDphZhfk9x19K0ARJGOeejKMyXLpuz1+Y/m9XbJG0+Mj
c8Zyus6aK+2w/iJ6d4vYmJ/509S8sH17ZrY+A3YpErI8f4rpNN6/znScjKzHeiXD
jnoRlmCEQ0/pGVc4Ea/MiqX8FNHvQIN5PXNj11EvQZvqI4IOZVOrMaOuIKi46tQp
fJ643u9tkQ8VOgpFvTyND/c7PsRUYSaZ8pFV5HMB/as6MHqX7wFcdU0Q1ZfbiSqb
JsfjHjOk1IHLs5C/mfoNBbGkBl4yMId7+OJa+PKROA26Hgmlj6pJSpPQBNwgnYXj
hbVNsqsFUM8YNaOXPk/LrNNfJb4eN0jduvyvtIeM1tDLCW0COhnhPXqOil1pMJiO
Dl6RcY22fEjo41c4dQammVhzKfCFjHK+85j6/Ijqb77LrDZ7B/ORIOI2+Z9dreNv
khYSlYkcCnsZvB7j5WN0yrO76qEy1dAudKw+ZPvNMeJQJ+gyX/oxjqk+biiFvO9L
zcRuWqvALneManvAnk26Ze4tG4krRBuiwSgpXYqfy/jfrA9rzdnvTmKYvSAOZrHV
1c1MuiVfq6zbiHQV3A9hlG7tananLrZdl6GueExFrZD6f6Puh9RungRqD1xmD7cw
H8MQTU5O6pXNhGQQCldbTeMnFeywLPQelIxA96GMCbTMdvWyufLqK6nW2x0RcM5a
j2XHgCpqeZgDnfO5r1XGiMhp6kTM2eKs0BN29quq5qAFj64I/yyIGF1fWXXXxvy3
hSl+it7vGrc/5wfGqsDKb0vaCX3cFjF6GC2WI9ylZv+oS7zva3JMAaCXJBoPKifJ
Dku9Jwuq41hnVeMfdXQ1yAWRRKWYO8k620xX3+wGe3fXEh7VcUmayjVYkkqK6nra
aOo2fmE6WZwPvhuyYOZlRytq7UE9vNwRf8kkF7ot3+Sdu34dfemTxnFOfzpzWaBo
s0lKrPzMcFVV6CWUSXK3wF8hiBXNtD+sDzuTwkETwqKhXam5l8PNr+8fjpxMoGYs
q8U0x51GhoEBaNxq81dJUd0teRHNG71AMuEDDcEqE6z4Bai1mUCCm7fY7RfPKx9y
xx1ytNJFCTIxAnBU0YdXfZxZUPhzekexkKW+P1OS3zxW7kIfVG64NP/KYdv+TYvT
OCcMJerDwID791GAM3uLJqHian8wnOCROAh5b8pssP0dBymfTkbNHSG4tIdZ+CFD
c2bymrIC7lmaMaYSb6f100zX2/Y/smfCUuhHdOWTcSxuG/hAhMG39h7UN3Pa5rvx
tJsH3eoOroNRfJ0RUlDWPZtFW97EOg/iXGMjCbsn83gZgRMLiAoC1FXWf/Squ97g
FsnGdd85syPQsTPzDefys01FUqB3q1+8jCjmZ+QEsBRFw0sXG39L+OpbFGU1Z5jR
B8qE4dyjPptKpdGuEYp9SBpo4dJQT1cJPW+pzQVuB3EgX5g8sFOOZOLQFjAHRq7g
ObtgB3NshbyjSoBE6IBL5HG9z6wbPcKIOd/pz7+grpi+jGvLHuarY3j2vomynkc+
MnT2iRrGcFBzRTf+GvzonYi/ytJAf7+l3nYOUjd9ntmOJaB6ndFSVL/nBquZdTkV
VH8L/Opqz3uKP+SriDYTH+8lHgG45q7K4qyznX3UyjtdG8kvtC8nvyS1wnLvcFKK
GTFMzKDJjmhnQHPrAiwCI0ho8P/AvXvhb6N5lZFTs/BAdI6Qdopxj5AqmtJN09E6
McCvFANv3FAWSVpXmhOKi/w9rIRiYMeQkKzH6kiv30vTTZ38BhFx5i2o/7j/X14o
jb9D+Aajtv8qq4KLBIgIXFqH3a3V+VeNjTALKOfTFt6L7unJVYN6F5i4uUkrDcEQ
9RVAS/lpckdiq/+30C0yUNeqQjFuAjCKYmn7QnoNnmAH1scoeKuWkzZkceFaFmYB
btZA21wX0f4AvlGsx993Lcxxz3YgBLp5fYELmZQlwghlodu/lsMuBJ5VNAtrtrth
Vh39EYhoUmVeWbXpYWPNmv/Z/ZdzV4kKUEoIwzc18PXpy7sVY+/xp95srociKTSY
DhqH0jwf1M2i1myQlgvgIpUPY0NLGNQOn7avFIS6V121OjxB3hjGWLW7jWJAG6PP
MOj2TRSdeGUCxtgpGFidk2XeKnKJQbDt2O9KKzudMAXPSIfHF288NxdD7OZSQbTQ
znGt3na6HUHDoaM2Z7yliH1N41lO+mmWotClaCUMHGTDxOee3kpKbY7ga0Qn4P9b
9kKFsMyv96J6WYMlfetGMFX5r9CACQD1UB+r69b7E6qOPfOWmCb4FyU4S1G6OnCX
ZajgA/Ygem39noRHINtiuO4gxSIHRkcWeechu4N+O9lzdc0g3bVDFiNithWRDD18
R9oKjHD0FI3LrFjbFnhgfH96NN/2RrUh8TA18NxtCPeB+V+hmpDO+ZnRAU6bX12p
xeInJntDkGsF/74YXMPe3Ly/G37xr3tHmQQQ96uzqKc9P5sCAxY14gnhxBYyuPIA
RsLxEa6/FGBKdp6VwxN06hsZw0Qj0ZzpzFE6mmEAmWl3qV9E0vVAyoTYgkAw6IvG
e9xhqPEgv186nX28IsXZSqFj5H2oFU1+8+8aQHACEaQDURm8Q7q2E6pyPJtwwid2
S4pVwhHxiAnBkuzJ2/4pxUkWtKmRe09IkT5qzg+qgufQNogqk7azB07KL5PpoWWV
lHM/0m+ZyaUziDta6fWhw+sNRQhCiPOXvmIaYtfKzmKA7ExYSjZEwoq7ZUN5ombI
Hr216sO+VZtJkg/apdst1lm/kOC2lrnN3V1jseOi33+nFOf9OGQVdtF4i1GtXcUe
NQ1XKM6R9bdKBRtYQMfeUuMJ87W1EKntLVgoiJkrpCcD9YEe5ar5fdnuH48hIVSY
mtv430VPVvGZpmlYDGoip51o61AD/fZKTDMcGonFylTQAEY266dUyWgQaLsXJ7lW
SlKuBzN792r0Hn7JVl89pRpUywh+lTmLmzBxD/6//1ViOY9PFsNnAGoUDBpG/ILd
IgTlDwm1CEEfw+Z1Ej9Lo371IOyUsslGcVD50s5BqpyGtONAEh2GTqdMY8wKPdQn
YUIBHXtO8KVg/1rGP1hawrRnME2nvJO15E+iy3jEKp+CY1nSEchwfA4SKpcSKT8Z
lyEu12ZUEXBRiFw3B+jxzRwJexNd0i30bsUHOylTREYOiMQxMX01nGehwkqaZ+c9
DlMdTPnQYbCswwkNFI5rXT55/+Zi7ZUoaGmXPwNHzdaWut2Env3m9ymb7d2w7/QI
XmzuXVrr2vILCe1fuASerr0J+A6LM42PFf/5yXTzVGS/1qXvpvASGkL9/bVJGJKU
nYPw80fDViXYUPm+yMDuzWhegTnepyEZToKg0RlVoNWpY2DuMXPTx9EGQ5zO54sw
36j8Yfvwap1Z07LNwuUCquqhiaM4i7y0FZiDNudFhxCo39KgczdwnUChiFOpZq6B
bvx1qVNrAgHOAhVQo7MgdYzN0b+w+8Skk3YNwdkcs9+TIwh2Jw4zFcp8ob0Xgc52
NSNKBZRj6cT4MDdmm2C/WGIxHIIvvEX6Qc+kdNmSnkn8hyQebMoVMzh816Yq+ixh
WU59Iz53Poz1y1YSsfrS9gAE3zwiOVJQPCXI5jpdpBC7tuKctNLkhWb6+w8ED098
AC+3jjsc8RPBaQS0/CRg5Kl4Sz8ZipVK/R7ta2NGKlOUG3ZChIR1hV8KU8TIv4YJ
S3S1jjS4QI2SmTp7Y6Y2rPUxW5p60Ne2CTf5ZEhN4idNmpybgs1JZjAie/ZFcnS1
tpULGNcubabUfKAENWdDo7w0ogMhWaV20Dj6jTN9xpCaz31utqjYoQm61uqfX10v
82V4bNsq1e5wJrw9kjXlKrcnsOMHpAfvWdJ8a8IRBidtWl7layNxZM1IQ/jJOn+o
O/P6hHgyuY8NSyhNt87UAzIfPhM5DUXSI+uVqEgK3T7yu4vfkEO0l2KZcGcZQ3Qj
vv2VfmkvEVZzfDnhGCCIQ2YpVTUFw6/g51sKZpacdm1HqH5bh0T/Qrt8LS5VtVEp
/3jOzt6/rY8v1irUTag5n6jPrGbj0ovjfGmMvfLytdPvlVux1hAWhlIGuZLWXfuC
rNgVXRXqyAciVJChS1IBryE/N7pF8diI/5PupE9rn6bpj0NQxC0Wi8D3vZfJm0do
RJ3rWebUGUmucIF+3HCdgWFMPbaVsUJwwTxnxVs+dk2uMzryC+8lRroOvUJDJFRL
cPq3oSIbc9WQ8hLPwn0v+uDiuSvUdanGUSvcY5ts7HcYgu6im/ytI+LOyxRJV2Qg
GifNkrUDsIXuUV+ilOm5ULvWbMVOVD4nM+BHKMFagCkwR14IWxUFB134TOV0+9zg
jR+n59NDx76zMb/G/O/PyYitT2iyL/w11VGxVGuFpzM+1kQv+IybTW+ES8afUn+h
5RjTm6ewIbzgM5GWZevmCGlQHxbb1rJtuygecdsvtcdH75jjwzaU2hCALuyTLzok
XmfLEATXMs565NO4oknc4HhqlalWqA/ljDvMACCzSObtuLIOH0uBxRcRji5XsIr+
xeD+kiZqQutLCFIyozugfIanHZs1hfpYQbKF9UttgQTIiMY/49F3GReCsCu1L7jk
4lUMD7WD3b+gVF1QoPmdi6e6+NGqN7fRD/yqsDeUN7lHP3fz5r1BRdf+DWKGk1Gs
J0TDp4HD1OqIl3pfcUmRAlds8sVhaPjwfGRrmI2StDCX+f4rZsTHAKLWeBVAepBB
BZHvej17SEc45R4xtIZ6rGhQ2sKaS3IvpL1NbYKuh3JiY0HFtIPRhI6ZxIfeRC8+
XNLY1fmg0+XO1E+cazHPPD3oODiMAMKTqcwU1nMlANcb7bsicMKJFms1puKnPu0t
YsRWbeO1/7TyXJ/G6nwT2HIUvpUrHJuSqPoWuJ8PXS41R9HUfyqAjefJa3VNF9D4
kTWME1T/Ho4EGGtyKM47eJO0Xy65ccPsrGtJfwuGEiS8FrUJSP9C78plVgbck6Un
j6l/MY1znln0flyR55LcNoAL7eFcjr2lAWY6rePXMgmvTK9u+IL/cZjjEfEAeQgq
MN90cJ8nAmogNYF35J8z0WDbXB1jMZtISV03bU1Wtrw8mBQnBQf0pOlRffTSPUTF
4WVSJIhW2ppx0N7q2atVHIBNn0rmCpy6kcqaIaS8OOAHBdeQpnoSiAM8o+rMo+lX
WTX/V9vUC0fHU9Hx+86yZU4feNkJnQOVuRRV6/YfkLsQ5rr/XuSJCYSRKh1GQf8y
QnzEq8pVtlszkGziD2cLNRJBKHCWGuEq0Zd2mauTND7V7TeZnxo4GyVrsHCg8T8k
byx41KXP62JkNI5zC7ZjxQlWVisRyrqMlvOYQ6RoWKF7FEtrK8T5DKx6CZOiFfEv
MvAl4OhRap+ODvS5f1m/Pu/mWUcx2IERaq+mPZ/OhrTajYzUt8BUjUJrZGcpV1BO
eqVA1nWuWwyWmoHWQsBXNZd56hnTDE+I1XmmgkC9Nh5WmC4s0Ym40Q1vW8oFGg2a
rXUPDSy4X8xWP9M3SCGcTVQGZ6VSb1JJNzzE+7g/KQ5A5w7vuIxjE1gJpZT6roJo
h7d5j12lCg+XpIB2a+mWj13AW1RJW9i0zSArIDOK1wxO1XzdX88a1C1WBObiM2qP
OvH47OrevDKj9XfyP5g2OqtjN50ufJsb7t2pMs5mfQe0lpqhbk+VkyfkHVuqI3QD
FcCiFJqrNUdEhUe9Q7vvaIPlCHqVBX/4aT4yPiKaxZ30GExPo2/kcZRQZdg7N/su
xjn3/vX5XBv1uVApIx6diMcwcIRXQH7MXOtgkXhDVkU/l6D5883wxBDrBPfm5ox1
pm4TqV1AeYUMJ6zr/xpEC6gGPCNtjwh9+3pUIa5t+F5AwKtfliby9WwLLu8+/APO
KCxUSlRy+ptcpStKRDpElJJmsRYF9hzSZAEG8XzjmNOpNJwrs6MgxKTCI2sMeKD2
6uoc+hscocqiatwdFtAzjgt2xxuk+WxDBtgYAFAmQ5iLQ4ZGnPnFLEoyZIcGnVDc
OYnh9kP96DLNacuE7tbeIYmyMrGtF+041DoYqOj5g7cV0MIb09ebyjS0iKSg4abU
vXcay1wOc+pvA4weneSh7gZHz1BNEIzFbHSzfyV8pRP1XAlorhmnKfaR1TdREnrm
ctESMISGg4l8ZkC36dr37a6gwr7RUmG+gSABALk00Y9+iDr+wz/2/99odBM7eN4f
a4NoZFFfdD2YP6tbGRd1RciHXdWdIbFsQ6nGNIkjso8hCwSSwHON4jXiDHDCw1mI
RHT2k63pmPOmevPQAVHTAaWa09FyXqzYuk9969lxezPrpSruvdpCcO7qJViIFYBT
AFCBIqoiZKpO/P/jT546cKhDxeelLM4RRvGqo4I506yfLV0kyY3wymR/uivwHb2x
wTmakze7q+A68vFrzhvZ1450KCX3MY6A+bXHWsrLUnbTOS3lUk8I/ZW/Vm1mWGca
8llVsyztXM7A6uT2OpGqK+5k4AY1Ks9GV+NondUp3yc+GtspizN8T1CkEAjW5c80
tLYaMKt3Lq1QHhu90sKanxMDYrW7Wr66L99ilCl8ueOu79xMKyLgkhhLbS+U3IYB
h6mDCNTkyLqumkQculPXRsHIADonYTvShwUONPXsbU6TUnh6tDWvLSGDro/a0+7B
VO0Y0zJCMxG8RXkSK81IZs7XG7TN56UnTMCI4CvsDBVf4NGzroU+GLLfORJiAOyv
1p3qmeEwWaOC9BQ8DXoiBMnLRbL/SdaxImvrWkUGdqOhpWjH2u/oIlujQvLmzL3S
CkVb3F72BIEbOEn7gjRF00cwRW6OugvQ3QShQPshoV2MrPb+z1iju33KOapYtu8u
AZ1qmkTvwPf7q6OojRaHxvBa9fbGsJ1tvQbCqD5COnQg70WyjQemLZf5o6ZboRh7
u9HUVv+H4N7/7UJreTx2mzxzyhdDzLHqKOY5bKMO+0y1p2/wKjxicWyD/Si5gEkk
SH04xdhh5WDRKdRtDPYSSSmbZg0xTAWQcmgL3R3BlDfwuUZ8icR+Hen1KmGXqqEq
8/068HiITQYk44lmFuGnvbGiMkLtk6cOKAvlGpbSiUBSlnf4kCo73kM1EMxGRdJy
ZYZOQmYAA7cJ6bvYp+IKAF/M6oasYMvG7rcqiGsoX2etkMkpKtM1QQk4hL0Ix4NO
urcIyO7V3Rb9ai2TlHKcle4xv//vIhZhvnS2b73XYL+AbH3Z+/Ay3/Ewb0NpiM92
l3HLMfHARmpy0TmKzaP8Fr4Nf1j2RphDBd3e9+YpSeXs8mD6hj8hLTcBmmXnEBCV
9OcUHUWX9aeWuWUOlIXgbz9TJYcCt4l+USxKanA7N4BWW7SwjmTBXvVGJq9wbfoO
O9s0/TYAIywGOSihLw2A69KX9QgT57jBKDuReQKlHVmclL7lwCOJPmzA2Xtq4RDT
pbP9Hy3yTe8+GHhT8tT9tbbpKLm2Bq3w7U2ZpzCgbZxjFx4b7lfLZfTBZvNqGyj6
P6SOOWH2Fqr55CBOPD3sLLPFf+Jn/Ub8prBvD9Xuw0V0ziNVMCQlYBXg39v+fL7Y
410o2f4xgYp4AgT6dwQGbAqXNhmjK0kliTQ/Kz03bLhBqYoK7sST5VlsM4T/7Xvm
P6rw69W54aEIMiAqmDAy4QyKX2noOBHTkkhX13WmUMqwBQKth3BP0A93RRYYR0Aa
4Yp4Xwxxeq8zmfDZXetHgj1CZ+KxhYAqAyZR31Bsh/KkNGAUI8pmXpH5AwbEF+6h
VIYXhzzpPLVLPAhNcs4PXDXWFnK6e5rjHf31+67Xf/5AIrO1cZfBEA4kMe7A75NS
0FmMkhuoYT9qTwbBYrzZR6E3q2ogDDX5ALeEGWpM4cquYFdCz24mUAXY2Js9Bngp
XTLnkAPd1ZqoOt9v3m368HMsrpA2xjn3x4zVsUdDbbn0mVdd1PMqNceY+dpeAJ32
b2sevCQ9nsbVq5EtgV4UbKGZyc/Fdsw0uXCpF7Hfuze6Ezng0517QeGWSx9xAYcO
6lk3TYVGTJ2IDpgbAw65xKDXia1MtVxvM0lHIcCQkeP5hk6yD7NUrUrw9+apf9S7
NISPR0Wq4S12RseCTfDxyel3rpQ4azJULLw+oVVmnnYzasnWtg/2j+zkJYBwcSDy
kUS1y9ygNu1lh1VrjmGpjfE4q72muJzPhoFTD2Tvsy+Q1F1yfQBd8iHGgeIzuQvJ
QkLfNBWC9+p4196Sn6h6juyTQuqYg2nKXg+wD/hpbbUh8A+OlLZfyDRTRy3MkYN8
J4Ilfi7Ura3530kCKDq2PCcJtKva7Xy7XCmM3GmkkhGFG3nk/0xmKPlA5DudixS/
o9R5hS3wa5LPRyG9mZTbu6037UPI9lGXKcnfAKSHWoPCSxWdntLrahMaUvhXSHGj
LxriV9LRr37K9FEwBYJKs9rnxohx7H6HLroVJpSq+7FdKL397XcYbacbULFa/h08
h/n8CXz+c+2M44SD8yAFcz1dptYffx7lmVoaSf+Xt10nn4EBkBBv5hJEHXeQmb+N
aqe+sbGthqf4SseKcqhltr9yyR+WhU57fEXLmCUAV9MUJrkEMm27jD8yxbkA2yOn
A2xOrUHxuOTDwU2KobHBN6ivc/PEf0oGzStonKt72S9jqLnKrVrnuCIMty5SN0Ek
CknmtQoAXUlBLOQlxOOVLtP70X/aZcH8L1LAhHWjBThz1vBCAgm3Ofgl7/9KHers
ajUSTHtBsNpMfVb2mKfQd7KAn3Czsxcf2hPKpRck4b1kLq7XTPdTbab2ScGb2Tgp
DJbX6gR6cSWjaheiy9Ip+iBNkL+EPtjSFY0QtVCWRhPlcWAXG1NOQYAfVsle9L6O
JTVWF1gW1/+zrnY7ssoPI0NikjR71sZFrtpeFTbXEJGRsbFAGPv2u8LP0sGkqEAz
s4OM7pGuFhB08EetLTIftfBNcvm6b+5o6n/8CDl7tEsy3NvWEvSqEaNqGCPyP2tD
Q16rBC+dTMuFpxhrTJ/bno1tVuZR2/fW+z67k8l51XkonLNXQIow20i4XYNhxrRF
qZOji6ooDk0iYgcN5XprrTmb6M+yW/wy9YYtxm6arU8rEs13AYUAIakXQ3jQzfKW
X5CkJtPM/G6QFl04MpAEQyWeaXdsh6dgEkr8vRo/FNEq/HaeKuz+ZwG7DEMKSrMy
3E+lvNVlYq5FcG5DXIu8Rb9PwKWbC7jldEBYIWukm6vQkuezp/NlWaI/03Rl+jRK
SUI/4KTEJ7PlhnpF6ai8tfT2jm9wtl9jb8OGejx4Z9VIAAWihyFPVgbgu5/CNiEH
f12An5xVGGeO5D5IrGiVHkTja0lQWuSm27mPkOy/9kfG5fhmMsq1QuUl1n3lxtW5
/VdEvbhMQUJy96L1lS0/2H+uecImg8E5Zy8U8QbqNnyoGDODiYkqAEfqeKJCN3es
v6zkmKYd2cZxM9fPk0VVTr1kLkG3LlSVVchvAirkdP8+st9BnsPVE2pDoZvZwBMd
RoNHl3kEpklZ5fT16YuvzenXiLJFAun0tHD6bO9f7/n+VmeOVsAR7xjYZDNkNkgV
X6zzkrC8QtsQy0AoVPSVXOouxK+OGf/5wGY37PD9Kg9TBRM2Jqfdld3SBpuYDBMt
Ep7Va2bYu0z7hcyAuDNVKOmSFJyLGD57emyx1HawLAXYBQNpyu4jHO854yajH6bl
oua5nPChLx23oFquPL8eIrdDGsfUltZYzOlWusihT2n/i6jZJ2vOOslLaIWiQu93
rBInGvokZRPjppgUlS4KMs18CmCw4I7i88Hwhy+JJCAMYgaEGDFG2AbzSdyCdsOP
chGefltZd1TgeOsKpj+fgcF9lM/hpXCySaAKk20keNPqB54W/8123gSvMwCc2au6
M2lT7C7e905be75J2E6SpOTJN5Bv1Kxzc7IyqysXrXNeBBwaQRN811Lq2LinKZF2
TmHlmv+thfOK+TDoAJDHGHyXYoNRx+K4srWipRWo0W3xDd3gFAixEb6qSkG46KXi
uW+lcBigorCrgIipYe4zeEzzrptszCuGdFbgJ36Up/o1gVYzZ6pjb2nmE/VHSEk6
LULAXika/I/amvV9KihrHU0CtD8zuwochHGQi9Zn8/+DkS6MTazHgYGFPqD5aGr9
HpeVbNM8YFhF9GdOIiPajqAAEORPQ3pMaVRKwAzXMJjrANjZ9mAtHujui9P03SWp
MgObU5QIDGZGji9DaGEJTM6xepZyEy/58Brkeet7SyRQCvBm6rmaCNBZOKBkO/RW
wy/idpfoFgEzV6u90J1hPQ3HIgNSdRcvu7PR+HaQq7THEdgI9JOqcqY9oftHzJMe
3O8yBHt6B6eOy/B3c2FYPEE2l+jB70/W/FeSJg/UwbzQumsG56xcSn9WyE7FcgqS
bcvB4ctGk6AbsTVIwR4A5MwHkDDXpLIYfg+JW/0PatMR9CO2CCHl/k1M+dZwbMy9
v6qqjZztmpKc2PPiZe5yT/DhwzWE17OufbOhSicbJYpJpk07QYmBX1z7grFTWlGz
f+dxh3bt9k6Y+436Liy27czkJGM2YDv4hnIt5768gcccIkjTwReg22ePJFSdwyvV
62+tTf5Gm6eApPpQ6iWbDUi7rtwhduPdFpR9pyn4GaNbjgyDAMqjelH0akEG1Wxw
yLAqnoEPCUEjupolDJjDUMTI/q9+kBvy5mgoxbyCrX5Bql2xRF7kj/2rwWRE0sFU
BoRH4Du7KfiNAkZ/22zgK3+U+1kP1lueWk7K8EmFDucC4X3pycK10+KBUKTqwVYE
jycYlojHDjvr2ME0h7zox7mKYtDKwpXign/DH54fAPJ9UinuB+SSN0HMLX3JRSI/
8pjwrZezqX7tX6QqAYbH52rPxmNxqnC862OdVCc3AfTxE7N79v7cbm3dOYyUX6ng
7HaGvpXOiw7y4PV++kQtQBTVeHNJmla/SWB5ZilNTCiWPbFiaQ873IJfA18X1yIB
RoB9A2+N+f3P3fd9XaxEx9wSUXddYo/oL6xCf/X4ZBXDvpgMWcTXE0G6T7bDrhh4
HnDRYLX6Gk5H/byYT7wSUs3q45b0BQOfgQWu6Mc330Pv36CZEr9kFV4HPXIUiYjV
gg1AyM6r1QhcW3LM8k7UwsdIw53O1uIVrFkewuGXNDEj7V6wgefTlnja3QniOZHm
Zn3F2WhGVb3JmQuqglEnBhoaH/ziLuJ8fZArN/K8ZqovyTBdlIoqjuPyE+C8bgH4
PwwI880Ak006jKeyuBrpe9TNblUl3a1+i0WnGzpeBh3BoSU187DrXlG+6EmxOHK3
+m6dD+OVCOUTT0wKP2ioYEPDlUPHKhglcd3V6HSroCzSIvBZaNMqXt8ONaG2S7ON
YxgmJXBsp9ng0wwWkOETP7LI3r/25yScQ0/I+i+MHHqOl2sV9l1MBh1q8H63iSMZ
vVUyjXE1QTacJvqGDq1bwSlGBb3fVtMXfBKajZID/JvOdWaijE1OCoM9AS5wh4IP
boVxvAd6pj1fdFSIZK4VDrld5mGRSGHhyElubg1ZYWqKHWExpwSCB9FErA6pVOyI
RWC4K7ss0P6/LaS2W3jl7QyWg4QjZ5scObU7DDGbUs7/nXe5YW9SfxmnrHHzabj4
2RkcBrRE7kfvL1gJBAF3HHOoBSd9e46dS73UthDPxBmcGUCt8AFjQp9QG2ZaVWQI
LYSTXmbMgBxhGuppVIIClbz2S/p8DodmjNS7NOZr9Opbhq4iDl8+qlvIc9FpYHJ8
ikLZC1vcuWcdEd7KSUpEAoLr73VPOMhfXRAo3rxZZX3nK73VeFLAuNIthXwnGnug
tJSZSDsYHtFHcPNMHbJTxkMDrtxzBG2muLdyYUlhWXMJOH+9EVSwkWx2ylkcNl0g
GABTCzjuzkLfDEmbH95Mzr2m2RCcSBCXrihxN3XOYhRwz2byOyF753A27RZTE4uy
JQHXIhymcMno4iy9MTDtUEjc7QS8w0VHgBzNUFRBIz2kZq9XLEs8/nOFSluWxFDw
6IvSgXi6H4yzm3Qs05roXjUgadrklmnmUv20Cwu8sz7lAHZiMuhlDaYPObG4vjuB
5yfe14vnhYi7TNLBX/o69xU2LoQ+l1bSXIr1yg/7ooU2eTdPrgsw8tcBVK2tYdKe
yKRfmNAamsr6M8RLu5DZw+OcV6gami72dakMUG9JdOEFwQTJWvKPEWDI8uRfjJ5X
EA47sXrtyLa7yihbu5YCQDSUpVsFcY0d3sOTQA7NiLySO3KLHRcrzhjyrkbaSfFD
5PiWErW1I/b0xk9GTYQ0+cee8rlRFzkK+LdOX4mo3qA7sSSVKPEoBYXAISvfip/g
6hPva7xnuJJkS9cK7Re7RRPDYTVjqQsw47xQIOqW7b3CXssJ/EFrP6lR8mNCJD43
LQ6WDHzNBBDzRAL+1Ebz/UQIGBekn0jI+lYwReAz4hf3Tp47nI6EQMrRO1Vvih7Z
IK9x43if2FC6RfeHQCiVitcRwvTFMhMJQeB7tFkox9bPAs0RLPrJ8AXnzN3CMf+Q
9KiHTVuxCYC/KN5BtnEdenrvuZNFPkIH0qMTIsOwGHj0QlsNshvGGcVMDMjfAdnV
ARv31CwSpcwzRJCNyj+JqrbvzettwituAwVzXTbrpCBSErD0lk4DVVh79VMcJSNm
H8NwChjvMRqZYNeMLUe9tfE0muIwsxob8EzAnojRSHhcRCpAdc++QmnrSi5PvVao
z4ee0K6Oe1Xmm5bgsAgYU0JqRmjxxEB57/DRHtL9F4fp45wi9zYyP0r1PZHsOcd9
DwYs4z75oxHmvLoAqc35DK38uhcbTbtJu+7c3cEgh0vAkeLhzkoDgmTzJAbDHnLg
yr3Xr1FdweD5fiBTf7sC1pWI9hRRBMjlvjkumrKKCroIozZoEtyVaRorzMokhXTQ
GL0b6YCNmadeK16nkGDc8qYTGE6KN4APGzgVjI3nHmGGWxAI+fOnKIrf25Oywtne
Xd0eYRDOBcmOOsuxjgbtjY/FXYMm+AxnOFlZ2pYxwI5tB20VkuRudi7OTNTOTVqm
J2bxBlel/B/+8iv9URQxyy9alSzWact/LLLuwBRugK1msu3jfBE+Bpw+YbgFZczN
1/SJW8mAN+2eZqF5thV+WKJ5WPvKjsgcGI0DrVMItmYLsHOnj0SQaQPuAvMo2uKG
lmLwR+5SNE1ZRwMxJ9M2sAr5XkISY26DmLLsYApOnAHT9oBH+Q9CKCM3fD3Pm3wo
00zfJkrgWOhG28sySh9P7vjPPfs4cd9nXIO5fY/9zDpgoM+2b5GgMYkyxNCIDMkd
+wOtujyjHzROMbeLWUCuPFWQl9w8uuhA/1SfqU1ZOusZZZvBit5Kmnt8oZ84/Bki
KU00lFPNSDQVB3sYwW4Sm6xxq7CLDE+dcwCqk4QOoTeVJM/AoeQLMxtipEiuRRrk
DJ6OT4jJGvYw2HSYcLcTNOalmDQGHgDoJfJHWmIwXGEIP5jsYGaxkmOHWtMMIHoX
gPjn3BByF4DZJaFJR5PCyPo5Ica/RigPE0rwlJoLFYf9J8sj5mW8eygUzhrb01I7
f8zbAAKiJZkgsKlgvDUkLQLoeqLRb/XczhFv2v/XOEbRrIaKW2PeciXd4ZvmbrP6
uM+rnQnvXYcQzmAm2ZoKw6YqRcUQf6Q3JgDk2shmrAAFSm5jQN3ZxeWUi4cyRZwH
D66ejLH4znnzgbw6QowZeYwuVPx5afqooIqLMcNOGgnqtYejUW3vE7SfP9s2ZZdz
bcCumkzjhXccHKG6Dw6gEBYt0NWQtyGiZIDRQ8f/aWzAfU3RebWCUEGdk7dzyWfH
LqW+qDY40kxRcMa2x7nGokCeqcT9SPo6H5vmcY/S3c56Ze1j0Kb0lUeMYORzrLhf
scjIf1ZzCW9pX6GIYyb3/2C8bD9N8k711fZEsNSSvqqyf2FExN9ZokTgWqupTHNC
FF7LiXewIloWMDYa2YFNmycLbzrefcCK6sNjV94AQd2Y2zxQwtyqZCXj9kFi3dMs
PemAI1Wlms9DkrDr+xAdYeA2rQn+N7YvitzRkLPXXwNY7Qj9Hk+mezsI+7JOMRCP
9UunpceZV0LAQ1Qqgtn+WzW2nYv4XbS0tTlnFGPgPnAv1rniI1Ns084uCK1DBDBO
NZPLDc/vuni9YwwiZKwMZwcc17PmBphqggAVkvReca75NLCgcdrT55bOpwUNiMah
Qu2Nck/kQiqwY8i/WFPdBrdrjQYy2nDotgICsuDvZAzG9YbJTXhtFbjiVxON4dxo
RkjvHCZBeiv+te6asC/BzKx/72rM19ij1M+dzx6LWEi+v3cTYDir2u9Sk76jx5RG
yWQsvsFMCTsjWfRqaxFtZeWNq/w+YOThfApPsEJs2ZThkl1XRVa3zptgjodNxx1t
DO8Ps/YRDerXnlebPqv0jS2UQU8BMAriSoRjed+E52u2/vmFxEVc8KRkNMzZf8ko
QjJKawRVxQSfFhZ1tyA15bSXbs0nQ8FbjFWHmQxp49UQ5lPeVPO9+Pdu6G6fIFMr
bntCfoJN1Ll+XE0Irtq2k92NSGVJpW3qT4v5zcQY6w9DcJgdMDV2lyxdv4RjT1au
yj1vp1u6XNP203Dmu3cX0WAGMF/DZ5E+ShYWQsIWGMYv/YgcmnhqV3WqQI7fqaGM
v2fv/x2pDzslvhecG6Y0RePx+o3JsbMcHZqzEKv+vrNtvY0SK/eMI7tIwtE7Ikmk
kNzLwoiXHrkfUGztIkg/FRbR3cFCMLmBDnVTbBSD7ZpTcnH5fKekjzt4KGPr9XtL
I4jlRdvyLxSRapieRrnc4l75Evk9TkLOu7AMT5MNg43QNSGu2Vu4CEUpEgzjvW7J
m/ZwlXM0wlFFlscjFS+MEIkyqZaPEytq1izrF18BgtrBCKMFkXFk4VwfRJadN+Gc
XgRmxU4OJWuS07jSJgxCrawg1P23bzgo4F1MXQuXiZUJqLYKJr7POM1aNcy6Dr89
DadQA05tlAe7NWgbqpstnoNvoSWsBJGxbDRcKzcr6tdI+fDLQKI8DMNhfT39EU6D
WFQW9IAhKBnVufM/t8aHlb+65iUgX3+SJ8ac5deyh1ZDCh0pO3SPF/bKbv9/ywCN
e6gJkvXZKmO5SHcwa109F3VifdldBtuYKcFXtkYQag2xADJROvLrf/xDF7whBlNq
BPuQq0QZLSF5ZdC/0Am6emoCKsWhBNnWurGqvjXvJiorCsZj+fKBtwRtfdYtPf40
rqNvJFfq82wN2KfkU3vbV7PddVUoCq6dRYyk/BbIuMAdbsZuC8B8PsJKKxB6pkYT
KaCvcLAfGyfnhNFbnYIbb9U3EMhusm3ysCjv1Anh/tbZ0bH4AvFgPsrAJszo673i
kJjRYgHDtA+qgdUyS2rdD5aKZh5cdu3OzkJpMeye26whpqWUd6zZHQg/FDhZ7ujz
4f0DXQkONpRiejdCzinMczCMBpcIk3ZtrRBssEysiWLD4iZmWdjd576vX7Htp3Z2
lApPTcfb8jE4EybQaNh+kzg7rlPhUmOgjl75axdEp048mDPwKaWNxXE+6paetqFb
skDQModYiMHEPuJ+/SZ3P/jfNIVYF94KPMupfkagCqSm/D+ZJ+HtN7oEoCt+i47z
w6NErDvCSYUxRfJlIFCka7aWC6xvPrT/x7YmH++CSkYJ1X9Wpas5fbby5XI7syD2
Xtn9fKfM9WL3ojXM2pVkJU0AZ7DzOVCo5gV6m7QSe45Be+MzYkyzJy1VR59btoB9
e2icyDEsGcvp9v+Fr+uSvKvbIFVzZC6K7CdFu2z/iRA37EVVWocTDk962D5LwqIA
NHKxq5ve5XzzOQAMU9BnXo8wF8DYsR5xrKsNOQ3RyboUoYKkybqs0HDZU2GSiTbE
JnvbaNLI5gbHMo14xLdp71Mi0B8yTwgeAeuh160EAqSAss8q/bbtGrzv2IVv9kyR
CQMCIe9Hyy6XXU6lpqlrdf/aaheLWDGd6uVNvgjSy7Eu7ZIs0XBjo1L2qwEky2rq
mUcftkUVkvjmoH3paAoQ4jkLL2wmQfRieXHYzhPHrnF99qAY8RGnBmMnxMI14+uT
npZg1Bc034zh/MUIhdwFilrES+KuI2r6XhsDejNiSFO1VaHf/yRVj/SzyUKL9iRU
1S3DR/1/OAqCVmpxwa4PTvBlVym92fYHYylodk/57oHmWYBhlqC6Hla7ydCNqfUh
0jA9E9tmAhge84lKxQTUmpruJwQKfrjhYgGCns7OPTlKx/z+G0tOshT79nrczSjk
uiOyFErs9S1sLRNvla26O+jL3MOW2Jwj8HCW93qVp7GUqfPyEg5900P+a1JFNV+0
NRA2s/WlOwYd4HUVHScS0IPhuXUu/LDuuDtFTzy8gwf66da7aCX4fkaQoZm7Xyc6
DhFS3lhiU4rAKmgX5azcRybAWUANtaFLK9UaPwVcQSw+OUuZ9KGA41qrp4ZHkFwF
n+hcupDJyV9xUjXLO510E9bHukYrVdJje7kP204lhJZG6TY/bdCuht3CBI2/uOPe
uZzsooAnIUqAVj5eT3OJUw4qMZ9ZsjtpwxT1tRtosZ4opwsRG34XrbJdbmuxvsID
v60D+knENBZnytTY+EGUEKTFsPmmajNYo+4/moV8EPqNa05EPt+9hJAPXzOScp8x
BXudNekg6LhIJamYBkqrDgXnkLbf2vg6c1VxVOtyZCabqfZJQwadKZasr0lBA4Qq
vl5sKcQ8SbadTj/nB16aD6RXc59NYE9uojo0AMWhlxfWqQfp196O++kpmp1UZWTL
NatNNKB545MycWMXsE6XZex3JvvRKKpdgctS/XQxgV1V4FSrl6fmB95KyaKxmyAO
ZjNrlgLmQeCKHqp2HBz0tFeeZw7P/WZhLp/Wkt1bIz7HbCa3GVJUMenGARfkC/Dh
NF2R5ByD/SlWU3NZJPzUieCYxK5uEg1DNc5dGD3mR5Y48MuEq4p970CEZ/v80Qs1
YK+oF417BAre6z03UjJ205kuwQong/FtFbNe78/kM8e+XYEAxkiu3n0KKs3Q0fR9
HDY16TH5Y+n4HHl79FzZEz+LhQFqGATtPYtnCarkn3BXpF6UQw6nvF8ISihiU/Aa
MdjaRhXOmZu9F13QcT0rPsRgUW4WqapL7PKUxBnq3lrqSXSFvtKj+X9IBQ5yVJx/
31XXv2VbDdQ75twOx2LW8FJBLY3+jfvcmBSdLCa9oCgSanl7WxExVsqddKIEZqbu
ZniJMAShn15FSbf84xqF7aUYDX2+BaVYHk5Bk4hhar5aw9KPrrS2FLAo3ca2cULO
pip2rCtKZbU214WeDNYsgOAdMvf5JQ2mYbwDiCD3Ei/9Y4YqxeFzspUtKbqjvOWR
AucmdGjylzRoRJ898KzoS8Nnrs094pSog9Yd1veXaX/29UCSjTTuEcAATfT0hF6E
yNXenBxM/jTJS1hu5CqQ1YBxQUdpiGqfEY105EbW2GuWaBjEYVsNVvvdB41p+bx/
7ZwKztPKH7I0ykgqfe0gIMoj1EZzmSaYhvi4umQSaWWqMe3WXSb2im3EgZ6f/E8/
QxsOiZNIATVkwdAIzHHl3321YyH2NPq9NwYqJehFYOTEjzSsn8f9y5yLbX+KXrUo
WOiGjBt8VNo+lWipqCjsjm+3uf1zberd8tM0OZZ8Kjv4vURQwwTMnpVj+q8m5XNM
aw9FD+3KUr3C1EBAAEbxoKXrxm8RdddT9aaZqhkxPJ49oDlKj6q92eZBK4I/h8xH
DfxFtpRiUxnNwwP+T9enRzYaYJfaoirz3rGiQ05oqOJVmuTJwV9jQhvIsiPEkqJW
xtQy+nPYISerPQzaq8VlSkpBVbkeFAFkqC6zI27XXjhHCDak/NGlJge9+LkrrwSG
wp52HrBzw9AVUroD0sjC1n1yZ8NFgpaUAGy40AwCsnLHo36TLvt/M4aUdFgrLfbh
2gs/4ETMOGlRfcyTVUEXreydXixG9Xeis2chz6TFzdYQFxjK29Edc2YRDC/XFkn4
S5ZriHhJBs5bkxenLEtPLxAP58uB1I8hKRcB8LhdJul764lYi3BEiQDbvtO/Gd0+
8qJjQPKGOlBHrFBrGNlqkp+HRFJ3dMXqCf/Y/v2PXYjbcyNhTzLEAajt0r6+OCBi
WfFpvaqA+0FRDALeoyaLA4pKXvaV943mvAVd8aiylZlCyWA0tm/SzUc0m7KwS0IE
/vgqHMWT8e4qO8JJMvlW+QuAwPJW3oeFFh0eUS6DDBDdWgrSvk4Oje5mrej4cDic
7hXixEXTK4bRYebVbpWkzisNglmqjdJVUfplzJJq46vh3w+DBEXiIqGvzCS0oNFV
TeQYG4WvYlYjjkainszLvaGWvYujjtcCA15UEoAMcz4SWyo3o1UZlkVLEcbU3drH
i4ZzMlLxyixAEvg3z55iZEqtckLGkXuuyP4ZVaktvYTKCOHVYBUNeBVS5TFTUJs9
u7Wx4lYPc4rMT+fcqdiLK/GPR7E0TQNDqwtqquZvAQF53m7+xfL12rrSqI40cH7M
Zig52b3K6o1jVdJPmDorQZ6nK0uvJPjLxFferPi8uBtbCFxkNcteeBJSb4/NE5Zd
GmOUo8gyFOcU7cU968+NYCH8Wn50sPMcjkgKPtVWMmuEx7AK9pXjBo2/ehSTnW6h
6FqO9RL16iZCcaJOBQUMB3lBM/HiRQCNGC2hWDi8KpaF7mFR7/K2kSXIasYEC7ni
AFX2g3TJrN6P8hj013MZd2CruNnHAUxukkPwrvg+aNEWcs/k+vYA5FtSChhFjGGe
4CGJNL5tCvakVeF86WOANyH8plX2YhDXnIhvaX4u/1q4J0QXiYVTEOHV1YLs4XYW
3tfdW+V+0xscWy7sNVkij+o+t0AJD4/GRKGSnz2A/TIHZRW0AD2GnDj5UN/XNPnL
mEDqnpGBgLS2UgUOWYKEs0PMX1QGr5B0hb9SjhNxNBzpmpif6qCsorr+PBSQ4aBE
TbMQoIUEboHLPgp1iOnzrEgd6EQ9dgeKdxUyGsqALD2Cu+Hd8DsgurljqjBFVzY+
VVzQeFi/++n4II0Mn6kUDomTNieWOCJO0jNYfZ5aLAK6tNt1KdII1bnV6c7Vb1Rn
9FkZuSrIPkD/E2VhM5Mhku8he3M5mFZY0nYTiB831zIbthdJ2CbGFL859LPN8gmv
sAMTW70jm2ugVQEUi5jIqB/ZIMPgdW/e2F41dVCTT2RnPsrOf6JYJLHZLY1FJio+
JLmVvPb5R/WqiN2E6u1VBelE2AKEQ9zKP6JQ/2H/8won9bWi8rsdKl7V7kRj1S8M
SubQqi3dAkj5ARxc0u+QhmTtkrItGtXrc0WNsS60nr662R8ZOCkYOLbJU00R1VkW
owoCVKDgaxN5oQrfmf7OFFR72C95OfV9n1ZHXR2WC9UIXk9BvMZInX34V5lZCToM
t8jzBtN/wSqSkM8xdoMJj61GPozRCd8WRGWVB8W8O1EOTgwKW9vy7DN9CNPtIKmz
17xsPXPuvUACNLIXDXJfFjhy/zM5zlbjMoqYGhcYImU+qBsLmuOZ4tuCV2lvHtC5
KLGwXcvGXmlhyCWnDDGLwuTJ/SBJIavm5nQxWFHmM3FkKarZXKGcqWkFGXiBwWRL
hnl8OLgCCkY/TzvjES22V8T5LDrM4tVSV1ezL1S3zRSknFWTXUjYc5cAMDWyHm3M
0iv4PGVC1kIcy6/YcO6guYz+pODuTEhtW/T35gRDEz9FmxM12Vo24klFMz2r6pNC
2am3K5WTxzug5DDGBimHQHJFEbH8Mw1n9Us+iWhtnlDRxYZnJ2lct6VQ6um7lf/k
PCLa5qRnWvmXUaBsb6KZ/mZVgjn97gY0GJnTFNIud4jL2voDA6PkxDBehkI7HHqM
7//Bz6Okfp1m1rPRsX+rzgOPLIjHbxHmKV9tarjfyDYupc3NGQBbRgtp9Xm9+1k5
k0HeIA1v8+HXGZTNkitNitPR4KrzUTXTFgcBns5IAXE3C92/HrR3CLQELamfd8lB
ij1ifLWYKCrWTSBfF1hQNPjj3EBi3J9RWdAGNkK/gRAAIJY8oTDMQA0Q1VFv9+Cl
lOYHx6j73SVkLr92c2nboRrnRuXonrYxCQrvKiDtwPXrfLOACMxou0X/pbFrbBK/
Pi7y4ESodQE78awuA0KXVPoS26jK7zhq60iLghvUPxlU6andBWJEqpzL860QkqvZ
Xgz0yz5NBqHHx94viBhFQDWDc2SgoADzXKZKsmVMFfiNumJUIjG2LEkKrKMrh7Dr
4lvSzV6WOML1D0Q16PNusYgZTj5kCHDHiNYVUtznn5/843YHjX7UhTbBWnyiazVk
ytDVHCXQsms5POn0b+JLWP2SsQj7aSHZmROuhJYQSTuDLkaSNR1L1/XjsvgtXXK3
C8HDM/jNv26PfUo9aFDmfNd2CtqgXkQr4ux4912UFsPp0+kmoARgocGf2RCLvCCw
EqMmHe+s/Fff6CZKotnLu7j9kcsI57QFHKTiHk70iEJtKOq6liI3TwUpc+BWgyjw
uiTnYTka1I14w9TkeA/2N7NbgmdUMdJUdBuLLmHRy/umFhayGDViqTQ2ZtWryNZu
7MaQwXgVKN9BC3twr/2BZU27uOlHJ2Er3X253OAMjyoqWVF6hMiZgvoqnnjaAZU9
WffHsLBhFGkz2S/wx6E1ExN+vYw0E5g/xXv4di3JA3odqaz8qiOd5mEKoSW0Eot+
RvfdD95tUa+fiymizU1kfXttE6GDWWiD49JTlPwIt/h7cuqPgd4zpCLF6HxQ2Obf
hnslgCUn1cRYvHOKWekDXrqw/qvlBD5uxibGda9xc8P1KMunSr5mEgBc2Q/mkOHM
ijOuXKKolEMndSwhEsF7+KMI+QE1ViczkaSBSTSpSiYCb5MTH7M5yM/LS6SQZLhW
Lz9P4QwnD2PWTvWpzJDb6mdfzPusd22SQ75y5lo/WztDY2u8kg6y2xD9NGam5SSR
Vz4xICJesIfIaxBIk6ohmJB59Q8lpqFww80Nvt/be3zJ2BBv86GKR+nu9hIidl9M
0DoO2znrH6NTP10zG7bx2Mxm6N+CLRrsr6XPYUvxhdSeOtog6lGZs+Cxjg2DugMi
Gtl1QI6nKd9lTfl4p0EG2rxpGhD4627r0A3VamzgMOEyoMJ3FcKSoE+uEOWJR5jl
krFTR7De4HTss/p8lvAJaOSqICcvUrYAfvA/FAURrXTwUHRXPYJszrAtGCNlrj35
8kc8L05sB1viaGdjzTjWQ/VSkWl2bjxMowM9LoWK7FGMs4hJxcdhNq3xfUxaWiNv
UokDL95TTpLoEmEgqxnkHhhcI8QsKg3IbJussCMJUu7jfYhzH/BVhEnYfmJWcYRa
xDLhBz+YbFLxGvt+/VH77eNPjJ0+rTsFLEf2upusuC+IHbi2CPFwtLBZAKIuptnr
pK0rwZcEOVtyLHRV4J5FWGtSFtdk1Ds+Z/ieQF0XDbRvn7tWArvUHIJQUeIqzoFj
oT9C1qN02Zzy/Q8uNa0tG3Ud7GEA81DTn6UVW8OndVOxuX3syjhmzEDJTG3xvqoK
AI2PenUBpWQ3nrh9Ld4/tAX43pJ2utw2h+S+dhR3meUWyfCl6MnG9B0bPUJS4zRQ
WP8ugwDf5tmMz5WJVwowx/O6Nq7osbpI8Frnx8nUEVBJN7/1Pq9TFBEFrvuap9lx
WWpqtixGZ6uYTmfNhxh/k9pnQQpiiWrZOaRhm+xuJkm1NPhjqkUB2CS/PHcHiq5c
HykBKylZ2Cy+D5OdL/t8VSA9c0H0SskLFTRmqSOUnzDc1+MCRBXNU4SWuvsZZf+X
hQc7MRz+w/f52DqpCPGUAbVj+gFPmumzLmNImXdOZz851t06fqx0N+dtMVUAlTXR
CL00b9CavyK8agueInjxgmsa56Xd7MwfqqtBoGpl7N6KFwEtkpHxpsYJDlVSuQXb
naH60iEqGizh72H8APZVvKoeOrIcFfSN1m4VtoH2iappqr+bR4SFPYsX12fWD+v8
N4kt2Lag008efOBI5ufngtA4dQy5C/4dEMxxq7hxJjJ4y2s6JkAnx0A2MQCcP7Oc
md8TkNXsxX4YGSptIL52fknf0RacLqmzYqbcDbF0vBo1R+cmtjD/PXiaenLvEnzO
pUtw5npiLA0k7nnR8BNyA0hx+eaXnUCb+pJl4kGNo2WTjkM4gnd+kElQRDCUff0c
HD6T6KrVCI49Kq6y804fDNTPptMNLNBUw5j5HD7mF2yD7J21hxCkCbCQSQi0q8Qr
Z1wl9EEQSJxaUmcySUp6QxE8jViHoo5u0lilnsRpBjQmv05UqPkPJ0R9W95+5AHf
64bf1j6t3nUghgVNeFwyIC7vNceTgcrRHKZZTRiYc8mg2fmsJdL4Xsz9aouSS9oz
YdW6qJ6++7Mj/CEmqbG7NSIkLztLtXHi7gz9wYDo32tomk4UP1vpCqrCfB0nXoPq
4hydH9wLpaGK0mpYHTjdJKdzfE2Xj2rCt0l8TtcXJ5UMzNSs8vM0VLbHz2MJJ0uy
6oub5gaYo0zaACVmKQSi6snvbpT9glYFYikbeNb+aMVGm6QAQYMENHyNKZsVyRs0
2iHdo5fH0Hd9XL2U7+2QJidTRVh5aMiApOcIRCKliM28+xWzX+D8pI5utENvQz8K
Ge9AcBTD9Fe/7XTRj2sy71Wl4K9/t5l0CQF/BGuaUyLZfdNshC4m09rF5UJeYVn5
PpqFHAKnOrc2+Lf5imosOKrq8FTm0zZjh07EcrI9dk/OYL3f7LTVTsil2s7K1K3s
t4Uflkr4ZN2a/Px7thtgFzp85D+n/uuWe1nXRjoIzMi/PFUK5IrpECY7av0Ui1ZL
uePt/yy5jll1yC4YcTm4TeLCKeOIcU2MfJJ+6+2Jb7pRaddJuTd2/HHNva3cbkY2
hDnfo6d5seaH2IpJjtNfIsrUmMKus1CTuHT6gkc7eLaz5v1PN97GEO99OO+ddIlE
M07dh6tSddeaET2oNIkX3voTb8yq/L5yqI/UfpIff+lt4oGD1RlT2QoDUoONirGD
zMYOirIJ5kBgaYGRe+KjRj5iKlrMLBXFbRtfX4Vr0DfhpQKWb9JlEuSHBPMKagqn
tjuZptajfYJxYBzIoymwz0jKyaM1G6qyAPtLN7qUncqhQdPiKAW8XmR+sA2SuPA6
U7cS7UBS3a5eUNeOwVD+7CDGS+hLC7llcnfdY6Uq3Vy7AaXCOg7xe8rUST45icp7
ob+brNnOu3kwMBsKEkqWelH1QDv1pfcxAvhUoyzSpr8PDDDSpfNyUXlq4oWY2yW/
KsJGrA6hTHTDmHC2wrILvj18a0SxcQNW2YGuLBmU0DisMHpYAg6/ouT1oX+6hRya
za8gmkULGHAkC6Pnewa8t9Jvl6BdG0KfSoN2uMspeixW1gBQut2HYBwPPPPD0cy0
K2BA5vkDMzFykrmUcU47qMBh4YJwQlIvyzSkFq0oA8eoYgj1fltcEijzJJMuSTK+
2p+T9x6jWxqUKX/e0/fdY0HIc5wu+asJIPuDv0++/L86BG0pNNUPZvUSbClsOR8c
57y/NmOFzdNqGQDY4jRBEQ+AAlDXqMXjNVC2rNvJEJnlvCtSovT2iSlFHDE6giWA
jgnqg8xCtg+toBTQ9IBnCzcx+A8gk702rRNHiC5TWd10gS2+CRuEqSAuyqh6uZxL
s9MYqmezjuLMYp+0mdtIQEsjwv7CfKhIueFcT5FYspugI7ENWjTO6kWLyy9aEfto
KFwFLBIdxH0C2ftOffY0rIN/Vb9BjkC1V1oHNXs1MZxlCfVR107lDYO29yIlcAEm
+aZxn2ybfETl7RRdvwnZN1MOLXV4JhcuTY/WDhNGJPNMalPKOVJhaX1Z8sC/QpFr
+m/4bu8e18E6YbvQuzV3eO7Xo78M6TEbpZhdAVfKtN5hxz0u5IUd5q+ehh7q5AgG
perxU4Zr2S5iipnAkrNWoNAVVl1LESheSTwnejr3CgQYn5hgSh4s1OetJ+anrJmc
+bZ/ycUJJhNIZUnPqyVQG+RPacFf2huuAqdb4s1bgfbG3sxAtXezKZW/W2GT4Y7c
WK5G4Io4P1SpbdvMe291K4X1p/J8oRjm4CJPDXm0VQpdzbc4SbkRg29gENemx5ex
TWs5ti8NVOcN19YXPYU0bZOsIDYRlJWt7SUCFfTgEIh0ldG1QhjuSk6UEHxcAFcW
PQ4THR3KoOKL2UK3iRJAVQHxaXp2VxvPzEmRaxOBGPZXh3hsvg3h3jOCyKFC02ST
w11zLw2lZdWSrz1KQsHDA14rGXolnsmgq9kuZCy4P+v/Xvrq412jO5Ce4K1Aa+a/
Y0JmvGvrOOvttA/4kQl5IJk2vaeZq8QVeFHfOF4wW9tZkxueNoQzP7JoXKtfXVun
LKUgZDB9LRSELPeeLQB9Yk8Z4G5fTM0F8rWMROaHozzMh77uky+n4dyfsRAiAyGn
LTfprmJwhPDUjzyoXNFsiemBk8TozJqL8AX4tyNf7J2oKB3xypTHdFwih8mzca7j
HqZJgmgaMjoKrZgzqd/73FSG1Bx4ZbmBozKgGwoS8P3JLC9P+gy0tsfVidIK+32i
xHy9GPn0KMfOOx/vlzs5KtXWRcfbj/kuBXrd92GvzF8CqnyuNKuJpt9APQ0Dgc7/
U/D3htwwRYonm99LiuFHtGIldVdMC2213nDBhIaSZt4twQG31XDkytg3F0G64MJl
CI1wmz8sjOYRKRyB1sV1Jk74q3ESyqSOaDxS+8AcaE01PENy+KHZYfgUpez0kNy2
yacH0ps5YMtNUJ9NRZB2nv6AwxtJX2G4fYY6ElXBhBozZHFrjc1GEU3xHgmyzkKY
eQoockT6fgh4po7AGOSXbo9vXG3UjpBF0zvE/r0jGU7RWdTVcZSxSkugAGWXjZ/q
fYmBmhnHX8GKBtlVz6IEcRVIHUg9yR+M4vTqxgYnflADX0pV16s2VB/z1Q1NpBhX
+jrOuVMRwlHkeyKhuuTmiH9dmTHFHBQt69R8kTLWed8H3t/Jje5QhyV74dtD8ina
7oxWyP76fFxbE4CxI3YmE0zK3sNLijNNMKrOrnrFLjvIv7qsvhZDlx9Yk1EKKh1p
5Zci6il4e3hBazk7o3t6zXndrBhGPov8H3XOGho48J//CQsCT4J/elpkNdFcjSvx
EzijwgKsnm6/yIVUBt6mWgkw35kR2k2QuLh9aojPG0yAAeP3s9V2dIu2yCY4p5p+
JeykA7gNdnga9TMKs6AsMObACrxdgqN7dV5O0HZJMWu13wkS7UPupvlYVTGSh0Bd
jNbcNGa9u9lWhDOYyLbbYOUChIDj2umxOczuThVnXCWdwW5hO5eVPxBFcN1/5rPC
iwL740t5suvYb0l9gBFvHAePNYBoXF5fcUfUq86l+nGW+MxRTpl/alRKGr6aoKUz
w6J53DA0G9W7YUmxc3nFpE0D3TopbWxj38SO4iTwgOSpThsV+vA43j+Wk+V2JUEY
lULkOQhCX1nFSMaoprt++gIQQpnzG6+ps/1tAs+ZXyg+ETGoRnRmfNjWn+kXhMfS
jujfxlh24eDjiZ7OvGB0yjMGB+mOoKdJjD1Hv57R68K9gmcA/XxER8Ww8CRWOImH
gSYxNEqinmAujE6uvdGp3jxFhEJIgz4oSnGqP9JLFMrobvHzTdFcM3EOLU4Jqt8e
BgafZvcCF8xWQVbBuxnSF08lz6tncu+gkk+uH4RpUrw5VtlCtMCHXxJtXPyLWToH
G2ET2Di8gtFdhoufWNpoZ8FPHMllwU6SW0BH27fA2TLw+xr1h2s37SH2H4SXLW6d
frMUzvWNGB0355GmA1iVIcF6Kklx6Jf3CNlURwQL5juSlFhP6uKBZXRb2vqmHtVZ
iTg33CjZVw979j5m3jFuWLrVLNlFZX28/zMa7i1zFNCune0N5Zq1WPg1ApuDZkET
9tsySMdEw6S4RS11HJqp+IeUmaFJEs6X2cXFvplDB6km9AHiXVoRDjYfYBWYOJVP
yTyRqGkpjtrwgSFBrFDeuh+rup020wrYscwLrAt7fc99UFDcAWKObBkJjA0OvFWz
c+AaeY35tmrS1YpLCyRL+MZa3OsIbj7Wqpw7H/9PKHVbnwVmd1fFV/OIZfal7LQ4
uOA/6gnYO+2zvTKgS0Nzh94YhMg4QSLSdp0ltD3gLxjic/UkK2BFss6lPgGlMuZ3
ZNgxPTlT3aHdPElHCaKTXc3LN16GLI6IWNnpXAPFvbGi6XMtu2uA6mBMb/S0lSr7
bE/WCPPvBZwLnbnIFgWNooTm5IkXixZ3JKwV9XmyfyrNitfPsnzc/S0yNk25J0HK
VFpCg87SGkLJ+040B67BUxpgpHIM368aSGcP8innnpk1cIoKn/Z9615MiZIgT4eF
SaiEUPfist7YRFP/NgRX8ZLLz6s4MuKN/pM5VWQ6IuqZMKvdeUD0s8rqzpJAAa+g
6zaJBSPWOWkcZCcg5THHyuH+cGNAWWCL7YD2onmvON32vzM+0DS93qjmnuF5F3Ia
byg/bqvMlpWz7Ivsq3goW2V4ztuEAlOROq9Ko+BphACYvaFj0ecd7MJb9OpHVAZE
suw39492vjTn+zj/RB8nr1enw96dJz/sV6T07DPAKvpbGFZwx/S2Uq5c3cWgikvD
NmDlGJyJm+cnddNP5K2kdJRrkpbIvjDtMkoTujozCv3e3F/RiJ5blQK/2rMNSov7
fbLFV6bazX07Wi+uK2wrAyimFHJmn5DlW/q632GKhJVqiHUIujWZcleKrdSSygt4
ygix7JMeNfYYHdn7y2EpbzT1FJKEtjJ9PxI2iN35nn0+R36N7QIDyGlhM3jiOInt
hWVXPNNfZJl9JMHD3n0v/tvIASIRYQOWkJFdG3FFr3ZQif83Gqg115ByBpW1ZhnP
H4TcVLp7I0rlRkG2eIedmpLJklb3ArB8mRTwFabp2AoKh1yuxqYQc7pwSoQJH+cx
88uBAHJ3YDbUjCWjTpLsX3VLOW5MgMpzoblLZ0V1WNYyvXaLkTioQnffldYhQa1N
RXOUB2NQ8AvSc7svMPw0wAsfkiL/hbH3Fk8hByITCbIDiGwAoXO8864Dy8D4wT9v
JkUt1dd1DJnrpaVy4moAGvRtEv5RNvFXCAzcawkM8qYJavRLxj1mA/bgKfQQTDF2
Ow/Ikez7gULaF1mClojL7kzy73NyQryy8W7FKc+/WN4smkgZFJtqdUEsG78pQfGV
+njIWxTaJyyQxzwZdCNJ6kRzu9inssP8U5fU+eXb+ffT8VDdtxxJfWi/552Y9H6p
YGh9prSmtBzKUReVkoVoUBDlDA0ow7pJPcT8QjytSZDtmrLslegcxY2GFFKmukBa
QndrjjdidE4pjIRn5y6/Dr1p+wu8wkRA1sNpjTWPq5RofoBHLvxTL2myNaZLRGZo
mDmCk7/AbCu3kNvKZ+ugS0PwU6VpxmmJEh4NmmBdL3tdaT/u5zGjkA9idvHB8VFs
M/m5xWH+fYSiWth0l+EsNep/nsfZ7w2wwnfinpgIbOEXLLnagEEFHb6lnsiYbdh0
ztoSEMGvKM6jcVIMjV744k4Z2TI9uBbnF+o37eSal4pgvLg5DPXtoMSv7xsfvO1Y
Nx6eQpAUULuE8PZT5K1VQha8jzUmQZYNcaHiLfrYHapt1REwl0PPzBbivaFusGpN
3G1CsJyQ5GxkrdQxJq2ankVcBl4nPTXNbBSFnp5phcwDR+NiHRR5SeY5ohcqeOpR
mFhcuBmnikQjsuPoC/FPFgBrSzKBqZkDjvmYt04iZOh/sMwZi1VoppuYGES+F7MA
eZTPugLRCb762U7B87oG1V5jpB0aRZO0xU0t4o9FPnLaQr64gFgbU05WxjIkv2YO
dgqNdURxxWuyjw+RCC8wetuMvaUE99bn0kzYj/+5WkJ17RmXPnSZ1ZiGvl/2E+yn
5DWT4MRZ5UBlhkEW6PVT5I9nNDuP1NspIIAYRZR3PmXOeS5ucfQf+cExg+nF34YR
yyyTF7d2nkZ7FCk9X7k1Q8gL4gqpAJt43doxdmOp639ErtZCz5HoDsTPt4S66SiG
xiI1oEAdYDv5SJL2BImMh4KJCCIk0oPrDZB9tS2srdflRq02A+TC423vaVtN0H9Q
zODD8lgpRfqULcOUW0wdsdLeebXccLxkY7uqkHIED4huk0iT2z20R0XD1lcv0qUz
0lp61apg5ruKJsILA0EJc9MCe+oIYhpBdGSwIX6/COfjnsIvEjlwzxHNMpqoeDny
pXVu0yBhwTGmjaUSEGlO2xNtTsY3HvtkqPX4VQEv18HM8i7AgDKRZKT8FLYj/0Jr
jHCwiY3k3uLFIXDbGTfVBeYRg8F84BnIceNnb8NtHbyvlKlk2DC+fXm+4hcTNOSD
nc85NyhiYY/FkztMCQJFq+8/En4KeYriHkPY0wJ4w/KLVkXsS23FYja/sFU8MlYy
eyJ7LY1iiWyvk2RYV3OnypR3zJwAHtQIu01P5ggvxFkuIIo63jGBn/NJkFTr+oTP
DBNsoLg3dqBZaU0VW1he6wNsBr7Zgl2I+YOb9vcCaAxkGg4AKy5qz1vSWqO3vIhT
nv9RPYP9i4Hmdui9qrkRZPCROUOmzT5HJWUQCCEt9lzyVlfdc7AQNmfa/5OQNQVj
2H+aFbX0KxbFnh6emCrFH7trBSjJen4FUymmsoLVjMrs+UOA2WIwGy6xMw6jN1x8
TrIixdGVVAly41ZsfIimFv/a6B+TCPMEm73e4orQeSstli1q9JshbJVr38wSIzjh
2YSb3OJWiSo4JT1Jsy173D10vBCznyTy08zzm0l2ht4q/jYFbeabEvuW2nm0M8i0
gRp3H4kjxoSw9qtLVYms3NT0TTIGc4mvFsjQ6dqKmS4kkioPun3rz4vbpAQzYl8p
YxmmxvZy8iD8p9qhdNZaE+uuErEdAF4ykmuSFjEwL3UEpSqbkjT0XYoi03t1oUMZ
EJal0v6dOzKDsNRqh2LtF0upKGFzGat0u3yDyuExYIs9irROzBVlqIvpbL1NVnh8
zp2v8iMxBnzsq4mh5jjRG0X1VISQtH1yL85NSIhXjvjFTWh0xrBty8wfq1nbOQ+b
kQUU1PQ64CuPOJQomkKuQOSOXTjK4g69fx1W8s6YSIEvgOWzTmhbDBRaPozW3sYL
cTVMigEEAxHXtU8d8tECh59kUET9O0FACoZOcavJCAkbv1A/wb8qiYmaS5cm66vZ
XxsOBaZeHWw3iwHYj9EkNHofpwjDb7OcPR59n/iq626FN9g8XAa/KwwKenn/NXya
FCq9nKMr5Ardk8RhVNVuOtVqAtPYEoJL7D4qf00a//FKa04PgkME8kJtT+3dsHhV
4EDdRi4aBFtWs0vBKJXyJX+bEE9fwgh+TQS4L7JcUq1rClQs8BLpD58y5NPfFK2O
0wI0k4Ocn4HbktRvPvmaHUzhke/H19NVm2IuK3P1nPwFb4GtBwRPBjAZkuxc8xGD
bylZnNFLVNQHl6y+UcTbCSwM3h6KRDBHghCT67cKEh9g17eyC65H5R7zUaCyVxe7
7l9LdmBKtMCaQ8+wI1AIZ9hPttkad/JGufrkX3x3EKEWAYMWq7dZ0nMU6EfpHkSP
sxunnvfMLiWFACzMvZ2E+kaSp3Rpc23DkurD/V22eyKZyLoq94AvXBmgCW4MkOcy
djzmai4QXvEAhMhDMRKCDG5XFuQpZj5SFlPwF9W2dWB+EbPpri2FNr9cLF/IETuR
t+ysNcigPeuWn/oMiequU/JdaMSgxnxvI0EtWzoz5KQ2zHBpGXU63d69qZTz75Hd
5B5qWnDNRl9d0H2/23wY811pbIziIi3imuGHONGb3BXHt+zO+qmfA+HqlcCUyCLx
chD5WEpTPWw70Tv9CCHbvadWfwA6T2wHDR56hUzbCEPwk9F/q9RsKkXrAfEY3rku
SGKFRCMdWbThrfcyCrZXwX/PHjW8x/mC+MS0OTdYDTBCQoeW46i9fWqSvif/mNUm
W210/mbWg5d4vO9KFz3E39cdOUzXF9ya99ccnPbb/rTmnpMECGt4VW/7J+p8wGJg
yyHLlvSfQA6MVUX4ns5i9EHouiOCrZ9m1H/Kro9DFQLW+hFAwNTSl9Ri+shyND85
1bcfGhG7EcnCuN9FawCBkPSmgvxfciS/Q3I5nahUqxOxdSEwsXipyMaNQ7i4C+ih
mObtEQ/9wBkVa7fhBsi+eovv/k422OMd6zys4fOHYUBbE0M9kvTydW125bNGl8g5
oNOSxp2RQ/XUidbNrkLD0kT0JPVqMyPnye9gGTLDvRxaA7nG5YBoU11MbJdQPx8/
G1tvWDeFkt/K3y6o+ZC/zOEWzYHneg9HOehNiMGkctPsIYOUTAqM97TKeJrk3gBV
bV2Ph4SGgqJPYegHoHvdpisdFDlNbt0/syM5X/TFQLKAssApnr4N9juVZNq3Xxi3
JQP9odSUYmepSuXoQWr583tr0iyInAtEyhq8yFV/ih5WBHakg8gTH+7Bj0Be2cfK
YROcofWhNeUsX4RBBSkFVRQ7Q/tolTgHBndW+s+rShV+g44rtJrawOdWakZWUVIj
ta5Yh04QhrwCja3FK+mWlCSGcNFK24fDM0YoI1Dkax6IzGdrcRimcVVI4WFCw8oN
Kqi4L0h3z8kcLuVRPojJSu9oyRqcuTl0aEEhuAmHZCn7W8iZ5WCaH93FwLvsE+NN
5Oca78GPvsLGrk1TAlcZe/NNHyeIQf2UJAOhGUdX4ruKQN0+rmFYWuENKztPjOkr
CrgB6dUS92QX5TRvO88tmYj/1a/pLme/qXfawHGBtjiI9+LSHytziAYPrEfGfR3M
loa+fLwRwbCvO66O3EiNemocLsM+CpCkaCKsdshBEGMwn/FMD+fV6AuydhFNOPZ5
Go9pgwZ2K8GAr9yDPDfRtFUwA8+4woJrts+ONvzevJHMWBsWwtlpUN3irMsB9S7d
qm56Ay9z09a4JfvJVoJq+Q1NqyhxP0RPHOU3G2+76XusFrA/x6Vw7LBov5+qt9MS
9HDafC2lDYzYaXRReFJFriDaF+xmRBjW5MgcLDB67v59s+YjFC6huSZ0wrdLiHPC
xo93NjWOHfqwK8bYwDYoUwqRF/WzdXQp9kfdlXNhCaqkGCB5P4ewk00MTfoHUuhj
dpScpyFbd2u0cWNoXJ+0uTMCJ/lX2DmGUhBfebOlQztc2abB+xKD6fS49vSJeu7X
wmADtWovJHK7z+X0bY7/gN57+UwbMkHkgD+8pf1e678r7MGA7DD4PYA1dgBRIhQb
ldOlY15u4hHjrNt8c1uCpVLWb62SDz8bro5D8eVizH1dZF3yMaNPpGn5hYd6nM1K
NC0hecGsNeLas7+MIOtV+FWRzhHxX62g4jltQKISUGSadcigJXAQ4YofM0GxlGzc
2yl2L0ZNCK8TaAyc7/PdG97Stth4lzSIEC+n+cFeE+O53J076ji3HfEAyI/utduQ
CNVAgUmoj178eSThwUMwV5C+Z6ZzDQ0mQBFQB/r8593yOTtsStRSf0sBVlpwkvSm
etIKNWaVWcFgScY655hGHODR4HlEiNInG+vLANJLNG2mwHviEtB6Z7Im009PMtb8
WSKajMS0/6Xx1YgoW/PEPUxmjKRN70b4qF8Xy89ey2cz35g00wakXBYG2YXTwnNm
XkPJr6VxKbMX7t6KxYgwkeMl1uwbYK58NZXmcCs2CwGUAgOBr244fm6JHJgGUoMY
lq56xd8beqvlKlUzkBqoxoHaD0XpI5OZWxcF8VwKXoZgXJpD7LZOxYeQPXX46AzD
DipTGe/9rPQpoLEcQTlTl6td6NsujZHAZIGeeCV6tsOL6jncKWgIqp+1eMnOWxN0
6qB0gckdFdjeZRVUZSJKZbeK+53bNqxwpX6ztVLU5eW1s0QzaMWQC8dSk9oJXVlA
QR3+Hq9v0qsKiZDmwGWhh+6T6G6avgozvvfe5mYz8dxk5tPrCp2JhCRJx990skAf
AcAmPV99nFhxFMq50uppoxsapu4dCba2O+W4+aImqn1pjMlhulRwYDkR/UcqNS9c
P90RqA4P7JtAEFJ3d3ysO1dfdsTKKMhCpDxt6y7JkSRms3IKuTsMTqNTBSbAnXX9
TbGhYe7P6524d2bqw/LPj7fcyopWQOxVAcMtSBA47CnLv3N1gP72+uA8+oSsGSru
VtXfSa4mE5lkN/BcvCzr/phTsJIXUalFgxH4zHktm+ToBYf8QhjzKUCcMC5j1IL+
UUMwIAFUvIuAoSp4cUDyIZQoSrqiAZ/IOMaLjSxJy3OarYVOt8XZRDFy18sS0LcF
atXjMEqLBkspIiog68HvzCRQTSlJSTE3xQyQ9Z9fzsMi6iey4ntR1OixP5oV57N9
VLuSO6lGjOFsUoY5EKCaBuDptiXqd6HR8U6kXoP8QiTN7gWyRTS2EFa6g3CuIP+v
gR3YZ8lr1AqCEkzh8Q/Q6Ive8QxPDVpe6//GeOmdHkciXJLk+EEL4lxjkZEyd+c1
JwG6AZst7QUYZSNAzpQJEDJ2zbNh7dHf7e2SEduoKo75LSP/DY1MNfmmlD3LXgVv
S8gV9erTG7ziWTaOLNOvJcO5vUEmAaOLm2I7YN7mdEByMEqhmXYvII5ucds8EYlW
AwccS3E/5aM0vnw31xIWDrjsy9sgjmt/kgJkx2WSNObzhvsI+0vKKzKUlmBInBLm
h9RdiCe2l70mlmI4+g0P8v6YS7q7OIjgrMMuH5qU1Hudo4R676E3HbAayMsKSJPq
HUYqKPMbyybvYlJZkYUsD8doix/Y+Aj5hRVwb2KJutWxEowjvg/4VVdh4dVA+exQ
AwpMAOpetwXechE7uKAOnXpY8pygd7VwWPnXAkYGYsxrvHlAwjkm9AaDayPfCdde
zp3ahVjqzV+z3J9S5qfrfkDCbdmqU7is3IiAR9wTWQFqYyA/HiTH5UDApICeU4KN
G0nRBmqnBA/X80T8sYKPq5Y9bJkD+u3Ga1Wizilx53JftpvDUTKXeaf+ywxJ7PD1
Z+Bbfgb7HCJBWwyJU3+3CqwqD3b40bKXqTc4vk7jOlXMpPVfyzxykFXnU5qaGshe
2TlBvuzoPvgMtoCG6nrtb47tk5bCqtAz8oyCcqI4ZFsWlGr59XvzxJb39cClcv8w
a71fEZNSiyobCj97J4YZ1OzeN5Ulgyc6n9lYd90sTV59y+A/CALdV63NWj7ZjMLc
2NUVnOtfC9Wqp/pwyEYbHHBuAi0StAOV1iQZ2j1kIAtkZZb0eyhDo7Mat1JYWF5c
fq0ufVJxTitnEPAZwnTla/xT7PkxNjSgMU69/cpPry4bk5G8VI5+g5Vr8MitIsyb
2KZxOHm4CxgsrtUat1dLgmznuR0R83Y4U36DGQJSfeYHvNqqArDEJBa/n1Ltre0y
j95k2wp+jm/e38v/POtir2pk3VzTkCUmaweCeBri3v3inIZ/eXzGvGHjbM5lSus4
sJc+2SuAT0xmCHKHeleq+xnAMLFRy5dmrp1coZmdBBfJ+Jx1306ssGD3DVN4uw5e
dZE+A2BCpfGG3cBQAfCJZoceCpGNaU/qswZC2CFiNPkSbG+tWaWFcVQMRDb4pgTf
0RTA/kaqoacDUummoO7RkQftvSML1dVBtjYicJ9DqysE7AWHXAgYxVuI9LcMefUO
//unXaC3ZhdH8LbezGYXRhkXb2SkhM+jfBfUD2uHO9jUbWnDr+DN6Dx1MTBs7CLO
Yy3BaPxGNZFTwR36WZb9ko4BxMoA6ULJ3Ld6ABinAYIsNkpkq2unRbtMlN4BMTyA
6IXe6wSZP+MoXY2aXh2XesJqIIP57Ljo2K35OfDvxeyTLXGZ8J70/sK+rnKIlF+H
/FOA/nw+fA0l+dyEyylT4oxAq306b3qjkNFEX11zOLK+uhwe2JQlI8GflQ8fw4IY
cSx6xP/Hp9JEkRUaCFZ3bPpbYiXZPEYtiJ927C3RJhJWPf8YGCp5A3hMFtFrljDj
Ee0q7KvSSJJu7g3ctSWBIq7ZQepNVKogcNX+jB6uDhxrlko+2YhC80ZovIX82I5R
rsfIWPhemIbullvRAhyMghxeRpymcGeLESToPWvUTWCm6ZUXVPlXooBqS6PuxoBM
csk4EWdKe+1yi66m0vpHeQwC6D8Qtw1xGzC4kj5xYDj0Xb26bq8jL7lQlQjvNIf1
StVVvLnJzDcxINBeaCxAqSBA55bimKmob8S59/4lZjomiMRmg8AClQR83MvQHoI9
hvqTIC6rl4LA3pZ2cleQWet//+2Noh1LlYOWM/6ugx3lY7ls8iZQu0poH/+usp1v
EP/C7WTctAj1j+CO+GkOF5P+j0mQ8e1PgxF7KCwKQrwiT622sfiTo9xFw3XoQhUv
u2WME3uXX2+0QfqqwCoixI221nU+nirGVPp2hin7HoQ/CpKUl7Vh2woEJhu5EVpT
3/NHH6DB40jfPYohPpiplP9Esxsy/wcbemjxbT9XOY1t9U3m/9urXthYTAIffDNo
98KfQhpQmj/ykEjLbLvLWgA0HtUAWC+Ep+t7iImWGJbLOc/w0d6sQK8SnOi7W7nw
PM9o88Wb7IwSAOnHWP9Qs4pdtGua9nWqLPmLzv1P7yi0dLkxbgrEmhC7pgxMj3gf
kert/XjXJYQiGOV5IyVuwEHVlUbLbAxaF/wv4KGITCkwEsrc54uN70Pr7wNDk7Vi
nUZB5VtUBtW/oklIZBcw5L1yu6UehnE3uWpMdz0etjlmdAGQ6DW7zo+19WypwiA3
U732us+dXfBeJtLhmht6h6t24iyPhizMyXFLqT2uMx4Zx7PPN7Jn/5wWZ2JQYD0r
Wokp6FQUDgM6k7BbxN1fnnovjq+/D9fsd3Ngw84Utcl1v3mceKG1Z29SjItsKw3n
8Z4z59n1svzi3wR9DAA4RiRAg/iNVmslo001yd3WWBZHwi2H1mMPq/IDq+UYmf1u
9FRrztjFBvW8LJ0WkRf70tk6LSh/Z9SZWde3K2apXs0KK8bw/aQy8oO00CRSTwUk
h0A1cypHnk+X7oxDD4dz/X4Px7ZM/mdzkkjETfa5hqy6jk9gd7hXK3x7f1054VKq
djbuTsji6qfLUB3YwitutsM4ILC4LC1ZUQtHMsVy8XKd63tgtidXzfi3EV0bkpKx
yJ5cWVZP0ZrTelL4IniOmokzh7kl5fvYe4fXhBIlVh14lszmVUDhF9KogHzIplHW
FBy8v5UZcD2QGZjUU0HabzUs/iGSGEcrKebkQ7MXjEg3ACyMnpIwrmlUrgH6TplZ
2n/UOEmEgnpwzrGwV1l7Kwzj01/kuCGk4045eQD40vU+iyA2nAKWsXXZz+mU109L
0z7b/sf+QDn7Azmcai+zlPosADK81I2+1DFAemVNu9Ud6WUpBZRYoEs9q/0eg59s
JJaqSbfLXFOZujbdgnUimGYjzY88FsDeJLvhBly27GgPQ0YCvhTjWpO6W4gQFcdV
pRl9zT+QGg7e/dcNO8CgPjZ1u3RR9xqNsoki71fTPEoLyRRKt4Bv5CB2/yNeiMDB
1XpYUWpi1t/7EeplOrfCL95q/mAP+tOgTZo3M6ovNyMwwOFqtoXAEhOWo213SlQU
AgUKxWVeWRy6A/CIMPHkw1xiEFSx0QaE5gdhctSnN4kCq4kumuOT5GYkxnh9nzXG
j/4TD00wCLG51t8IrClatHpJh+FfBeHHSVMV1UDkmWexPOHJjjGxjrBUnMp67gTr
TU7stCjmshRxla3VUkXm728GDZjPDFdiSpeFyBRuibw22y+7mbCcID0hngxu4JPQ
DRN7o0+PGDxSh4T5XxhTWveFPuOa2hi6FFkTHmXdqRtELdNDmxDNPzZ93q8sjzjk
wATB5zasgnz0Z0apijmN2LnlhzG0b1KjtR/gpy5HOiOg/QsGkYdSsWCDQUw7Mudi
gfEesI5DyYvEuBdkNoGNnCRLTkbO4eQfe9FYegO0KkhxMtSltN3197qjfEZOB7BW
BUAS3HixsU32jHNZuQJc5E+UaS9H4/srhfpRVBDgbqNm+YjwSHkKemOi4wuFWJF9
xiVgq+uYQ7sSEcRZ8vYVkuU+7WtASaL9MVLezUJJawfIhKoeMGclPla1uV6rNv3T
3946bLM4BNWx0wVRAUOT41bZ5nta0kdInpcmrrVcnFAVOCyJg0kTsaq63WhXkrZB
BTHGEiquotfF/NAZcQ5vIGeFIncSAlvMt1o75oiyS9iVM09d1zFzZjdPGPv42NrV
pp0XjDATaCh4xt4gEybkWRdga3EEqUN/rYFOkGr8Y5nUbUCRDwyFhouFKuxmDSUd
8uklXGGdNB1XT1M+wOraXYEUPEXBLaZdxXnQsvwKAQqw1YeF1AK1gJIp4Jl+9d7w
wFlHTDQwmtTWaxJyjzq/Mob9K0sCGOLt7e0w8MZg6e0GR+BQKswSSkMCFGHsLaA6
nN0RzQQBtDnHGtDwCoB6UhfKxDVDyHG+zusPdFmHMcHPGcwQIr2pSPNAfN1zjwW/
plxXmqpy18xoJgaDBsY/EbQIBMhl9iXLRuik9keaqTQ5RE/YNkApUCdGWY0tAz83
KHHNU4LD2psOMQzXF7p8yz6IRTzB/Izpc5xJpMBoMLZBn+e95O6wGGjMvFg8Oml/
cs0RXL5dEer+Q/KFijsPdWJ7v/70nYFtt9uQ/t4YYOwkDodnn4SPFJpFb/oQy4gX
u01s6A06Gmz6Ug6y62POqwJqlWqWF5Rc3JIZJ6smo8IIfshcOL+cSZjY7q9H6h/b
ZLxDJXncJT2uh9Jo2ZDsY5TMlE2pqRtrIjaAMWwU9Uw5P0eBrNhg1bPWYxfyzQd0
H6Cvxv35a/TifgS7Wp56z1UPLNslFH6gVIQxjvl21AxGsB0HNF0M72rGjIE8zC8a
kTGFlAPtnn5GJ9z/k2yx65z++CiujMg+ZwKUDehOw+4kVh7wl7kQbI7+jcDbPJKi
E2yNEvxYck8Wu9vdUiXpkjtWBFGMfvbri1eZL2w9sR2Q3jDYcLu/VK0VoqGxMKZt
iC3ltSjsHSMN9pxwMjLv5Cb4/HWmdpo0uQw5aLkrg4lsqInJ2IuwqHNuCmaC7FXr
8Ldj9TsbH/Z1oB43hThyCjr36VdZd5aq4aV/cvraUzwFKtxm8v7GrUb0TfSxRA93
V/AyAl9fpUyzwEZYigPgI4z4lf9eHhPsi4M+3zUW1GBGDpg2M1ilp8HwUkqIVC1h
sDs0jK54otBrXDor2uy3PXHN+LLK0LPar/CnzAvchZlcPuwznyATiU8FhM1CFbpN
E3oXdmRgD33zvhotOtsn9evA9W67XpofLmhWmyLDjyRHvUs4fjudRD6IslHFm8i9
D/0ZP8dZIlCui/ppmNrYaLgKVBJb+Y1xqRdh7zor5gYoEWRQUCRAy+eCZltxdDTY
CtTmoe/fN6v0uZRwxCqmg0f47tYnBOYUZMTllcPZRCyUQX78soslzKhgFigm+ZIN
mWv2ESUSIcoXcN3BCzN2jTa0Y6folg6Clr9czsBRoxpDHtcx9QVmesPtcpr/DDHl
oswy2tWI8x/Lnna43f6sqhT5I8tacHYvw+HQC+CewuBdytkm00XUkCSgMfKqPDXk
lkwNbNrNJ4kbe0zTBPb47WZiphVTdKXC6maJ7LS1uCFNLJP/25o7eVgkkjYoX6DZ
/9uhbdnw79jojBlsCkAEo9gR6NZIEE1hCuSPiJ9pVVLQ9NClNtfIe8SSDg3mU7hY
DwZNCDuOl+aofeJyZdmMskU72xEiDVwIabpvAVawAi5ungj20rZnkhtfLonSahOi
K5H8VlzypwxTDtsvPczLJk33EmidkFDQYPsS/X35wizJiRty12ZVo76393OJkP4f
/dmKrL0n4cmeHJn4FqFCwW0FlUq0+pQ6ijXWSiowqDRqVpp56lkKRRkSSPg2nA9A
15wOQjyLd6ZyvXSRiYLD1f0dhLczzwgQLci/807ZUoyGWdHWFF3tr9bnGLmehHuM
u+lkMYWiFCcJtm1PSPYETzNFj/aUe2IdG9fNX5c6RT8m9gAp+MyC/Sa/pXcFmbZH
rRZYOXAfyyl+QSi3EgNlO7lKCISDg4j2sEXzHni/cLSHksBUTADxH1GhSx3ilF05
5rRcKw8930PEHAvWv+OsJfxRDeodM4W+g6u3D0PLUcPPhkVrjFzhmbLqvzPRjdE5
CXKJabmss+CQ5TAJmKsnnsMYSTK3teq+0kQ4xezAf/MMTzlGqhxe+/rp7lLgeL2b
K2izCZJWe22jEyXLOAAlsP6uZzoGlrV02wB3PCabULEogjpW4zacJK4P9ntah2p/
N2tIBPxZIFITTLNy0hzT/AqotH42heXLZwV4TWTpNXLAlffTqfkYISyrPYuacLo8
74S/sG/ftKf4JnyhpXZNioHamnXo6EUEHR88AUq3D40RIqIbJyQF2l1lWXO8Dav7
98SJYNmgTSuCQiMqC6Zt6d2lhnmj+fPUIpnGHJ8mDXOiUnKh1FsQZSeOzL8O1sd9
NeV68LugSlfWeJ/oMUncc3uW4l4fW3Os8PvkYkHru7upISTjDluZTe2uiOPmtk4G
xvQP5vAF1rAozbuT+apDKlJagElu2XwENNzwkcH6Fd2T1LMCfdZcxOnum2ReyMQJ
Ab/6YmP9nbVSID+Gp29PuK7/x/zRJOZQOdCn9hJoSUllV79ihHl4uuuL0lsDjmyx
MShi3ibz92sr+O2Pl6BfqwhbRWuCWI+rsqY1qc4sIBRudxIYztDg4CmpZ7K2kDz9
2cvHFytN2HOpx0dobkh6iQTOvKWZqLS5sdi+ujeTwfpRv/hWWlwcG5A5vXBRL6XD
CT2V9ZEtjMkB+3iZCmCUP3dNLCZ8zj+CC5VBzOqhmtMiN3E4c0z4rqsuw8NrhzUl
uXZIyEwfFXdhlcpOb8hZOgmUmcKBBOCHFKJSPxTt+q47e77mPpheo76+ry4kDcry
vjGLMiGf0Rctv2Wh1DlcKIDvjP+NpZHSdp3k5y6C6yZi5exb5zQAxWFibgHGqUZi
L0q+JO20UFDcVabAxJaDXbiTlf+J57s3w4nHkGoEzHGg6wAHbz2fmYY3TjyHFhXB
kGHzl/SkeCTQjTKsmeVhnghrwpOt26XYrxNvdFHPtZNDFOx0n0Q4XUgg5/5liTYu
zjAvkV2EAJk5XGb74YHLtF1XUwQcHLjyHVQyaKuZqgn7i53Vot6Hj+xqGlRefQ2U
/eq4x5XUl/4GiEzI7EW7gDdnEte/n+viK2mRfghPJscq8ECguukREtjdsGWafnUd
2BryZJjwB31u9mhJypsEzuWVJLp8Qq722w7ItSLrJWAsXHK0vSzZkQbpInI1JVnF
reAVZFTzKCS2VSO86o4Ek00LXJzYiB+Ae8qYPg7k8uKwvryThoHNZdejaRhbA8Bn
7d7hVjdxcuvQHxEDB5qqzLFMOoqqkF1Vp1KmPDK0eS6072UMjZOwFdPgROgkY4It
CtS2mjfrHN72+3knh4QRmJbN+a/dcLJ1mGBzm7m6lv/V3O/PCDK+vcIUtfEsYyBq
EigIBVaemRZ2frm5+xb7LX2Fji8c+MlM0e1mSx0MR5nY3p2CfC6GrkB7V0+znAWF
HhpLIMNJ8XUAUN+4vwjCaTEwu+r32iDC8OyHOZt2EQfQK3dlKLsx40acY27mSAAK
jV3mFzPrpc7aqyffjEyIS9UPdNLpeIBJ6/K2C+ne/laM6j9LviOJNXgDWQ6bInKC
ODsUQLStnhGKGCHrwrx0QYfOgilnAPLux6uKJEVOMJJxdqKjEa+Dvi1IrVTiDw1d
91QJPa49zAHpKGi0AUtWvIsanLaIoMwF1RtM18tdZ6VWWXEAJ4XA+t4n9IbSAkNH
lEb9UEvYhz5p8Tla4vOt1MbQaa7eJJB7BrircNVzJRu0S0Czwz5Nx3/XLBHQfuY1
40Lr6Tx01VaKF5xstA0dI3JuhBwmvaf5fmKa2+7vz5/DQnYJ+YcOez3Jsv1Zk0wm
Nz8dFTI2Ov/bitR4SA9SrmnV28l3VRQO/d+5j0PPyWYM0RKCnh7S9ZAMHX5UVD32
bIi41ny3+PrCw/hfCgU8mIv97uAU7Qyw1Gtn33CvmhWm7ssE827SOdgn9jHxFvDi
6PGihMnptkA6KtB7Vz4/OGAXO05ZksnlW2MXjObLRWFLv49RIOTss0yRfo182Ywg
Hbupwpd61N8dqsAOgNwTIMTCSeJkrQKvXBbCVCVrRn+DSfBF+Ya3r3f57FDpJZvT
Om7nZt9rvHDjKly53MX0x+KZXobzJQasp3gvUkFwL8Assch7eGBaInE2aMaeEl90
NoSNurQmyHt3YO+4xtP/ZMSao03lAoKO15QVwETPgpiudgDhAzswqCTRBpZYjSEm
OBAgcOohumiZyEQErMvBjhQAUEzu1cGWE94xYK3mjlB+46axYhBdwlUPtZ4Dsf03
bu3FJAN3ZvFeIXf/yN9uVuMM4MSai57v/LDy2VRpJDdG54T3z/8TNrIA1seS0KRJ
kJkKLpyId9KtnsF0zmTcP8iLz5nmKw1Y1OcWRvbBSs4wZtZlZj/aYzXMxB6pHOxT
E6EqUMGNcOPq1QVkUMFKbUDcysJtYS+mTU+NZ7TdqZFD7iOycZ8/PYD+wgv7Tj7W
CcWFhBZLIP0By985QoYKAylLAfLHNqc7S1swqPKc/BTEF12MmwM0BYfESowFfXto
IohULXAWZsXj6/xWq/4lsR86+qMqk+yfuhJ9lZDkXI4re0sqtbVgVwDjHU0xf1dZ
9+Ob7SiiwIiziR05QPBP038x7IucVjBjtO6PIDfjHc4HKRonxy5Ajyt+tEakvplN
q9bDPwBOJepGByXaDE91J4swIldaLigmBi6DqFKloqyP/QJ/OpZI1Dlii9W29TRA
Dys0+5Norl0fzsmFryRcsX+1yFpCw60jFaIegKb4zz/wUmkS8z0xKaWSMqDQiIWR
LVcF7gdWwakIVT8Xcz1Qzn0ci6gTWK92v1iV5x+BwNduvJVLkYL6WhrKsWzBH8r+
0mx4DTNUdEcS1Bzf9TGcfRPXecwlGaF0E8RhCuxc1Ef2ktx9+QJf5o/XdcUM7APS
ItI2kISAoD/Gnmj2y4nvC3lgArmuAa/E8wFQmwTDP9jcBUvI4/3Mr6mOG62xYnAb
bdQcA3IiIXFj4LFAV+52kCvgUQAKD/Kznt4Ym2fYikWz/rtrmcvnirSVBtn+nWwc
y7MfZNVJbUbq91YG5W7nyLuI5+Hv85bxo/N7iswZ2DrxgrSfwDormtQwIZW5my7X
Gy8PZqXOMUwERv4To0kEPVgraKTOxFArCX4e004nY07J7INi50RgL+cAQJuNi1vP
MNm7sv7UH8+UnFSQnAF6OVzNigWl7kFF/VLm8Y3+YuTlao2YVMD4y+QaTikIQT+p
MUhoLmiAzhj63VLk83Sft8WkcmJctqr7kayWdULwTuYUMizM7avMbvqiVI4zxWCU
QbxJqDlXZD9UaCF5id9ec3gwzdM6kmshtldVa4E3J6fdYNTJ9p0t/AljY9bZCjA1
qO/Nhq3+ItszImOU7PBjojmjYPItxF1D2rkcX9iNF3ddjKSve12p3PXyfKAKAV0j
F7gDLYh6tBTvGA65nEKc35qG3BU6+yNhYDyOOKyhUg0Z43oSo7u2oMtzNnMbKUFa
1LbcPuj/RoKKuFWHvx2lEiyeYzqtzWFMSYSuEPqpfoNz9xwNEeIhx+k45aA26Heg
tYev/aKXNGobSmKxN5QVKttiXA8LDcalnDjTwidblzGTQa6MpE71LTQS8rPXgV7o
jxCUVefbOi2R54moxVhX8DSe8jhgIaCZPr9m9wHJuLK+SAVzjespe/fJtbNmMMSl
14rUMen4l4MBl/XO1/ZQW4xNpOiamWOhOcB7X8tleKG/Jk5O4wyNijgGyvreDCow
s1ch10cQi9BtLRGb8FAtlZeISvU81EwSZYo/DaI07iwsVubzq+I+T9WMtodaqSXW
a6rHXNyLKN0V2w5nsg0nJt+94jZm/HhT7h6W4+mgLvX4UsLaso3XUeVt/4CSB/ia
wT3Ss6DM7B/Hp87UPXwkuSqX5vExLstvQAAJzHOJ3aRaSTmv84sShsDf+g/qK5NO
i7gJu5IBB4LZ9N+OTC1XIXLto/x5dRDgEs8c3A2v2nhLs9+n5Dln9TJC4jujjFqk
f8EeIIqE2pnM8foSN4YS3BqGtlqyZQDmybMY4W8OCw8G1thY/uQiQYDIHzJqt053
6S9AepUMsXxs3nLKYJAseFl6WRaBffRjbmo778cQ2JmCFNePLpqdw9DLUKxOXZAs
9FU4KBW+AuRXOiWlIMaD0Pkt1zTatgkF0tTFTbvEurrzebEtqbScnAbn8TjmFpGn
ni/ECs/lHOSiXm6afxZ70/Vt0kzM1YWUTTHSpNRoEVLY+RKsIJ+QqMySmOMVDMiK
9OmhZw0r8DrOhLxUpGgpNxC+l82UD/7llXIeWvf3kdaIxlTkOvZ97RwLt1t6Pw2H
EpWgIYXXp7pWSYFQ0HNHx4hV8vikg1GtwFPku5TUUxMWjEbGs2xhcpvhI3T8lNOw
fCgdN5f+fsO6dE+di43UIvyzJTe+SEo+DKIX25/4l0R0qJ2bGpK/uJv9Uyft6KWf
p4Se1dxCTH0SFPJdg/CTpAFNkEFxbFE8ypA3rRDY4KrHCISXX10THpM9UOXtEuuW
UG7Xq05Ia895eqMr4VxWqt9+o183IAh0LMimeX7FXZ9S0wM8stMgeptyyDXdjSuD
GhZgHc6s5caNfykE0Lb2HqqVNbL6Fp5g0sltolzbiBQg/OCGmUpnuu5WcLgPu3sb
fajhPa6wq1/JX09GtR+9ghhbnbR7gfH2kLicdXrLjE0gZzwuaVLjxDzwCdvdNIGS
fdH7A2/ZznJGk8w2k49WkBWTqnuizWRYbttZ5n8NAof8HJ4X9GWH+U8g0rRBsSDN
ZQ1/SfAuZppEIE3184oOACN8lRnrP1MjkQIvda24Swzqap3wujYvk/iSUMk8AEfz
d3BAE1Y9oKG0tErDXyz2Yh+iXOpv1+cj3MbQkyY63PqOz1ZlbDODMfY6PT/xI/X2
Mh+vHcTjsc8mKYG8w5Bz/rgXn7JufWvoby5XrxW2aB+hMdyb1Z0ZTYWsr9gkKAcN
Kc/AIX7RurVbrNbf/b/OyVFVIlvxr3dsTh+6paj0XS9vRhoOdzNj3ax8qU74Oo9o
w/EvyAQxjuxW731vBpJD/3fxv+bK1S0DqlWrNu1cRTZBGbdahf/b9KxOfL12fHAG
CP7gq8S8S4/y6JaCchQ/zJ6BLkPJYdl0NHHIqej1cHfMEcVQkZkM1GwwuEc2/DpS
RD81+56dvUqhf6CaqF6IR9cOccpWvikGPxb508D7ilZJBlPgLE1Aal5ag1wPEr0F
y/enJHg/crBqHLn85YbEqdBQ/Nh0sjZCYhOpxvwchKPJlSXy65+E7uGPuYAfF66Z
eKhyt13M/air80Px3wn79T7ydVdOxbqueul/E0oltipmOOVDlqLAFTr5ze5Hleic
79WtzVzONjH/6FF+6ZhVIDchiFe491bw6LKD8Xe9Sw9an4z46eME7Rf+zLJYmhsV
9s/U5EIk7O/ethYJyO4CSsbxMGg1ewFIPHhVeVrwtq6pVYchahrLbAdvQ3e8KM1B
NLHQ1ZmQaqckAZO5+EgvG3D+b2iuT2kewGMJhFaJrFqtsydsF1NsFWtaiLT/REtX
RO4ebrgnI939eCeA7oWPxAjO37/rVhunLJRijh7EAbPDQ0kKckblOdMxf9ItLK7X
OfQYuJRBE/b8+ZJT2v+RHT05wrT3e3enz+6dHPmAzqT7bTajIBtnW8+yGclxQSaP
WIzyQ47GceXunEG/ZiRZCXZsRNUB1mmPDBNHhnwXZ/ufNCfW6QGB95Y73R0REOQc
xRDH3JHEC8s9iXqZGxhaCIMVVLPbQcBIuvlXBUw1lRAo0KLpgywX1bUocX97arAx
sLGKBI5sb9kinjHCkaQnwbRJnaA5CxNUIIZwwi4cOSY8RFW9n77la/2aGZ9x2nV4
nPmYx5+NRZDQDPtIFt1Pug5v2wS3k/3x408a7/OpBMBVyv43e82mSp2EzXMzEQnC
YK+xvP6rRrD9W7bWDtJoRz5bKkIndJUlpO7XmVJpRssECKc3ugitiQ2pGtUx7Qal
7r0sWfb401yaGBkDdhtMNiil/vlrs39EScZYJynToPsbvuJSrBxX5iL9/EaHqE/P
eWqsmLBNpJSDJjaqE91WVJbEje06JaU5/UHiqBKQBxh75EgqBGCWuYOYaLD4w2rH
WRuSykuL+3z33e8K/xNz1PjAwdXHy6/uTtZJgPpFZtaciaRjyxdxNWdEt/31E3j1
Q7A2eDAyCs9p1sf3HKqAjjba02865Xefl0JDwLtaD06krQr5w+sxWmG3+uhFdmcw
mwDBRTRoBaaMZoj9zGX/pm/pyfy+5T8IKiptlXWfYfiMW/9wTErDiIXTTVlqg04t
p9dsCJA314bGwH3hti35yvhQg9KhG6/vn1ngoE1xXa54Cipqe6tj9oDMCBKIPU3m
/Grz8RrL7WBqWSkuRSd5oB1DNSE8z3YnXLU6ZtkCwezYq4STRowYlS98nId+WQpy
rZcEZbWyRtSIN8tdPf2MZLTRa0byu8ng4stj055lSg4sxOr9bMJPO/htq5JvmkJo
h8y3iSLAqknr8m2zsdbFf3SqGGZrLMzKYKHdc9NCJYTHJkW/ogrfDB6wv1kOHMnN
ndv96xgQO8qO7sRTu9NGY1KE53vfDKPdluB/gFNJARIenqgfEZkE8LiBoNyP1ZJm
IMMRK263p51BXKqJSjxsDgkOVOr4Z89v2oqL7peTderJX15CZsOMYX87K+sVCxf/
F1C0LJEUzndWYAH+K5asVIxARTxjAflQtfhyHtSj5VGIj5cYD2WCffSULuKgGyfX
f69oURPWyOpz9W8swvsqPH79ONkAyzDCfw8ktBEhzKkFgZUAiIPT7kw58HL9TJFk
ghBcgK8OJeduIc83SKJx1LcYQdIOiwHW9IKfPXzeoOVz84SNYC93sXKdnU5dvYL1
oPqky9GTOJEmnfql31LGmv23QMZfryIIaTZ+Z0Q3WPPpmQzrfLwQIdINm7a4eF46
cBD6CRJZYyEeFA8ktd72jxHZ3rIOhG/sqdSbC07yN3KOZRgIB3WYcLsZ2tgtqBPT
1YOiVw5X4zqhtbtqq27rnRqHuPaOhBgi6Dj6wvEHaHIP+2NrFOAQ9Hu4MsxgJFce
WFuQa94o/u0CvsR2f/4xga12Wp7Iwdz+7CqL344jDPF4NCIfw28d5SEhKvKKgP3P
eCWzC3pl2miTBAWLHafAQOZproZvlKn83YEqFVXB9S60OzP1UGt26p+QuGr3LWlg
q+93Z27Wg6q5vSrWjtuQCAyyZh10GyAdYxDAKaxxibcBgvJHz+0S2lA2va0Zlp8V
a7vAaRUhMIGaA3ciplgB6vI+BNHGxD0kAq0BaUo8a2BxMeON+PiTfnGjzAD9H8i9
VL1rO6zeo920gx83WZPHmb5b0OdGqXVGtQpBrEdPfRn0Lse6gtpV6TBCn04DjO3o
1xCnSzHeLmKqunnvrh/yHCe04fqWmj8/SXMCd0JTuVcfeEQ269IUWhZ7IwgZk4cl
`pragma protect end_protected
