// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rl3LjaWzWC6xm4ytmCpij2bbBzW9O1BEuxkmDTKeUF1SwC0mF+KYu4j53HZbK5xw
RD3MMUJ6c8YRdWPX0BxHS4Tvc4CW1gcN2gqkbjyPYW+ZQaEp+pZNEM6Q/E+FcOTd
534En/kO9MJEYIztqhB0mR2lrQXx/4c/ZSfP7UE9v7I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1760)
oj7oCos82z0JWQXGASXiIWgbEwsbKfOGV2PhGO5Qa+iFyxyupCbIsc5FRam9n9oO
BGZhvT7IkvzFyCjoFm+SpdahMXevN3W+3zya1H0iqv7Q7QFV/CDRDchtIDqsks1A
uBBtttlLOE9DSzA2SmLpgjfe6vBrtbfdw+A5rdf4szIB+vPykh24HgeMojAcvxOe
tEaHOYC+PyUd4kSiNn1Bs5BowjXvamKj7S67MmKLnbw68EWZJOaIMdE9dIT3i1aO
MOh6jyHzpmYmT9jsUuN9sxqlUHjr3ZJCQ2S2uN3kV9qwZRU/WcvI70AqeqCkiTei
RWnEqMa9a+VzM12gsJKH7NnxB0Us+aJP9SR+3FjVckxBRjMGAcLDOuuOw7jxo4wr
ySLUhPvP9QMKesG+5oL+JDPwR0RyZXsswaxG0aBY9j2N7xpzJe+KKgR9qzSwShDW
ejmnAGfKod6EDYc5beX67u2WmHgAnwSM7LOVj6zvs5PSNL2Z0bDDwkFSrXh0Wakp
3z/j5buDZUoPLb5R6riDUb1mMcVsVI5x6+uVXhMuyWmMpyXTGQCBIBzv9IPm22bJ
3f11SzNRTKrkupajQ9fGbyCXpkTuXkpyeoBAvVt96omlezpYCZAx6n+Nm+ILs6hZ
InO46C7wRx+6ZGrjHqS7i4xzygUUlMaUDjMDGIohkPZdrRhsGUD3fZgrhLxBHIIR
vXtGcV+n54hf5HyVZ9pyBZyzEn0W0hDE2kpBxrFslH4d/mHRKJReW00ZL5bGQSKO
IaZFbWxqw/oCC4+A6xbVU83tlbkJnsFO96jvqT+H2ajt5R2uSuLMAnRVzASrayRr
sdbjZKwmR9FcxkU5g31c9zng7rFM4n51SzwTTjEOaO4/1pd4oKY77iyRxQSjSbr2
cq2RqjR2DAZmtdu7CBLBY26X7SFWJaEzsXllmuBiZV91tPPwAvmULeeTRLh/KhAy
+K7RzM20SEzHtGTji0/6nwcb3YZMg5ZiRcA/epGB7EoTrTjY6jPoewpy7Q1pb8kT
pp4T1E/clU9tnxrjKw7wn+dkq6fM3ZiM5Xk7a2uvNZMvVZGwv0Wrtn0DXISrXzL7
NPglro+HB5fDUPcpcPZJdzj82NCVMAtzS4ry8b9zALxrD4VQWq0n5y/Cr747yspj
7FtIgGNUYT0kAE+VjdMDAkYVNT85Fmgv5VFo77nr0NgGF7SWqHtp5ENDzheLclYz
46NMlm2YXgTqkVMT9IPIhFvWv6lIhlt7AG6wZTVQHc9oTtpV1jHSa02o8EklVBZn
ctLzQeVpENSgpMJ8mcV5j7u6DTUYsdn221gviAxKTx7UHdxsernqw9oC90j3Th2Z
2iUv40hwnhgEazleNjSTvEHvxhxq/Ay4ygD4crJ+MZgiG2cxJwOb6e5gyWx4LHq7
37if7r5PHd741q8/SDNrIFBuB1n11lp4EQcl8vSQmE5DSg8AofBJnIGlaZD9OEw3
XWOMBZpcvcnJ5KXuWsOmx15IDPfKG9w3bFkNt1wVslpjWVbbLojsK7iWhuPIJyo0
XAdDP/j2EoE2CSHsJS1KMkwYkoWwn2Qmw0vAPRgIMG2QrW8A/IM5v9dLmzDy17BF
dfCsYhZWYjtbes438wXqcDZFo0OJPOVEB0UIeBfj/MgicdfHdgI/XbLhtS6iltrE
GP9vWqPDZBOLQqoraEpqhpUBv/2rx3/AAl2T6PVxlqUgwshu1A4xiKLZrZhYOMZL
vgG92u03PyHzb2oZEB8lNHEDEFW0IY5Go/xS512vdBAeMHvQOMHbIul+l4Lt4ksA
2zMUk+beTtcjP1GLwe846rG7VZknnFFPRoaZ80xYTztHuWRGDuJytKI5tgEGR4P/
Ur7MYl29uWardc8uZo42ztYRAqgwDRgeBaUkd44O5m94M5FQ/si/qunw8rdMvcfw
GBo213+esH8sBhylRbuJOTizng7KB+6ToWX+1vnm/Cf+Ew3WBUHOtygLBhjWZGwE
pgSoT7QePCNmdMAuhlJ2gaS7kJT+0TeIZs2F1ZsBdzBjmDmir4ObrOoT2Oo4v9hm
lqRM8N2kOIckAZ8huCDynt45xUwExcpZYziNoSL2MHAexoT8OwRylLOUo50F5D4A
3bFUv6gSBJ4eBOHFTsifkFt4tm5RsrQ7e1/BkOYC0y6xHF2o1Gd+gPvGNsrbrN2W
kiQv7EsrDJZwylbct1QoXdZl7D1MuNjA2or2BwKz69PqtqJ/V+cqrDffo5lpLsRw
OP2nOkg1jytVI7ivaMhvjQ2SsOGdpiPTDMA2cude4AS2cknThEbx4NNLJgo4vtx+
p73GzoIU2HaCr+deZraerljkZOX1qreoV8tBAqM8QCo=
`pragma protect end_protected
