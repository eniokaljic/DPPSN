// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WBeAk2kceVL3ObdmWfOHrI5IYQvZ4rTqFuvkuciwyAcNWb9pHEznEq5erL27UPir
FWHFcbWcSx5WItxjaaI5mDv/QyKz10PmME1yD0SyFIajRJMgC//+k/f+ijFX1LYU
oYQpf0z22Z+uMrBXKZ3ozVypnNzWf5O/277eNBtf/mI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23744)
u5g066bXjCfhrtdIKiv3Xazi7FAP2PjI6gxIs6xN9lOXSjCwEYOUhTBFTFGI35q/
FBhXzeIxWLSHNj8GNLmFfFyRP87FgKpvCfyGfciO4Nr+HwoQa7i9xiZGoGKYyi5d
JBwNghYEvZfWwwWX7IbalhxyaQ7EO5AdmgrRZCE7tRxKvC0EpeCpTqaOxYOQ7ODe
x+wuwMlR7tRx/DPmcCP4/xjIZ8y23Bd4W2kftL09ejZJGVGjeaAgiiywOAo1a1q9
DCe1iYtcNHe0i888DzHTg3MRnqnfDF9yDUhSQRM2v/gsZHrTLwBTgK7GF1aXghZN
g6orEydvhd/ZCtDvZT9nYN0xKJsZLFu69/KAaadZQNN+BzLUOeqV2lXmV89icinZ
XCQ3XtX+/TQBi3drFDBksemGFwgfHYEe1v6Mi+liDrebNljJYxLkC5l26epAPa7g
gqOTI66hZrcbSx5+3wTuszVnAVb0QFBnVyLe6tclcg5EA7ksj456d9PRaZSqTk9N
Vv7lzAFrNNAVxU9bZoxZQRN9uJRdK/q42PzM8/jDfFsCFKmVBR2zNTrPi9U4C3S7
PEns/ZuitoAbnpNO0ng8d6GRJKwJbzawOnteqXy/wsTktUar20a/GJQn49LFS1X3
TvZjylIMwYx7YuuXSno6gtaqt2JTcWfbPZ10XROfz2cHIAxKfXFi5kgLcdOQwXVs
2JJC90BeV2DfyVJVPC5C9CJPsxQWhw4tkOvfmxi09ijkMFvkWR/xLHyLNFTvNsmf
II1L6z01icrbInAkGFGuLqcNHcNhw15hATqvlsJaeI7Uzu++WbIzv6cD7sAfZBIo
AU0+0iN3sfhyzYBKv8LORFNmNYQBX24wnt5tyDFQA00pbSgxub/6P2N97YRLRHXr
4ru0+zsnYsatPHsV9mHwlytzwml4Og0joLNKOWxvzFPHOYRvdeqU2H1ywOoj/XTg
54cc2TBJTVdspCACnJOOG9renWMZ2i++SYPNJUKSa1bA3g7lD5pOadhYB1OOGjON
uEFV2E6CVDPChlZyGZGeaSzV8Pelu68zGpm1GFoXxlNdkvXQGNQstTim9ytKT8He
3in58eUkb5mfYtXou3oZB94YNGww/INIf1nsfyRJIe+oCZVs44f7WX+XIpOJrjb4
QZdsNJG4peCykulbG3lgCf8mlJCqKYe0+ikQLNPffqx8KV1IvO8FtvohThqi+D5T
QVam97NORXtJWxdzBSUatXIoEco5F1tw5hwN7jE22nEQJrKEY3eDinNNPlgi/F4W
Q/hdQzEaqM4cb23EPDBI2lw/jrv4jMCCsOcGCbf283Gjnu8Yk4+tmp7Y//QpHaql
rwC1w6VTWbPRbmUdfUUTQnHBp99waPG+oxMszchu5nC2tL6oO6uND045MHeEor2r
e+2FQb4leTjGs6cxacRKoEABDciQ9nexgfGnHfTQNVzh6Dj8h2EaXmJHDeDfYNI9
7nxWlDVdKdEb2aWr2G72dRJ4dtIXd9WdI67n3Va+sUPz1Pt8rWDyIJ6PkdW9V0+t
4DVA8F2bu46UAeSos/4HQCYKmv+/OFeWWG9fhqT92xVxpGT8kcjMHwY30o9Emh4s
LID31zqU/iltrg6cKn3cvqW3II2WyzWzrfy41vwyl9DI0UL13StKTukp9+qmSNRx
EN254bD7Y5j79r+5PUt2zlheZw1gapZIeLxipB/j7hlHqLgpkwH/3yi6YePBWZY+
G0INJC0ULvewe0hQNQwD2Z00i47IczakFG/f5lykNOEsoPWVvYHhIkPQN0D3biFY
XB7t+SjrOxoPSLpcj4kGX5WL82H8WhvxDIyAVW1+9MUvIujGRh36lWTL4bkk5mbJ
UeAyvh4Np51hMRUk60X7+g/jUOBCMoejnv26YaS1N6ZNBiDd37zvNllhrZYqhTTb
0MeJl6Az30pvGD8oBjmaWQxxyIYrGrBjLh51Lmjr+AT5RuPaVA/RtKgUcoTDllpa
aOrVF8XEaUVSk2Fx+UYIDQo38qDvQHircf+V7vqltnG4GCClDgFs1224II+tKLlK
qlKYHQXrfVLD5euvQ9QiLZV37pbg2al1Ak9umxeL0IxGoXqOY6bOBOAX9DPnGXd8
ZAmupObVqiStTDn21aNZEm1+umwCdjno/Ej9grTr2unuSuNMWRCqCrQP6KoNXW+q
liXIUpuEmmyFTMxg4IpbhV6pMAjEx8GdrHZCkghZueOq7iQSAIJ3xHkPAcaaKz5i
Qihr1DqSQdnC9laSYXZqSYKOMQiDBRr17e7OAioxsY3O8yfhx5Q7TlXYAvRU1ZjZ
xnCzopNMc+qGpNraiuKN7jJhhCJJmSq4dSLNYTS3EucD0Fhqi1wGZDpq1H5Ycyyp
WAYcIrNN71Huv2gMXZ25v9wgVVCjhZo07QWlvVBuB/2WiMj9hhyHPxNlLa1kzBer
T7qm6AsjIgAjSL9WUEW4YsUcDty4Oz+kdCMABb1Yb0sfNUyJpgbwW7IWWozIoNkV
9sv6v5BW4LS4rd4vLe8r6ZDxB84DOWrkiGUDTnRd4cLgEMr7IJqnhppJvaiLX1/P
oX5LaJYjkgpHhuP3bAaqmIv9Mlnu2/YPG1Cfthk+iLv3CcIjSXubTHg8eR7mEt7u
JafAXhVBILVLGAu34O+T8gU4zbdi+X9+CcKI38BKHzbPK0cMgKeXe3s8sTuUKgtQ
8M/JULrcOu+TXGL+2fvrum8tWdRW3800/L2uselpSUNPMZ/clY8gtT4zA1JsDzu5
Zb+9e8wbLPk0qN0ota6h+6tlfQ+zzb8hXcVr3PnkGMf+/2eh/zPiDC2wAEhQuU/o
cBw6eM7G3oXF8NzMrOTCo5MTVGMSD3N/w0alYnYV6b+U26oAD3cclVqRTjA2nGch
v1JvNJXb59H1ZMqjPgdMdkOun0AtOirXjvADtrimcQr3UyxOfwWpN3mtVCGsvVgI
XwvH0c4BNUpBPB4HggFjtf2TF2eBVKYSDe4ooMNRE7f8BRyMnI8/jBC8UcvPQtXV
mOVq0zgzKXIhpG+CjFYWSciQ+G3pwoc4a5KCG/DrWFFd8t22l6XWHyHUTHOQgHXC
XElcvHc1MyaO7j42/+Jvp+LOE/67bNuKLXROKLsqqnvvniE8/tjNgwcPGxkreTUM
xWYjjmwMs8943gyv6EL/6eZhbTVLrRIK1PZAuts4OcehghV8zCkktr0s0PHzHUZ4
zwPOW4d9bIZCxTsAcd4hRd6Mpczf45hzcD8gGkisF23xsTaArBZ3e8YocYm1OHk9
iq7R3BBbYBjc4/oq1hVuNL0qdCMfwq321XV0Zl+CU32aJeuD026BfiMJEWxpk/Ak
atQBya8mXb6AuOr76UMUL/Crsr8LIwhnlIA82cDHq9UvlM1jwvI+Ij+CsbRBIQdQ
/4vVdPB8bowUQdDn3InFneXMRgq0Uj9QHsT6XWGIpkV0K/CTJ1sT1rlG5Z63VkvK
9fWunKDmjOKY/Ca1cu8a4RgpQEg2BkJbQ7C9IvUw4Qmev+1JL4RbhkMeqANM20Vw
tSUrb3PIZyfKd6VxiJtkaEK96wcriCdFluRZXqQPWMf6e8IinuxM1GOK6nG6mAqI
hHcTNgmeWwTVJene4qUtErMJ5VOsgt76lVyz5w2wPOLKB+f7iRSDnsKqnmx24Eal
jf7JLaPfF862ql9ccBXdHGc4Vrxz+7T4FSnr58EP5vL6uQB1Xi9+2IHagaZXP5X6
EmUfHZmGxpJHmPOumcgBMQd+SY1DPi3dxUPepAR+YpsehCso1ej9X4vfQ3/kCQAi
3Ng/ULe+BdouSLzXnzemxfcx6uMBdwEEaNsmfmnv9rX05Lug5tOPcjJpTUo8qKyc
CMdIL7gAzLWlxO7zslTuvkvvrSk0gmImQdXBgOLtJ5ENDqfvEd48IQWEzhzHU6kF
CGLSvHeSdj+0ZHEGT3Sd1eHwT1lyR2EZWyqXE1e6LDnnSwoeIebytIc5idC+pWA1
M4gsC+Y4UG1cWl/5mSpBRhqyT8dNKDnyAkxijb30N0Hh7km/wvYRp1rtKwAdx/Y2
PdqpSp+kC1rmSC8QtQzHYPAk7909obKMqLvigXL4lBqd4xXUaksWdHaYYMVXvtrz
BbSnCvym8teY3SWE3/CyFLqGX+bo4amDVcLQW30+uiNlwQ1S7l3cDb8Gk0h31exp
FwZhAkFyUail7cLz6TR1dZSwirywa3H73NeQb2UrQmCL4zp21uIhSbZwIdO9o1Ce
hoDGhCi6b/QpC7dANQnwTvtSKdb/iq2pWZVdFVvIQzJlUkWwyTwCO18vXpuXt1hn
rKh4h78DuQ7fjYCLwFDkUs40foGO+TInm9raTDZ6wwTdPL1OpOXM4XYngXZAfDd2
5jQ9s1TdVGJc3nKe2bLpl89fnWiXqKZxssOZON3Zbf86sw+LoHw3Egx2XYsBZkWo
EpcKjbpgD8XSnPD43UnC+j/WEtyxvX76sBNaeSwjn2QWG3hJR3whtUPk1sEa1KUv
HD5pC9CEYpJlvbfnzPD3+eptW5YI8oFYj8QKsWKY6wrmQRml2ubdWYLQPKvNvdpb
z05R8sfcceO5rrVY9U2d04XbV6rtAtDiSaNmnWv9mdSNf4xyaLZMOtY7FMoKRS93
G/+O/Qd5CJzb3MWKFhtivFjIODkFZ8GzaJ1FiMfVNZIyYW9vCiSAMtL2bS6T1ppr
7CogrKK5dpYyrn7qy2y98SRwAhOVEg1MX7UbjBhRrxtLtLijCrgpggiiH3i2limv
Az0Jh31hAfCNYHA7D5JScaozRaj6qe1I3XcjK4Bj8w/RYE9kqHdgpzQ2JpSqzQa4
xOncBkfvQ7cfvktIB6fSlxamesEZCSNPluM9Z1I2CaWAtL3m+rc7KpqDv6kwB6AR
g3HBjuIICvdqMhznC1gzCVc58yHiwp9jRquph1sSaBAKA+Wy3FsDTx0vNZltUCuV
Wnk6q8JTNOAqjwUgtDuluYoO+NpGOhxwjeezAGWNW5jEjENlPLKbykd7pD+9lBu2
81csWYcKXvHncpo6hYnB6CJ8Hw1MF8dyTf/Jg/hi/cJLXkYfYa1MucjD6jgCwwsN
gwWWll3WNLTOAR3O4VYVF8+cwKK5DMUXGBn799zvdLUyk97OdYhn3QPdI0YzHOOE
obLEjqj+zWB5apEaT2mhWL9Ax2MN34Mhpkrfr5F4ixEKCmyiEAqlPEujNO8TxSgE
FAd4FSnNL1yV0KXy8M+cdZhk8Jg60nOwoTsrOxskjSLMzPHAuR+NIAYB5nvl1sgv
l38aDEQ5JCmECa/ohpG+QZBoNUTBiIwJL3evOeOafmLCNwdws0t1GHuIMbQIPt/a
Q48z1ZCIQ8pu7YSyOzEGeXjnFZnWbvp6XbFqX6z3lF73etII/TiOMCeC/1PjFWoZ
wwoRd/lxEs/zToQgpYMqdyfR+FlbApadBkb/xn/TsvPElGMRVPXmLsdujOGIVF7x
yR06akGkuf+lNBO9fuVV7pbuXBBXsRMAfJivOGIFbDtV4s6recleLsNG2BjOYKMu
EXlfiVLPfGuY70PqOvuzUBTLP1dEOCsxiCkwq2ovJS/+xFu5dZfdzAj/PLAegLrq
I/uQSooED4WejuPOpfojL2a1Cw4JVZZk2WoFLqZGjArP9yreRu9qMTjm9gS7XyOu
v3ulMqvwicwmURIi8Uwj+zoFHfzdCg1rsgF/Jcna7qYFU02gPRmovWELxwaC5VSU
or+O7pk1kSyUuoVTVraC1+c9yrXJRZvN/u5D9Kg3ZBZwWaKJc2RPzCqjeLQmbFRj
w0sTiTyV1mKmOOGEGyHmNhRDwHkjMAUbX6OvQX3aenTeaDFfgKYeNiVJya7PCBTN
SmdsYZo9VqkCHinjYsxihOGonCIzADtvN+xrkTRbpm2LdkwH4D6KinCRzBLib5gz
MEsGWMkp3In/l3QqDq1M9h0uH/1+awnnqXwy90G5+jorv7KQ5nqZBR6zEUQJrMZp
Igv44uwa4o73dgOCqynj7MP3aZvJsw7tqRUfiLhGlUK/9JhTZpGjQFbo5p7pz/kL
OKGgPjEydeNftK8LKj+S87FPT+SA2n9uQsscXyuMw4z+dlDWxvAiMyXrd2y3PNEe
VLXWbNeMc6+AME4joEaZ6j5kQsK3tZfVu6moXUCORPAAdpIKJIvVEVWBmvu/MCfM
GXpJAsJuEXExzHWRmHnlJunxx9yb1tt2rTdrW5CeE51d2fUCfxXFdX7Mp7FnQpqp
9gkcENu4zMpuThHEX3TpuvLJ+zmSi2s3bbZVzZQXoKMeiaWgvmdUqK6V9nUJQJQW
UNF+gmh6MjsnG4SPXiRzZpQYSys/kFuGqq9gfmkK1HgmfcSxn/LyrXX/6vri9GYe
tl7g92VpoZ71CFhRqLK5gMrhZ8ux3FDHKymc2e6UBNv8F1DVH0oWAROtvOoFMXYy
osVVBzg3IIWbddkfiSKzLWEFxa75sIvWXfIE5dBqV1mTuLvcYttk6KkIzejBJSsc
G8WNqjEHHFBuG0BgdkjajPBHE5WybrdvSLhWs+2nsQKLMvNzxgUVYiB3LzgFTHD2
ExayvjCQPUES/Ndaf4sr6m3TeB3lECip9URXbJrPSNoVp7OX5cbiCyiYhbD706MU
fROzO1Cze00PAUcEAtwUqo0NcXKL3w0BZdl34Tk2GuUgzW7dnPWfB9V6N6RiKEvy
dh4gqeqk6wyHPPiRZe52Wm/byduB9cyE8clDUzvmn8cyMhz5nnrSd0n7dxCVcepV
38I7m4EUIJjOOIJKc8OjaSBDv7jJUKBUnc/jPSwXw0CtcyZa+aYer0gp9qUcSCob
bff9Vz39WoiLWQ82DRGq1bb6ekqHW5HkGG5nnwheY0e2zLzb0P44vJrQE3z63ozC
vLH54Hb+yKANVpHaV3wRahVay9BlUqT2dhlCNQBr7/taQ5ViPYjOGiYyfCwyRjOZ
6q9NOp0jJksJLEby73kjw1NpyHt6CkPvIFEhfRbFdVgSTleTIHP+tZtlwkJmwC7f
RROXei1Me5ZmU+ioIbH0VHWbJYSFUNIepGWoSCmj6G+8wgTCYpqKQlPuVvblSzXR
6LxbJQ7RKI/UMjwelzQUkCt0Zxn8yvo5d7XCnXu+VEMseEqb2pOzkIzqs+G8fwzm
/EOJIlh1goO3sJWa4epmg+Vb+Sdp/Ix+p8EVbhrbfZz82kAIBwoz8kaSkDNv2CNt
Hlpzci+c4MvVK9rNF56G5z1Soa8VfZ2a2slKbdNG2Ugaa8cHgD63Ln7DYeARPJQo
01ypFuLs2MbFG70+wdbBAnIsNBfUECvwXb+G0+sSeiFrwXAtbg026nCTUE/18jnR
o1VwsrtqO5XiE0bia33AybiJ4Np4G28pfhhEoAN0QQTdP6xegkcgU7Eg8xuU7M4W
9kcgjDSZQmtDXV3JKcUC+FIICfLcD07IdzmZB8AiAXtOHMWxJrUTa2H4YF+nYFZJ
q6iPnrrF9UQkMGIG2ugWXA5kTTBSjMM3OXqU92vCCliCdCdBwYWbffeRGGskH0w8
363fjzA5YCWZNhawvK997Lz5tQ42X5LIhSCuUtxBFs2bZXCT+lNLbgdVT6S/Q+pP
9V5qdkG3T71ru9PTxDdpVVk+YQYnUdRm0h2rmT2q0dRMMme0x2f5Gua8x9pEPLsH
bPukhGO7lYXPzHycxZX564EWXIQuDPYZk6tJ7X1ryFNqZtDGJ2Zzwv1u4eal3uLn
P/Am6RWaldZa/ATbRRRqu/M3Pcti/kFVrbjYUwfWfoMBH2DlAHhl1MYxE1G8CfXM
Ait3vWmFETuoe+smmK3K1vGh6yVo3Y9+I5qISof2ooEzZyRolGUUAPWjqPtKZBDa
lHNmpU5QzB6gMbDaZ8JpJDhhVV8qZfP7RC4ryagvQCnDz9IqvswG+t4yL37tju9Z
lmJkIp1+A5v+m7UOmBJIOlW1Dk0Th8BbHgWYMRFBB8gDoQlz8HU9+1lSDnA0B4AB
W5dpgMMXFXkw3j79+O7GCiNiqnTjnBsEL8LDUf/D9IUgOL2iejrMjusvNhnR9Xv+
7gnPcwD/KjbH2tO3gJkR96b7MMRCgXcve63+HEwdlm6qf3zPp9kxtQ2x+rM2T5Q1
eTPvb5g+YE720/IVDSpc9VRRYOy/pnVP/VQDxVpAw7OMqb2ybzU9AI2gm+SAwluE
lmUETyqlbtoR+2nK0w13PzEyQRBe4dNrMoBGKcfKGslEXtYGjm/RglBG8L+OC8Sz
9jC2Enxru9+7WxhrBzScZPK8oS46j75LXZcELSsDkchBJz8BMcz45nDj1+V4xB3G
rV7p2C0fJJakSCCqpbsKncsV1XxxGO/BFNXQgCuYIFP7QWqv+ug1johyR3w72ePf
9XZC/r0LYkojIxVR/1aIHEfLJPTqkWxVc9HQxmFrzVxVmY4dEWHzL64rY4ImXwQz
ZNoed7kqxjftd9pKjoLhBQahUguJExoICZr5KZn6+FdRT0rUtVP6fKadUI+64UNi
vB3Frg66IiMFWgRgGKrQp1PYpNaS/f3BK6/NNyac7gpMeenuP+gWOOmbPo7FpNSq
+TO7/X533folBH6fsAXnJyIMloAg/YaTcgGVB9va2wH3IfUT6PXlmmolzyxl0NUc
qcQxA4k7BrsIz76/Lt58Wh7EBWeAi4F8AWMt51JyhND9ypevmO1bEs9NaTIUNI/g
N3aB9fqq+rt18Et/w8JszJVy6OfEmgkh30QOFQvwhEGSLOuyeHXI4hrAK13APigM
sR6FlNEo82bGQtwMJy8SS+ntMuO2L+67AK0q9t0y9K8xoS8LxEanK7obbFEzRLob
gnluqAD28ACWsxZ1gX7F5uQ4H/EM+u1bdXLPYRrVnKFsONGKzpUX7V8/L+kQLs9u
t0cQ40p5ZKgB9KulSYA+U5GVHpYE6UaxoTOQbLQTKs9nIiWDk62zMnOS2cvTROfY
q3DzDugGQSM+clq0YwYfD6EW9giHlQzpzKGQ2PRBGBC/0OUczoa26z+qFp02/AYD
P//bSRb+VmcLlIZxHaP6fhaB2IFnTc2sRImYuzilq6yMqo2acMrVvMGH1X1CKeoB
krL18orDPgNVodP99n6sZxN4Zo/PK7WBl5o2bxBTGYuIhfTeIWWlgFIxfNPePfVJ
WDrsYDfrMjXQHsDDuI6VZBwe4AcGWLx0csh1cOXjqN6zbt4Ok8lMmf5PvpKggxVC
ijoIfMq6kr08emnfrXPCd9RnKSA3oxyUg4n/Zu9hZQa0rdlYSV3lV4nG3vASMKtH
g+huHi4R5bnXtrHHpSTw063Qr950gPZa8DIHVJkRwC7KuTYH+nPU8YeZAyNbGV5+
4FbsrSmkeGDD7Gw3VPlDb+cqky6fnPyov7qhodcOQkUQcvE3jWXuFoRQz+joxmL7
kjngDj+myUyw0FEght1YUeIHkfa8hwqyKigPy7LMxDBHj3UxE3sV4wc2xwYOMW/c
XWbwD9VrnQmrEqc0vBSJk3P+qK3zUm1tESMosCVeIPN22lWo+bvFyQbgMjT4Q7F7
DvAGlguPR1Izadr9xzjjJNc0R1YsqzOwsaxN/1AV9QWeALnmY7ns975xXai5j04O
KiAZhjUE/2GkplnzoM4vt5jmXzxKyuZP1FX3Aso77NQx3ifFDh2IYfaz6YzEoAwV
yYLlrl6sf4w02vag4jHR3BAAM/s3fDDcjzheDo6oMsiyiOMOovA7hCfi8q6Un/WZ
Z5WpuG+jVucmx90wVh//qsFJaQjXosgZvfQXmy0rlqlidSicPFruauV6Do3VUMqh
zZ+JbOvgaIq/QJUgQmfGCPgKQrdp/be+2YeW+V1boGzphxxC6mzpts6twtM1SSJp
mKLafzu8AcNfbRIVZocldbKjpm0lv1Ed9ilZTecfG8NziGu3+YCyTCbTJrAhvCUD
o7Y5VRClN7J4jgSwEK1jP7TW7xFwiK0DZXnGVySr19qEUSH/7V1al82jCGYimK8C
PX4xn+kn0ww9ctrx4OE06qCgoESY7m1phNsmdBTDzpt8ZlVXKLz4KMWrSBKnkAkl
vU1wXnW+GKUVQHVigT/mMJ8Ik9/sbyuxaThe7gWgprXLUMxP8IDK4vZcMWtZ2GAI
/IgW0IjmgMjQp3eiKvw1yFjzmTpu1bWih4UR1K6ifX6EPjS2FEnXoS5HHpI8WNy1
QfUClPmO2uHKTC0HXBRMowoCRyPj0ovzxIjrprxScOOXVPJZ3qhnK7ssOMq1nuUt
nWK2ibbXbd4nrXEyDiJ6v2ulWW2LryGMcelzLlchKxNgAnsiirWWH6IA5zPckrUE
yXGQH2JNE6U17OKzJqgW1hypMQJsiuw6vkblfXFAcjo/siw4C0WXwdOAt955etTf
JK2yun+x8VC8HxhGAbFBIA2FXRQM1psDLlMA0NpAPJOAqMR7B2ANr71jMbkUDRgs
zrpkyKR5KaXIiIBczHAg+iUl5g70aeHIIWBgVmyEoo/VmqopNJT5jzRCCjah3Bc+
IgEwhMB8lGvk5ymbD1InNBQUYI7AidlBWY7y9t02Lyuy9SQmfMJRkdgGDXSGP5fl
InZAG2+Q//Ok2VLBFajLNYj3AO/VnRp7PHj7TH7K3DxuQo0umfkcs2qcSgn98+0Z
0dZp3HdkbY5HzKI9IMPkhLgP2onczaP43knD2cc2QuuFLrStac8PitEIwryK2lKz
h3JEEqE7AaD+fMssclkNUEcMFiTQHTibNxCRgf8znSKJJPzoRNrBX3mff+FLHaJk
tFKh/fWxxV0M6xMSIPQ9NFPl8JARdDmcXZPw4zejpj73GLEJTwd9oIRALxdYJy/s
6DvYSWCS4sny7z0AmcQOVrRozLW2PFv879wp+qKENKeOcdpCfHokoRJnG1kHikmo
JGkCBWpGXUIWiPcBOxerReKMEWJczmtkKbYTIPA/kgJnKDnnZ8e7kf+hUKFv0py7
B7hTHBWHAqra7LjhuBG02n6h4owd5XaDdzSzzuhVdvT1mGs3SZT14yA0iC3AEjtA
Acr2Auupy4Q9KfmWRyg+8qCm6eljqFAZBz6RrkLZDMTxWPjfl8llvFbAt3wlEx6S
Pr+kKPM52SaYvGPFjkTREOjO9rYJ5hzUSDzsxx4hRgov41uv3IJ6Uy36sXcfETgo
Yj6TaSdzbQAjt4D2kXsGbI1m8omuy690kiKS8I68OPyvmLhUCzlkqE4ayallwWrq
3jM1HViHiVUEgqzJHz1DPlpt7eIsBjQHVQPMVlLXzuT5xgYQrQv8F3oM0bFlGImy
Qqeim/RX8KE6pcD2Q600caPRw+bNVK25cZ6pxIrUdWqJLS9KxU6KimpYgNV8kLEc
3xXsHiLObPYzx0EvWj6qS6+0bK7Cy7YclhVFeTaSvGu9kVSSwllVcRcWf1naoIe+
kToz9QJrnyXQdWBQct1I27Bsshw9+TD74Hf0O8KCUjVXj+NRiY4pQMVFkz/uEqDK
kpwzy9I6Q53FuaPI85J0PcHaRcGeP2x6vWOBwSPUjbZtO/LSitMnWJ3FpV2S5GYn
ogprRGeDRel0ClEE90NGyyYd6eFRgcQ1AiRL4nWP10XWC4nidRaOApN3GZLd1FCG
PaZre8PBM9mJ9Lf/Ml4RIEZpjFDpVYG9zKdFKT86jUhzWMlzlSbd+oGQmAx5akMZ
Xwo+55QaGFRK2UQWnzCM/Qv4eQX3kb0f2KXXSlSWlWP7lRcXUMouZ2Bhy//IAypE
Ipa9jDKqF82iqn6EJvrddqOXUNnazgu0emPafG9IknzPA/gZSvejtStZUnF79RNh
6tLa63joT1bieXuZOwSw0Ei2i72fw1XPgBluEghJGIiO2SR6O/y6CuSZnVIn9fqI
04yYxvmIYMCclRfqGIaZtFIQhm/gyYCCs2Yp+KlQfT0gim37ssseOnDmioXLLqDQ
9UFB3iJBWdphhVyjdj1zOeJdbb8wVAQgvhOtGycqSWBZFe6NaetY3WwqMfkyyn58
TacGk2Z7Hng6AV4ywy+JhoCQjt8Q4OXFjHZ7BjGN4UM/P3IytexsyQFl8A77ppmC
MW18Hdv9OwJ+r6IWsqEKehULJHdwxyjMxV4Jtkr2CpCuhGvPnK/3eS4TqiBjUTRu
dZ0tBwfGBQfLY0JANYADIDtVlTrlZWE/yHvjfE5sMSWBMcM3HIX3uY833kmzabY1
cTI5qX8W4t7WHpcpMnd9u6tPLidc6V3rlyTq39kGPhEA0t3/nNZlRE+vZYM6M5pW
gelSkc8pKbHLFCLRuaep5JzAUzrLnrcJWo78wJ69FAz21Vy5qWtnBjKNSR9ZVb3b
4EJfJ8lYJQfcaXh4g3jT6vPqBRM6W0zBtfGBDWRaRQiMUwWpBLvNEq8CNZo4nBDn
wrAwVD+V0Xh71de/sSLCfMlEm/gSC/z+drIhic01WddR463ggqiHYn4kmqiVr+EF
/ABkfKy5Du9T4Yde1HAN8vhSPTL3jMWWiWvdk81wOl/lU+Pp6SZMBy7IvWSk2oxB
SqxEYQdT38JP+CEFXuDn+7OoseR+zfpqGiesl+yJYwjDy9+C6k1MfzmWCRubAdwD
O2LUqwNj5DNJs16t3fTb+zKf7KlRb09b9eBo/WhHEsnyZecHri1MkKQ/BHyOUDEL
3Py55zw/zeIl9ILWWE2zD3N0GRHlWC5BFN2dzBAxeLZsnT5KF+wZx2qmP6coNUC+
kOjgkuQ8JUP21MnYDmB8w2Mg6FSgikoGvJsj72Yqes5gKt5opbUByPZYuK3zvgmt
89BYl49uEQvbu8l7oF8HdKM/Z+0MX6PviN5Glmq5Qx69AQglDh2PmxQbZZP8P3C9
jrIG2FmS4qS5NdHEyUzMJMpkos2PArzjF6oPp3iLFgaWa245/h7g96PLlrbioHuV
P5Oqsnc538QUDXyvt+4FWU6OMH+G6vTH2tunx4ZLBuad2lNOCdMaXcboDyhUICD3
pjncZkr0e1RYH2LT0uWpCToHOslnzerYdR7wSWd6vlN1KMxuSw+l4c7Gyhy1B0ai
21bXFuGMPXAPKUz8g1Hag+1ITNDzoYwjo2LPxd39Ld2iThbSgOnc2IUJKkS0f3vk
eDtbZrOiIt0wOJWQPvaZnWhl1xZ8SHqZeZjaDRfMMYfw+hr3JEvqdyNhNSuyG4o0
4WiU9UnHXW1EjSJfb/qJpU6r10pMw97uTH8xJVXgEpkvrft4L3YAjFpsZWln0UV9
8mRWWbwhahrBdDYqvq1WhVky3NhobUKxgj7KP0msA8YBvydewoYkYKLm0aPSIFPl
6NKUSkU9Xft64pkd99gQeD4A9MOrG0X4LYB6i+HKM/uevVJlEjw2TMth5QNfhQNU
DhG0aM+/m7Iy49IMIqpvG2t2WYZAqcUsFyWbgjNZusRtibDVudV3IUfaS59ixqSD
JaNt9+bnD8aguKUFhKhYhxrXN+uHYmcvexVZcnb+SnCehfFwhY1O4TBJ3/IM75kQ
LIcKnh6MQ0uws8RSOJaiJpE5/okCNSKnWHNf1J7CKo21e2HRUfyDrlaZLp/wJtV8
Ehsz0QPL8rVtxhMxe6CZ6Npvq+wQaMcGRFy2CC5JB0DA5i/vF1Z6p/1gNhBdnXea
lrAhuyt1gIpVGGMgZo5JVG7jqgcTGnJ2thi8RghTwBVLij52ZIjKhgy63q9lgnQe
/5qNzs4KG1RMKRVRbx/xNC9zz0Tumc2omHEWXlL4ObyZzhgLAk98Rb3B6Q1eC8Uf
fpEb/ls3yZWd/fUlaYlbYEM8U0b7cuj/2C3aPI+MaNOoFfb5PH5GkGY2siLrhTl2
RNiP2Rk5cayHBxisd1FJXYS8n9D8VEL7GPI9SE2z6XB15EgZmn+mOwBxpfqvIpMc
KleHUNuW9D8YtL5eCY60rukbs4MZzZ3kF6pWfZfbtcsCVXP24VUbw7NUMYVngpdM
YPBoFHlpLh7kx7jEydd0soMSy+fnJhEazSX+ORU66AlyB0qbt6LtZKzOAbdtcIQo
0M6ljyuSGERIJmeI47B3oDJLg3N9hc8nFb/CyTGotLrNO5wcVoH0O6oN4t2x33b2
OCd8+LLAYuWzuvjqmaxTZZqYeHoblS6FduF29ibwLBnFbdgi1J1y52Di7cJ0Z/8B
ktNIwZm60tkTRyWPGpoS768R0hvzmZHSSOTKJLQpZfHjDI7KJ560vM30MqXM/Eys
uP+TXoQWkjREPW+GqtKuSyz2WHHm/MgaVn29fXZEqESM04Ft50TAuD5ivnXgvVy/
dcuxkGVovAsuyozJVAcSVQ+sFCWKTPdNkIjaWJAA9IxzgJyCXVc9Bcfs3qDFaqTy
eKUxwpy0538iTILHFQ0uG9OhQaDIHo5B/kXvA9rMHIshvumiD5v7zTLPQtPGy0xm
SEoqRKz7+o8TgbGIu8fNinr+gapL7ah11SxUMVFbeTutXiaCRhXQ+BW/pwS+t6le
2BEzZkIGRoJXoPi2PqS4wBNGyxZ1MMwpgvvTqd6vUpOTtkeyVvB4SS16hcRrkul7
Sm85TGihKFatPuxU8ATqApHlB0eePvIkNgcc58B5PVnnT5/HYzs5TxVqtuSDyIOW
r6VPhakBqLaBN7ocINr1scWl3tSaIO8+hqNxo8GS6QilspUMgMPSq8DXB2e21q99
B7s3XjwBp/xnN/GQLOAJAZnm+/NhjsBn1bBTw78zPPAY+EjU5lDQB0S3N8ZT6e59
x9OGo1jaYNuIrGg1NAT4hZjnSrxTgENenJJt/gNYplI68M6NGoxYcZJS0exAH0P0
4YARm8rY1Qh/qzQ1sSIAsFOu4SyMz3tiQI7LarqqmCsXVjdjacENJS9t0nFQViXP
DSt6W/MzuTDdJEIjbg3rs0+cbfI+H19DBv4cSAZ/K8c8z7+uko/cjSggFnpEBHsc
gDMYBvUnP27OjiLGmWRQmNV4AViYGp/fc4JIGgs1Jlw0++qQsMqYE1jlzIcIfrw1
Xoii2T71f4FQVwPL/h2Oq1YEA1rddBlOnQOI5WMh4ESXm11UbDQFyREWGAreOX9F
avtkHRNieP0edbpS6mrHJfHt7IA25BKC5rQ+p2SO2NZ3oiNZT7KPQ2U0MGTtpFRk
J24Y2/z64R1XFvEJfxOXVFsGXxdr5MBLnDpAHfcRv+Uy6KMsubF4gjTl89HlCh2S
mzX0UIX8kKCKKbmybTnqfdxv9rHKh5DuzchHgiUm0fLt+v6cZ45TwI4HAe91cZzx
PNcK4vMcSZny2JkPI4XFfraBIdHEnyGIYFoRaZr0f6M4Yn5LGnaljVx7isiYfrqJ
vZq4LRxmSyJbqO5KXc4GPSVvXymPzIZB48L9XDZpJEZ3ZweKkgj+ASqZGtwkQVAt
6AWlqdxJ4QKOkLh/k0y/M+Y4rXxDZe+YET9sOhrXpu7V+QrDIeFYHOClnsFG3Mpr
u7Z4FxA8EEzBNN4XcXcNTHxKnaz82CcEKvW+z97prlsAysxR2MwLHmZictMHBb1j
c2OmV9pzXAUIfd/ERNtb0mKkmLS6iCWIOQIXSpS3Xju1J0VnwAYwDqwNXmoPYjVy
gSis/2nDcMLzQKYir43jU1vcZ39UX9KGSDtDSjDnMSrH9S3smR9smNnfWtsOUPGI
yaKGWzOuALjGGSzQpGZDj+DzXmgKxRcLVWM8GLrkoGa3WHTD2gg8/h0azfCWFz8L
tqLLMEkACujl3iwoHNrYa4Eu3npWiBTMIgmcqBSFTNLzybqebNj+gQS6QHZQq91a
Phcjb2tfTsKD1wfE/Um65pBPy48XtEpIxfjStwSwZRTXgvrosZB2I0lAWoNvphxy
107WRx/EblyB6Fbzz+QccbdOprh/91zXBIzHSBIic2f0Ej1E4HqEGxRrw+6mn+iT
Unfmf09gQdNE3SFF61uWgbY3uMtdd/JqqgWO52e0CMoVac5J39uA3O2GMwZ90Bls
VlMrCgiNrzWqWUDphROQMtT8gE5NNm3FAYiwSEgU3d9kz5pNJkfuubOLPZ1pg8fg
37u4XC2NBoKiBKY2+RGf01qR1tUSZDrC0tdjQ+lEZ79ltsiRtmrhaTl22Hiuml9D
oz+oaKTOrKA5frUpXfR+A1tSMziUCDgJDZIkmuep3IlOedFFIIzHTjyoCemXGoR/
uHGH+LeK55XiIo5b7IkFoOT1OalIj7fA/lgKyGRap4nvu1MXmLISgEK6yIUZ4QVc
0oDnavKHU0xfqVDO23gzoqVkzN+aPuw7ROllpP3to5g0MdBgsG7TDbt7kKayOKLn
H6WgEx76ftxJ1+PPIe4Av3TKW13hAvH2VKvhMphQUsKvKNLedLl0g6DRoHeTvDAJ
t2xLqLVvMNg+RDyBrsa/W1dm0xq1JE5rJ85yhHm2ycruFDxkZ5Fgxg17NSIkfRFk
FtK7XHQmT7JGUpBhU+/bVidZzEV1Y6eCTNSLJL3zIEgzPwlJ3wXwZHWHhJsSsWWH
9z1mYlc/vFzQeJ3Yga8/Df4ltUl9GW90+Rq6cuprwozuJIzFFuqiev+5TwngQ1/d
iLUZuxdkTmOQbpCNMuQOEYGldMZnm2S/4YkgexyRaJlJnqE7qZQHWsikAC4ZE4wp
TYOppIn3I17ESKn+AFZqkWtmKn/kcAqjJo5ON7VPVYdirPVjBcYzTX+whedReaKT
dsxtkImUJUN9p96rJNRyKDpOSYLuKcRrSNhNUTnC2ktulzbnhIqGntw4E0Bt2Qw+
DfzM8/rvgghaa8hxJZTD+wgC5S+wFgeDbrmRtyJCsxFObgcf8qMCERPrX7VMa9MM
N8suWU+yqULdRaUtXXbxQiVT/oEQyOXW8LqS/aSw5iJQmzEU7o7z2ZIJz8TutgGw
g51vb8c1zVE4SbzDSt9rAJRsXRrTzCbOW/iQru29Fm7jIFbKF2hlTqopkDZlNnmE
Y8XFsHWkrtC6Bw06ARs3jni6qBswo4MSwiQ24qVUai1D5vt26y+r7bDLUd4YY9YO
L4mdY7cyBCV5tSz64uakHbxjUyefl5t++vy2FqCd7mq+T/o5KELzFpOxjDJ1dO46
+n6LNv8aY5F7RIe0VlPnxz2ivYee6Q7/s5WZil/t4AZUqswYWubzfNzandkUw8KZ
+3TEYNo6wuTXIFkiyi43TTP5XWgw3SCWrPg00eEXM5I272iExAVFZ3ez74fyKtfB
L6vrMJYelCXmD2neNDz8kQwkM3xy0l6Y+4Rjw8B8cTq51FhEEvGtTjNUG53jw3+E
NcrTikhEnwnxkFjCNtqxHWxunHCQbHmG4X4YbUZ+qQyGwymBVQEXiHqtjne3A0rO
MADhqhQN3dsTRuiUx8TFUtA5F/UDKa+V08LP+y/JJ1odXXFXMI9cA1td4qTy12br
4oM9vsdrRSIXfgsBiyUd7a0Ykq3mdNwzCAqJnAYK1kAlyQUoJ5+Jf9E3OiSBfEVV
/d+Dxz4CQjvkMyULzhDwvO0M76dh7pnGvzxoQLDs1UHFyJVhr7SqK/UihieorvCs
x5T2Gv031qD/086bjj9+1CTkAI9zZdO9MhISAQXA5vae5CKKNwUNKUZtwJKdsQ8x
CIDJRegdrAkBnMe91HebextTXdfn6Bh+TlJHXgmDAg7MxGR2YH8nI7sQQBzRzitf
gCJajWACJJFO9oQyyiXM4iv2DG2PNXexO5jtVX2YOe9AGNk1RE7SGF6Q9kDy+7XR
O+ybkFOQY3e4AgzGpysUz9jv6M6NcSWn5RM9lhRUvr2rkOEMbcy1BpWV2xXR46Re
SoxtOM8eo5y8tLHgJuJHrW3n4EBRqY85LZMNs+IOiEpELVzsrdPIbbOefp4CHcXx
SEmXROSkAv+GdxwHXzcXbTqFv6bqacx5HbxE4qP+cMq6Xgc/mOqofS87kitZGOik
ukBkaPlsnrV1CC5J/7AjyDWSH2X7MRQo+oSLBS0xmAiYfZvFGutJXS0/U+OdMcmV
YWr2TJPyp9gafDLP6Q+4sdUSpemaJhFcNZViR9bmpVds1LVYFQp4l+gozYdbMKdp
U9F9DkHjIH4hmDz983yxDYlRplXv+N99jBiXLBwR/2yywOdHvetVBOifqbQvDK5E
ARvJJujeXUcW2nQoTGRNzrktpk0aGilTvevXSd0OGl6HZzE0TxtrJVJ+Ny19+1ke
o0x8CRS9HsL/z+EVdFoH+RX0ycVzLYNoLu7um6xgu/o0CawJbuA0+nQ/rLJfA+wk
rzEwQrBDWL+Rqp0xXUYvKuZh2LbJIcRVlz/kcaVhFPtfLt0u0PQ/DfWZ7N2X90zk
gTiPsbpWGXs5ONQmcMT1yJZjAnmbPBKufcnYLd/Zu5XiylS0L35ZH3CNuj/UpAwk
5qnNwHbbArpmCSwi3cvoOFj8MhmIaNmDWWFAKwksOWKPpH7ieO2LfsnVC8R9nugX
vlFdsjFLgilM9n/Nxgb9O+0cdHl8gtcAntySvAms8zHYX8m54tPqzzl34w4jGcxE
BEaHftkF0A4uhQ12piu4soDd7XrIsgTmArYPTDFMVYYZX3hOkZMMcqEGV/yVDBPF
Ky1vncIIQiSngwu800XtVQE2IHd6uHoPmcVnleIAgORSFmp02iN8mk4Y/4gxWSKk
54qnhRhEfodGyr4mz0nsJ16QAZYVpnLp0KCjpFQJ8g2dOb/GirUHV3o8P8KV3fDV
MXIZeqcVLE81bu2VLUE8XrBe3jcHTD6K3pjJr1TQkzFvfrZDyjYHaxHk2AjNk8mn
XsbgY38tCxsfM/lQFhaRsEk1EzRi66OwLTQMPvTNEjx03whKxFhY/RU4jx0eBpbf
hX2a/UyYC1lDr+JoGZWM2m8J/DLdLHDbWyMM6Q/EFi8LAm9eN0//H7PJG9TuRmwg
Zf5/Di7961qkyaAu8e7z451hItbFfZie0qj80DIPp9h7gbYVosqnG/fsitsNPOP3
gfD83DnZngarxul8B5M2Tgh0Vz2/tkXAxeDXLrnlLLfwX2t+YGGvdcanCgf81ajW
9fD2BgrVjMYtNKdjEWqotyjMeBcOibqSuUnks5BFF1ujfPOyEbMRKRmULMTyqPJx
XtL07K8wofIKjlj7RXE4VVeIW8Vc1amMro7/8pcpBib+d4F46fr3OkHv2tFSfBGT
tUoLaunU0VlR4gYfN1J3psxx0Z19qkzkfxSJCsBgFZ93Aes+QONZ5LOWxgrjiLIy
xR0pFJnPZDaee5bOyZNRUbl4lKlNDsVGMTQsgI0ZVO0x+g2+PbNK5EDHpbWzZynP
pxckFLkKrDWajFas2FJ+S+xt0S1pBaHQunLAKGdXJMbSqi3NQ/+iVJdEsSBUsPGU
57LDl0y3yD70tmJPs0c+hci5Zl2ZJb4EHB/xpfET7Lm9lQN6Pl8J0njPAOfEhWtB
0RMt7z5FJkaET5EEwnFd+Oo56Ehqnz8RzAIdHKybh1Ks1lYkLoQFjltjQrW5iC+p
Aipoi5pZCZ3Pom2v0R8YDfeNNvKYSrZ9bMruWasMUKjPhtsHs3oA1Q9++4KXmYOW
tFpW5UA+lp5QTdlAHLFrCsXl6VRKirbeKQ/KQrQnINgpyWEa5e7oY3OmoBzd3TMf
36WKyFdjL48kKuuTt36DHPG0etmBfCOofnkhFpiPfOwAs8vNMlCKFbp4ia0dfinf
bUpyXAqnHifsos+vh8ovFn3hYU85dU/J7FVhGcRrE3bDDlJUysAt96nJ7mmvpYi4
gGyKGpUzHs04k3gjsjCwPfdNgwZADcffE+R634/zkpXpcV2JAPFbtiulr5E+OEkC
WrjH6kVbRSJtIs10Q/mfp3XcglGAwZuKA3gnVwdXxH8rVrav6JSaU0tYh206RzNX
pN59C2qVb2/J+jPpRjZJl0E6cMfCSluMBYLpPKBVdzEmK1B1RGuq/Jy5D8Zmil9h
ossElXi1hz6QOzady11zPa0rq4PtZ44/8lHhV1smDmjO+TfklXOdH8Ci1sH181lf
mokmAfM+ins+bCKyDELJRHN+4UJlPU2vr+pb2hsbPvX80VsR9rndtiPcShpBbSL9
5JwkqGx4MbxBLbaUhXCFYuM3IJnIXf+ereN4zCvIM25FqpFetSZFJ3ai3WnIJcNn
LPoBgbDj6OqsoFqkg82czPG5DGHbC4UJ0WtJQn2K+kC4ZVK5EMwmJGF+CaorOY/I
Jwt9k92bnPxJuJ4hJNZrMWETfKG9ygFgobEJMfdb7UyY7bHWRZ5B1RD/IZResI1J
SoGXUDd76x+iVsrMxD5AIjfRU9k5879QIEOJhyuKkxMYcScak/exk9laPBo36O0S
GZrf3KzhVYcktA7tZ4OPaC4IdNncmEodmeNSAvZ8yoxHffwkDpR1FSZ34KibvC36
jR/fh0Ep2aH5TxDqg7OXiFqO1809wD3arVeSITg8GbjQJqUE9eOe2dPPF4gQmJKU
wEDN5Xj+6tdEDPEXqR8vOOh14/MLi1bBwwzP8C/qaIL4NOR3FA6okqmfyLcmxhyX
cH0V4xJCeElp7/fVDuwtiNHQOxtaDQT7L3FpMYK7QB3gaxV0YdHxIzXPV1Bc7dsZ
/JcxjqJuUf9nifVyu40Pfcxbg6CCNCoPP9HP+8Jys9gRZZ4McrkNNjctmI9Satl3
OolmwvAsC9A0hiofV5pViKDP0VRASOmt4O5wJ5Cm6mVgObvOBmjONa2djKjLb+bL
/hQxttoanY20jffpawfzZGKyfsigw5/JGcZ8HlsDvaSfxdTE8Z+LvYngJs5vBueG
yBDGzQks9NGfWAx5sPMgS1yns/I8xRqpL2KzqmG1q+/6ozomkcAh2k4Cy4TtodMu
oryMrMvR7viBdb+vMqKOU3z1EbX7XlWMrGIKV3siXf17ySTLEmmSuITt6vBEqHyv
nojGo5fCwxT56uTgPDZIFh9DZKNz46Ee9n0NzRA1o+fBmuQX+GVXyVnAYRUbRly3
ZCpuz5HEpUGUjP9vux/uFt9opgWjulKdRddFBIPrQ+UpW457xTVrzrhNW0dESuZd
wTUVxf2wbMLXRxAzMNlsSojQRgERlDjeunw2ukIzw5f+265gdobn/5N8JLKmllRf
IOo4kX8+p+6xNLTWh1aV6CzA1jFD7u8r2gS4S4jZ+WRPNXyAyqf8XWFJyXsniMXe
+dlGPUpVHSGPO5BRfeRirwDNZFRCO4w6eaijks+pP6pbo3zHYxRhMPESyI17lRvV
s+RC6avFaDBgiZU5/a6bKrls+RD35OCGXlbly7rgriTdXfwnE1QB6sKd6+qcHRsJ
hlUpp5ic1SeK1DPpkQd0UYWSN5zfCzvkDxk2ys9zAzC7/9savhHCuDNf4lMwpZXh
GZfasIj31d2RBZ4vB3PxK/GF47KYHC6iiDN1/TzlaLV1qbs8HUXDH1p5MYSvyL87
A2byQpnByocgbqL7qXGfYyBee0Qq79MXU+RRP3FLBBO33w+YJhsA0cyBd5wYzIEb
ub5Lqh6O9e8CYRY0Fkg18ZJ7W3tGT6QGJqm/IcSCKCNiR6gDAFz4XtEwUW+UXwpo
rXhvSRE6cq3mpsXEnU3uGVqDjY1YCGXnXqKpLjcvLzkCiVd+O5xywVjdPQ5cRN/b
nvU6jYZ0dYSDhwYXsjDI4FCcnVfoS4UmfJWrleKRUw18I09uIzY1SZvjIpjoIPol
iaWdSSByXsMaSial+SIe1wfKIKyNO/X+nkKuHCJRqUuY8rl0Yzc9lBuuS9lT+GyT
hj96P1sGHLakZKTFzQiH4uuOh/s93/NMtFCtprl6ZgpKdDwDGCUQILIW07hoA0Gs
7NFi7lzJ70uI+fuaA4h1tOaRcjw2G0jqlZ0Xh0lIoJjAuhynn+mOW0p7nHyGvqGd
8Sbqr5xLmRBwDmY40vLmwD4BD2yPwFRemr2vcglB9UCzGJfZmnEw0+Kha1OFOYpg
RsiblubJzW5EcYfcdEl1fdtPuHZyFqtMyle4drn5mjU4M4xqEs4Ng24T4M+AOJPO
K9xAh7vMS2eDeny7c5rLGnwqoX+9R8o+etmvy8AqKs2gEPtyV6sL6cnlMAHiDuMT
wP24PxFO5yvQQs8h6eXIdTehhbQH2+8ISGnCzZ1iBZNnKIYCM2HMoOVpT7NgPZoW
/NqZfNwID2YPZxI49jBhu/QdHVxedoxG1k0WVXLZf/kwxgvOaxOAwcKuqtAjsHl+
Vsv6qtGKfDCTRIIq11ZmgfP37X3HOK/ZAxLRFMpM/nNYgur0bMMOZ0P3+Yw3xwKH
9KiZ0HHJKULWkzqHWqfWPm4Cy6HLe/68UcyBUnByP+5ujmqpU9qoyt3zuLf8hTyu
m9z9fh26FA+VQ9mFzjiktbWVmknt2X+VH+JTv1FmxYGqN4u0I007t+c1iFJk7FKr
s0JeocfXxMtDnr32kz8RmKONwBEg+6MJHPKCu7Fxqclhm5FtGLiXLT1aZQmcPQg6
SsU7yeWJqX8BUoPure2EShYHU4ySqwr2taqE6zbYtyqHQk79vwoIQUB8t87KyFDF
Sx9XXcgi6NJMjLeTyID6v174ytCpl0MeEyNuzWDxH4hM/ml0OLogUNnO3R2x7ICl
mR4qFSBa/LzCt0kRJmxU1j7UpZPM/h/+FfJxS4/MJNz+95zWwO6KNyCmWmkb56VN
odZkgHfEICtLhBWlHODfS2iykxl+uui46cyXffyUxpGAVWjrpTXp6uzsyIusPhrf
G1pCBmJlQf5+FZY8lblaRLED1zLQpdYqnU40VTHEVzzA8FZQdTUFFDdGr1v4Vt9J
S1eKrz/wSzlYOOlLsD5IlS90B+izkeRzYVCDdflxDz6S+NWB8zXTts+VeTO0uQ1o
EV/PHn1Vj00ioJQIatqnZnpUhyv1KpkgajNCbhWHkHCoaSzax8LOV6ftBTuTVX58
nKwjIluJizq4heMBJ5Lckl4eh7mzQbPncj8r1nwYCWk9MVvj3WCKdSXJaBDW8UIs
eqpw896pnY2eHXZthoG2wsQNcVLJ7z1UfJYAvysR0sV5DZgB0x8NnYoAi+wV4Wom
9EUP1dM/kkn/kt0PahyOflNLZgT8NJxEMahbDiW0S3xsLfIHMllGd96I2eSm5KOv
w3ijGFBlqKJpW7RRnSN72wCVlkigbxU5zOwHGLR+Tek9Rdzw/hkyxtTmGN7QocZW
6TUvAVKieGJBgnuV2RW34rxMOS1KblscbnM6kuGMg+F67eOXK9o/9jWXI2RhkV/V
B0TjAnbZweo9AROy8hd8A2Lc0vAqNOVVi3P2FmVVcQ9oe8GSSUeqTkbbxUi9MUkR
HP1xsUJAKi9lRXIbNItQS95xLPTW9MuNlxpx6IdqaiJVlze2n/5yuYFx24dW/B4c
m2kofHVwbDErB9WSNGhxKZV/9hhMtyaiMzBZyJpzrq5xEgpZrrNFlnSWTatGE/zo
beIb5PcwE+a3s4AUbL80/cMy4EsexoN4HbsEJWDzB3zSqNmpvVLSm1m9r3f2UPDe
vxAZNHvUtmrKy33EgIy3KPs6zCDKfaApKZkxcPuyQPIT1y7zizajD+sO8U1F0Pm+
jKYAthBNfU6UAcNiHWVplJ6fMqxnTylQCw7XUYaBTbcKjwGviOVjOErkfIYZKd9m
Jl3uZX/rgQ9xL/oOt+gguO+XXcNygN06jjYvtoU3f6JbXWWlPJ1nmTYJlb1hUJ/v
3zFNJzKU2CFZkW+8Y7JNj1XJWRYEOgGb+BSdxRz9g2hnPVekbSMk/cifz8Q3LvLt
GyEmD9BLmdHtl/YZKpN3It+0S0U++O9aZtOjshQIEcRZWj6kxFAEv+Iwqfeby3ww
7UAczsHOVlNhWysg4tL1/is+1ipJ62VIYhAmM6YI0MwJHYXsk0qk6kTRhv+hvTvm
w2S+mrckLGkXBElZk9ueNag4QYdaDPGHIrBeQTpb4faMFaHrzt3BOr1IaGG+6iOJ
k2mgL4WSD8jfZK/UaQBdbq3FZwjZj/NYZjy2Hb5l3bmP58J1Jl6M3SoyOgdeS2mW
U3bjoGUsBjvIP+U/BWyMrYuzCgQezD9qpDG70v9Z2R2iG6/tA71uUIEwJM1ow+sW
CKzJToyFLCXlhZrAs/PFFPKXglpnX/FQZSo/1MuzNE8CYm/K1SN5MOP9Coi8NO4T
SFAJfOwg+VAWhkF6SI0Bdhu4o/ubsC/G4p/I7w/9q84fEvRsivMHyHTmLweY4T8J
GtD3kxYe7VUwdf7yO5o/syMSasw7aAYN8NuTehORh2PGuhaROVJVDdlylthItBCC
dnW/t3w7RSX13Gx6d5XT4yJ9x2eGemNM8Znpj2RVFPWHhWepKZX8Hd1q/LMFYIld
40XtzWU27uKALVfjObgD0wb8bkGCdadMMBQqai/ps5guEDQKwCiOL385O+aY2l+2
8bTPlMwbuoJ29fCt207gHSRT5yOAgEhN6l5fe1Lb4OtZNTfHOwG5n2SSyISv/k3I
pYS5cFZEBeeTmGrOiV9PPbqrQUrvTUhPd1ql6TIMgbh31quR3Xy1uFmxxxoShvAo
V9kQRk5vyFUJRVj+/n70L3zDl20rA6hnvmrwWhQNCXqDUz5MBWp4AfbrmyKuY337
IPPqtdrfoouM2m9ZCnC4ZY0strIQZzFCPtg/RlwhC6s3DX5qk2nM1DUoYXxX2WwH
mD02g0XKoY1Lbirxq9AW+9eWd4REXpNjemE318+E1PTKQKGnLaDAyIbbgwe9yrWk
peA3kSEwrrFFTo5wsfCSu5SS41VdkBHqDmq7V/EiTzvrZRf/sZ+B5+UN8E2f7AP7
S+v/UYUFt9YMFJHq7lgB+5yAz1uc8RJ2+oB3F74/EHT8Xr6dg3basEK7MRRgM6OO
dwVQtOvQ5IrtjrsFU5njJZj9k7Ll1vWMVwwiSdopPzHcvzgON0OMnpC0JuE/86Kd
AaP64HzTFYAUcl5bMUtKdU8iT0DQzX6UP4XBpGnYyEdJk+2fvfq7aBVjWXdcBjA0
NLIGHroA6c9HRx+wGm3ZvZ8T69wjLh2eKMScMjPL1apjQWYk+rDQmKmGt0LlZVL9
5Trqi0hagUPCgp2ZPqnvfRn78P8vAdZmbpLWfvoofue44IaPhIYvuxgH+ZAreg4R
uAJ9MiFqlwE1AlkGsCG8m9NthqJVFuO+UmLtJrDOkF76H1gFtaUYfsOSbNJMZyLz
6zJtM0WconE4wD7YrlyQTthg6Ob8a3HiuOA5EYqEOTC9WvUA41ca0wYqYZZcpbtC
h4haQP08cVE0YXvuerV8DaQDshNNSWCpuYsz0FXvbEslGJu6eeItLweW4MS13g3k
AseBNWHPQaSBAHLJjqvdsHd0CQ9EKWQpdh4cXzmeC7xuWWtHJrUY9JRgbLZbeWc/
JmkpShVpM72jMZkmdAn4qVl79BQzGAPWxjyQIIlVG7+sKEWtPuf3k2gRr8oqRuu9
OEzz4sd7IImfBsLpVFi0OLpY4/mtsqsZqPHWkRQwfUY5t0a5QnnMa3uXyuUHzlQD
9nOZ1uENgZbAqEkdsiZa+yt77d4hsI6bRKBKZuByc1wlcGUGJN/jogi81VvGJ98n
MT2SpZKu1gfB4Inj/x9OdET304WykADlD4WZXUJvE1N+ZFUCMp9opjpeketWlS1E
57mYiENSM7eQgqD9ac/uWHx+0yb9zKB/h1G/xPGfmvlKZ0+s1AVTQw28g9JUdARN
NiKjSiuOrPUyG808tja2lnWf4wK98yFTp2hd63qnwGaM0k2pAKrCxQwtDOtSdweP
LmYk38H/8b9PWp0Ce4pn2Q6CM2pH3i8d4t6oMefp9wf7S+11JAqtG93R5VOD8YWj
SZ2KPZjBuAqQ7+Y4l4XvBl3SB/MJGc+8PSwNnzt/P5NsnG2vSOSM7jjff5d7/A8u
o7i/E66YETW88TVDovgoxZ9Rz/zrH8yTU/2rd+Dj9QVOsHReq321hj6JrT0ehHvK
F2EiJcS8sP9D5owkyArT+cunfD5xOVISulHO1191tfUYzNvJCvHj8IZ7B7GbTf7v
0tsL08rMcqzOVvX0kfhsrka537Bmu9xnQ+VMWeVwBmj9RKi+2uVTnex5yHWGLfdk
TjmHPEjXjPEGz/01hWVSINQEf1oTuhiJYYCLw6MekA7kg+jdR6yw+mVaZ9+38dCg
YsWMLpDQl1P6uFIrihiwtCCgOSADD9oaJSXUKMuLBqa1SUAZuqqll6q9w3ilYQvJ
ApGL4c/N1wg89VD2UOZYJb8q9qzRR0GAo46op1G2aOznlYLGuokysDoOOvLcjieD
vCyUC6zGFdebd2p37899ClcK1CMEOVQlBZVRu3LuWu9cVkzOMymNntEnOY2Kukpf
C3xz4f6cDAOC9acrcAVLWb7VoCZcxIKUUtwTtOL+fLLcFOXwiQirBg29sCugtWCZ
fTcxjJbUKShgmYpTA+h/nS8dfPehEM+O6iEe2ggZUzDxLaAJMKYTvFQ+k6Fcw5Rw
SCCy79QqqAFvuG8+P+yjU5z9Q/Xo/ez828DIg7k4WK1p2jntPjAXj14KqkJZ5Ypa
eaNZMUATyc7je8qXrJVpJpe8NNWjB/vie4QnuLrB1FCc8A3Ai/ggVZS2ndRtoq/j
LHvrb5wA1lLVwFutJRvYn2QmSs/oYx1o0q26bYJCLyqVCXXswjg9REVuHI7vmMpL
lRN6XDye9RyaqOTs7LnRN2NmBIGIVQfnC+5aBNViVZ2Q292lG5uCz3jNCEEYxKUr
1wB5w8qHgO3zqnY9nV1Apsz2KRWPjCb4v7C02lUzWl4w9hO31lazt11TjhVkjV8H
26iup+ZeB6raOkgFzvLZnbPIZe0k7nZoHzcswfyjDyiYsY+AMRAEuulYfF84hMdr
wfF723Izy5U5igb55LtCMU9qvQw75rMWUEXy1/L5VPBXzJwNiMCm44HUm2PmsOAW
IJ8OKBkct6Vg93Oy7qLtAjnJhhox+MvCR4tl8RiPJW0uywohyVLSBOd4J57aMTIN
1oOdwq46Yqgtv6FzNt+nn6dKHeIx/6mq4NHXxYHmU9DSgJSJWlkIF+v4HNPrx7LL
kud+YUGbYlZHLdhe8p78ElZRnV5FHb6/Xy2ZLezvwzp2l/tqXAuU76yUxqylqrZE
skLW/+1abLUO3PILz5NyDXBVbExwuQtLwr13ixpd9CNbQNLHXUoRDC3iSS04srOT
ZWap5tmnpQGWg1H8T2N12ds/lOj+hrVe3p6u0l36iwGlZLZNfN35fBGqfsRCat8Z
Ne3Pp5jwLNB6xIe0vwxT/9MhZTUYuyVOCJvIOgeSPLdIEX5Nmk2MSFvtQ+WSA/yN
8FbOtCYCcv529Zo/FEK7tYYDGiOXK+lFlXBpYvJGwR0SMVcYGIBxwoe8OQkwbQ6L
dT3Q3N6vX/VVUsuuoeMcy3eeME/DGYdcdftynIeGk1ttTfjri0W2HviKoVQLrG6J
MQeT/AWp+x6hWUxQ1S2LpcpkRyFKY95TTQSlChUZKJFoNdlRQmbhzDEofvTLxhGA
wEGf8DBxfY2E6qWx87RSEhzNlbd49quhDf2f7v+ZrRXY8pT7/rmsriOFDGVo9Krf
cFbiDUp32xSE9ZkDJ0IFjGLGFJuSBL4hz+YkLgXwfXX4eHpQsdVfvpWmLniBYZG2
kbdibyXuxurtBKrzKr/Tn6hPsun4e/fiuJbCmZ+r6EAORJy/buXXKXjMpJPqnPml
BHRvuja+N050lyq5BSI3WLZKaGDYbXstBlkWGY0DbKnNWpA2OCIHgR+Err2ZwiY4
ci/XVKdXM6mrNezQLu7oCjXJNAIqu3a2N3hgTTvAc2TQ4CawGq9WvBnUfS6M/XiE
t69x+XKmLkPONr0s2JMnJh2BTP7Zu4MEvGtMU9Db6k2svrvhhMcIjRH6oCaVO2vK
u512w8mTjDPENtQJcOkheEYi/0nrN2LkCwroI+bFF9k78dsdKkjeTylDCEwLz3rP
EYorYwtMv+sIrPtIijRc/IolUrU2uE9DBuI60x137pkM51IclAOCRRR1Ha6YvbDE
C8CQlUIviXssRk/xI321WO5ZeBR8O8Yjz63DNV1O34cl6uSD6P2xypbMgwtU9Gey
FLMfR5DjfPACX2sntR+yvqhcyPvCtP5dNBml1N5EfAKlwkcdRdA/EktxCrulyhFk
KPpquL4i5E09HnOmU7AdzgK2ix0txQaWTVcDR3dgD3fskm7sqWpcxtOdDIT0TnGH
nLIjIHs9KuVcQrPf0GZNdFUqFzWf0mo0osE/eVfNcG5+JktboEEhQlG6MsKCi4YR
dd9nCqst3bDzCLv6cSCljVa3DLt4Jw6QX0xZhob3lWz1beuAwCF5hrZm3wccEvCg
/C7Qoumxb5vI1qcbvGlTT9q13uPYEvSAsHaOrDjpDCBBd6iqtibch0TfxscxTrO7
ONYky2dVonELoyEq/PXA3MMku06Xv2WxvuSRdT7hCXu1KD7cfCHDljeYgbVKRqS8
7SockNneWPw1ROpFlgVfz80tqsYneHju80RmdbSv9r8YEypOfxKRMDEFKRO0NZzB
A9DLe31mg3IWstqDFwx9Q+6qaQzOFbkEn7NB/Pf0BMuGpU9DmFnACacex95oH/kR
YhFm2YvkN/hTY3dEO3cZjS6ZlYrZw1npDffL2acEr7gWJk5V3IERH7C2zOR3ogD2
+8b4LJQijqr+zXQX9kA86vxN50GlI9k+0Ljc3+cQxDuNOjl5lF4pYT7NG+FEC28h
QZX7PO6L7Q7DQYiERdihlSWyv3Qhma5+Y+gM8zK09B2dX6CPvvZZHIDmEA9mAVJA
crGGV8GrvjedwN9X1xcgsihJuJqAzfauXgJlm+uKzOsBa281GVTuIFxeQoiCrQ4q
IB7z0ungJGc/ki8Xem+9HPWvnmXUUaVkYVJunZXDtydJz5549Sp/N449N6T+5qsJ
eyaV5r7aIp4xV9prUE6wYN1Bgsu3VA9HAMYILfUxTq2sfZJln/naRnqS3IR/ubU/
lRZVd9BM7oi/8Wu0zf85uqYyKNhN3nxhCh4igZlivEAqKboXzRpGPZTEJh0dDn5W
2rDY3qbsywY2pJIaHIeWqSFbF7SAGbyfuBKvspULZvlYqeESElLQOu0utzWAhZBn
nOvBlAplGMsFboL/dQGURV+NWH06T+iQPsI1HjO2gTNa9RCF1kvkJJlAOJOBg/Oq
m8qb8/nsjuk2a1S6L9UWDo5uysVN1Dwr21do3qbpya8TC6ek/i0kBfXgI0XTsK2V
GZ1W0HDBFGNfyfkFFjQ54IGM+k4rIMg/ssmuOFeilzWkdyfc7TkyASZRz37NgQDp
ybc5v7fglVL3+L4tM6nixmOc5BsCTAHONdwXzX+x+QceSseXVowtTJ7HhCdDCF5h
xaW7qY32oPk7Kr38hlSZyeuodh8c5azsGZZLK9pXBhQbJLWzLSB8i+kuHAIYfwJO
m2N68Y/elFAk/ra6qkvYybeIebwhTPJo/2OyzMoRbSnLdYzleEtPfxiPwIQoEOgY
vYRKL/JDjlHNoPJOqvDiS4u6/c/jGtYdlVzMcEm2JM9FLn13lwNTm+ZPT5LCTxnA
/r95SFDbFJ5W3+InwJQLbCT/Z2QnUCM/F0FlG+z/oiB2XlGumOqi3v0/VxzHCbqC
AVFkl15t8xNpeGVYJ2KZatUya0abAjcfZYbDLTlUhj4E88lFFKFvA2gqSV599goo
5MUFr/oNwhMsY5Z+QaZx9wK3Ud3vwKAOf0X9TI4N+2z1mczjHMGlnC76UNJvbFGE
xPRkVG4WCQnwbhjhDiD/xkrALDWSEJV09UCs12hSG8mMB1d8Hr1BPoRWbph5Nzm+
mDWRBBlpPT5gANLlsOuHFCo0C49yZhLQtkIuWgI9wbUcBulNDkXeqd68D5DTZcmS
zpgZ/4Y1vP5L51+E8rKgJmmYp0N7PN0Vix2vSYzHESNdvGoBuV2CfuQHAthPgDll
Cq3npRqzAjYw2Knt9RIlJfnOwms5ypPJU6FMKfvds76q6JGs0ukoxRoOGfjClNaZ
hNaxTYdoYj/mMFuw20jLDB5MqtIKdIQbA5Jn5A+IWSMW5F+wpiJu5DS3ReZAgCJg
lvhZZpgWh14iq7rI5iWPIRZxGbakeoY8WAZ2Xky0SygKiIuWdKG17kaOnkqdWTv6
v/MHOa7jhxi6+PGpv5Rbp1RfYQB8Tw0OLOpcfg+hbA7cexmQ4FJet7lmsWqNjoxb
Fn+VWnxSU9lUID2XtyeYsGAGBTZQIrVj+Ha4BNkQbmZYDgY3MA+Sj0dWu4+ASwOj
dDh2xP3oqem4UnyphTZFkGW+3a3sGtKiNAjLccbHuy1nL5SNyHCmqNZ1VNa87ghR
8si6T9pyab4kXhT2yTwqD7uZXmylU67P9hlZLamf6jpwO6udrFjmFhIGwlXZCXM2
xFaq3dJev2o+AGTRFtEX+OBLo5i1RDRZq2sEnamObH6AB6Fo4v57U4ZkNslPfc7x
sA1hVblWzmKviSUus5JxMxygEJsIrn3wLO2elPJbPqoCaBOotnu8D2sOWhBBfung
+jLAKNn043+3IS6GKmUQy72PRsxpq/tdxE5RnWytEzqMOIrDmhrzqIuXC9uwGJkq
CP5tmMxGlyxEyiz1xsidPnQPAqv9HWk1Csxblvm7K1/EX51hjzxZKsW/qcz3iyiM
077df2cbgn3oijsejsksXqOlVtnqgw+Dx4XZOzJKZT6cvKBQA01P+20oGDunaKaZ
pp3hFHfacleq9d8Ixjl72pYvKUhHlP6Y1pvk61mm+K5d2UFXZ9JsyfKl0FWqK0vC
m12nEohzj2xI3OgKVRnaV4mCO2r3l9TBiPYV8ezRrpEDSk8tap5IO4lQdA4aMets
+hw6lbsFgEZA+7U11AfIuWx+1xtE6I0sLNLZyY/rkCx3DEhK5wh8V7Da5nxyshO+
H6ls8G/Gdooa21+iwSudfyIcTlaBUNzXTk6JaQroQwY1BWIgdzyeZgH9MskyZoxB
MnWxD0CKqjQDkdcCNmTgw7OQ8HPW+xUG46mtUDCvRiYuuIjqxkerXyXFdAHqKCcL
frTFGwu9iW2oplCgOWuM1N3biWD/SxPetHkztI86+sflnP4VWhhH7K1tfQHEaYBQ
eA381NjvqIwrTPQ6nVyY+VtfZN7dx25GJiLbldL7om1nzzlZTBRDZNZh9WMs73yG
SQBzRnw2cjBZvHvk3Xr7ueqJ7LY7kstMBQ/29U0/aGsKHcyUBglO9QfRBvgMuOha
0O8cg5yKSZsMhpspsi4v2KoGQRLlcGJCWbbvgm9ABePSzP2cY/tEFZ1hxJAVo7Qo
aCdlnu1xw6bid4lnYq1D1aL4hVjg6Ujrl2SYulqHFs73UQy2dVRinXaXF1lKZ+hv
1AXAA2qKlvNYunFP3eZDrnkSF18XGYwS9YOHrLmg/rcljMFTsi2ek02fnPcWe4vY
crAHTnMPVBGJtKZKYeWS96ZS50EQ3kJuQwcpAeKCbDWd/6oYUy8VX9hKpSFkm/uX
AC7mIqeiTKV50o5RRxZwmP46CRMF0Lc4hwactwxF9FMlg/qS0dja4LUS04/wFn82
yZN5BAwqedlpDUawEO2sD1kQlW3uY4U5/jGWDsPm3M7NRvUM14DCecR9hSIxmhzk
Tfbsxlbh1FYrbdDoWkJTj0vi6b23377lWO3C53kzoqqRoquUgw+mCAfP/sMVDBgi
qsYPh9/S7PgBHDUFRRTGGJ0/uFApHNn4LGZ+X/ZodU/ichjGe+3E7DoKDVS9Voyf
t1n4n51RMo6TwIbwopZChGUnWS3VKTy9goNvfwmUoQEY6wpm8PoPmuJfsSPqKYeU
TBYZoOM3YnXe5jiGSl3oolLUXaIBBJ/wi/f0St6W91xJtFUkYwY9JdIKqfyhNHaQ
lHCmbuOtWiPnxX+8ABCJOUH+qt4ptDHNjZjS41rOuIw2FiOV6skZr73ALJ6WSGcK
kjX5J6vL15iC4hlvZKXuOpKQGh1L6kQEyiEIqSa5cGA=
`pragma protect end_protected
