// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gj3orzPAr7RL6aMtkGOZQxRzPPIY+ZtnzizcNc/gcxz8sRyeNk5xdUL1VSNxN+5w
8cLPm1aHWQS3HwOlzYZaFfRN0oX/ay+VxSVlyI1jVp76g+ADOpb2KIo08nGqJTEX
s2q6jcRUfVsTijXwPejIQA39Akb32U2a2EoZorFNZ4c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11856)
kD2/tIUOp4NOfSbMYWUfPkSz6J+X5TsxX2pXtyFvhcLwb/jOurHGhviK8UNAuwLg
RUNMGQhHdis/PWLr1am6wR/krteukshWcO8ZS2UM42MBmuVxVksVGXiY7hwxrfi0
cHGG0FEAk7QAbWelUXiDmq/pp2L2etj5rJGEp8gjx392yE7+jY2mP/T1qbLuhB8T
lCd2veVKa1/SJvWr/eXPopahv9O/36/XPWNKk0lxE2uzHZMY/F/7Sy3wwE268gfV
hAIfUDDGX6IvqighRxRSYbY1b/8iZruVRC3NB11ImrLqtSFI6eYyuAUBKxr3oHzI
O4vQu+mPirPz13QTYBmN0A556C5d3SxNArfrwiDsgV7jQiG9TvVXMUjav/KZVCF9
ThY08F1LXGzN2ZnY5RcwVbCfPwiO8ed2RAavg4ntZM26p7JhjDg0n1astvVrp3Su
YXhcADZSFaRiepMow1JVKfystX1nPdKQtWPKClJMpeZXNRPjsQs1mR5qIpwLPw/m
UDVr8hu0E87bnsLEi0n7mE2gsW99VNe8pLBzzCFl5zN/lPz3TO05fAawNQczRaCm
gp6Db/nUnUo54UGyLjFzcxQ3d73Jg1wsicipx8/UUhuIc0W94GtHTDWeX7wg1dxG
9hbndwZwBGmJx5L9S4AgT3DieAxHDDJOzTBReLR3zRbucLIsaKmRiMOTLxGvay18
5BqXGtSYqfa9Ace04f59MK7jKwU45OJftj02IMzsiIINxYXc6zn+FcPbMkFQQPMO
gDJarD1SWiCs9oIqcnBiho4duge1rm6CAVUvkORoobxrZ+2ICEYtjTNob3IKuxap
JcgTFpPT+sGxAkJYyGfpe2ctjqcb6TeV8xr/+tQwePOXwb3KV7rc6PyeQkSkz8sc
BzvsY7FNrfDnukg7FostHJkHSxksQjXzcfjG9ZP4WM9QZgdsznV9VKvAjtJ+6WbB
E02s2S1EK3BZfkk9n0b/iSG0+foZ9Sqky1mZrhl2KWtnRiiw/1Ooxt95hufaGCzV
WXOY65p2VlqCcbevA4/JYBSU7i/UCR/9Je6hIcBo1rsOlrszZ1JvZAwLgTNq9ByL
KfC4sfiGtONyOjGQDiJ9cpouhJIRRkLiyA9470VGLEnHV027e5qZ0lgVp+AJUzNK
AK4NDufgHLFqa8pKrDA5unXfHlJ5uq1aUmDIhgmt1CXIRBb5PimA83jzg89CaY4A
kz1lEpnHNm9OH9CG3LCyV5Y+8pGKUtG2wcrBer2wMeC4yQvYMNoOGqp2xE19xOuq
KmS1ZuRoaKOv4K9HdnVGapFWRJUwusJEbQjRAPzf+/QaaVwSuUvoakrIJxkZPFW3
t4Ykw6dHPyT31qHFe+FNWH/QWgkZ3ioCuYcFDm7PFtpMwPB7xywiAioeABCbxDOc
sydUYAa5TVxpPQ5ocm/SNq+FJsJmH4XDlbpXjvABK1VRq3+gX2DEpW+UV+GG6alu
xiz78QveBXAMW0CwbTAtrbnMsuGKSzaoqOWyd49U9t7Mjs8oUMPBI6S8ipe43gAs
C8ReencW3lMJhaG4Ma8OjS0qAMJKHvN+fGM+Ai2dXWoJU/UT0CH6luF13nbn7xvg
W2ea2BWnToxeHsRSLfQ6Bt88i5P3+yiyzAxA/K2052slFhmX3ospN4HQ0YGb7stn
cTWNB32wSTmJMpxP6MKD6gWSRLlvff5qQoHYNMzLVyGbdTpZ0VrQ0MMZjz44zRb0
V0yAcn+clPmyeP1QRTfuYzOb5uBAfz2q9pM2pqo5c4u0O3GY/092CCUhALqcCBDJ
3+cWregTjWhf5Y2JNO6hcn8LBBdSr3//+1fSsz5aT0qviECSL1Lq4iw2e2ICKo0E
0Vhy7jzAIjdLPaq2tjQdngh0FZDAHK17dcykZNY5/JzaKYHfVY53UgySyiVxCK9b
TG1iN459LMyrBQstnc1+zCFe2msNWJMgPRsGW+52JsnBjHFF+u5KDOskONuHS/+j
ucBT3OKPC62IOswTdWtaTx+JadykN9Jz0RBNn2NCRACQtcB8LnmCvjF6b9ZL3x4z
84Rm2d/yOrlOmR7M9QXWUXQ5fBqMreKooLbMWBEbe4vISP/KoRwqwGZSX9rwaPl0
aTpoFSzqCSwLd97+AU6KwhOWFNb4Q9p+e1D5ZvDwylWUe/p0kdIuZ9uYt4Pu1yLl
iM8WeMqus5DBW7k4ZjThfBa+U3AB1jFnwhS7hLWGBc3dU04m6SzRFjq1zl/2Vx3r
rbQrHoz3L1sJND7GfASg35VeK7fv46uezA5/2jOiB33kfR9ZM4/JocfOuQKEyVam
MExFRJmT+fiITI+pOzPexoPnVowfB1lQ4EP/eAjQ0gDdD2BX+9fnYKYToqGEgHZz
i+H6IJAVob3e/O8WqIAc/1MvD3HKwE4p0v8RKgIBI60y9+z1vRKg3URBah9wl57s
35s9vowZeYIr/A1a8uSsf8iO4iCCj6Agssj30kQshrbLB3swmbYvoUhtUBaY3V9m
Xzy2OwlywHMoM8HRZV14sSsuaPM2mot5I767UXdMVrMzPJlqtZ/k41yW7z2qH4VG
4Ox3kXNiD+vX5/Jcv8ZHe/mwg+9APAmBpyO/JZGgCuAQG6SKZVVkgOy2C/jUjGTJ
6HlTLPOQ1QcfQpc0r/+cIVIVZAQXkE7C+sB49erZgPFOxE4SFmH3bAe2hqL376iX
RoCgpGvrSmDhQlJVdlGSfZ4kPz8QdkHgDgCtFDCSXqcYcWthH8at3Ol6ncxCtDyh
oDmiTIZm9V6mOFidFxZVrM9/P65v5jIWBy8Loyd4FU62IqEl56gz6Hyms7P5F7Wr
J1NX3yNM6PjGnDxvKnDCMdGdvp+9xNh+uHOkrUbQ/lgyGsvg2+1MkJh2O8IyiQ/a
Lr1U9SeCJuayeKgcBQXgCQIW6mgGrCDXRJGv1nRupbq5rZLs14qVE79lUPlYpu5w
U0JD7rgN6Pz4nGRpipV95xsKL2sXJvqGIHJeB/GiXOiLqL6qKaYGvALpD3M01hRj
X2xtuR68qrXjIXZfl4WfndCJvtV2tcOSy6elUs99MDIBM9Jq0ID0E/N+UqsTjgMU
/v14vApCEriYhJfbWuZ9ZBbZYNu095utdxTRyZXiUid7Uc4B6WAB3pXbvm9pICvL
OguoSXrS770pnh3kNZhyNH3//dx6vyrSqzGWOHr64HQ0OUgiGsEPfSuwIFLMLHTB
zC6+PaTmM118Z1ic9R3rjZTFmBCm4mEn4nUnHZDQMXmg9YEO4mejIw/Z0gip1AW6
GCVcq3S2gd1JNaDEX4bbi7XHAyFO2R9LGFqcs3dZJnhnXtNZHDYLvIGnwpJRMcOT
YPH5qEPjo2C6seDLPviteyr9NF67H2nbEcm9Getv0Mv4dNXr2DbQ2n89rWr5FjX6
nHsf3u40MuSMYCRyUXODrEx3MKrRLSuLk5YhB2sKk6/QWOtaBRfou2M/skebS52j
1d2VkXc+LwZV0jBVTQfAEUsH2gxcwad2g0R4u491EU4mAQYzOU318pYspCkxsgU6
Q3amgwoZOZMcGoyAOaXx1xRTir1d2wyl/i4iqS2OmabmZUfpPGRHeStxUAyUdINd
0PcxyF2ce5mwdlRZ7//6pfB1OZJTls0B0Gve4K+rJfwtbC1n7CqRXRHSBBKO2VxX
/aG5x/f/KPGC0impHmhU9FfLP7jUC/wnL82ae6Bcn4W1ADKuiNgsPJTi9P9Cx5U1
bVMXm0W7AqXEn+SXZAUnsHym0Hzszb6vhFGVyctlfP4eGLdUFpduvZXe768qqVtQ
UysHLh+IaemDLJZVVWCXNmvymZRNTh4pCGKZS/kEAQsShaPUQd5xau1MFDzz6gln
HIUij0EynfhivX1BfB4IJZq6zFBBDKD2bVGQx3ZTO2PHqVSzC65d+xccsxT287mB
5z5D3W/9VWqA29mqtVGknA/Sm7zXgU3b41yQpt1uNjCHcfkxEonDpaRpqwKYd3z4
Q6tgx54+nTJa2PgCYihtNk3d/HXUppp/tqhLqzO06hSnh9Jy1jvTRQBmxMsXMM/z
CJ7P6TsB3Tz2+G9KSTtVIUsBH77iYnS4wRz8Op04njRVQTMKHNxfubOiIL6EUplT
uXwWLDduYfXN4RRodUau7ZRaK9xqFs1vcbVbbfJp96TjdnF+WUT8GA3Iwhm7bIQN
1Mmqu80z+V3A1slamrr6bS87NGVgveV0rj3wREKDMiQjn2nc0usIywvsPK/M5MK9
8DMYxzt4swHIHXmWzO8QPkcruv6O4OrHLUdJhHCA3d68lV0H6sR9b+yqHhBlBxEf
+OZQnel3P4aIzKGOKDxz7jyln5lw9NXmcly/bCJp2AkgjEUIpMHz5VHkbJe28n9A
xuhzf6y98V0m+IyUKT2wHBo9l1VtpVJhWLHo0RS0HS6rdzddxt2Jh9vKfJ6NxYe0
ttKyp1MspFfyJkelIi8aUOpJbVuyl7w17219vRDSCLWHo2Bl1aCFa8/jO8lbMfve
I8LujqYPaRH/hP5Rfl6jLYjQpwP5r5UioweMQADMtBEymrXxw2Aup/s59YNlh2OK
P+AW6HxFWACI91hf10f23SRC682E2esQzZCbSa0HUQ/0ZkpSarYJwX7bkO+eKUvO
F954NjP6ubqf+OQ0AJX09jWBlh2rvWX8iwrjEDvnAgkfNWDTXP5oYGlaGfrApziy
lFx+eNKRpV89pGo8YMxZN9zSUVfswdIr6qlvOE+RPxYOSncBXDIts+EaORteX54z
XcQ4JHSZUSQ7JwHahD882uyXtIXbRKgiuEibzEnQYb7Bhnbzbr+vHyaq1619m10s
dRcrVkG72F8aNWXoK7Pq57W97PrZdnQYWz8Zc/NxVM3tA6XmGbdB63zOX8D+e8/a
GoF/jyEbRb1h4pRbpjuwi4Z+XhLKYEGI1C2eQ+LB9WNSLHaZzeb9JEMYo3sWu2m2
h3381f+xfse1bU5oRJhFdUUFwr8OyJ9uq6j0wbZl5fKQ2yNz8LgYqTiWDR2pQh5H
gmTh4uMfrpqObr07vynt8gUS4QwufhcCYtPApdH/D9f1PCXFQ1FQbWhHn97fEfrm
gtlWUddpCbV0yHApQAnpYjGmMn86VgfP91fJ8OyLYX10deAnWJiwGz0RGH0oNR0V
taq7hMN1cMMbpz1yEwD0XHP9xNVSjN3mYjaranPHdjNzyiB/9e/nDtdvNRpFSXhO
86fRa0JHBRrxjE+JyufV6BioDRWBjbUN2lpHAdOSz+8EChSZbpnrqAQ0KN5pLvJL
onUL4eDrlhmZSNEfFddjP8jJpCQzLOwVsQ3rfkrMqY9NaAIE1S5wLoqN6HZmtv+3
g5UZ3CqrRx/bmX9CqditdmHmfRjhJ26w+38nm0TMqg8oxdjMCTO2F8ZzgAdegNFe
IV7vQl6rcSvRFadIcEnTB/GGF2eEU0O+w1GNjwfRAvZKcU2yUdAbuTR31QNzjLI+
WNSN49fQaX5nwGLmeKs6+v5NuJ6I8RGAHOJHVrZRfu/1sLy6bR7PPmZPRvAzb7wz
79Z44cZwJmzvaS1xFVsqSvHKCQXc+Qdz96tLI2u0a7ogv8AlJlDloXN7eovZcFEa
HDYWfCVfJ1B6LWpDTmVChayBDMcV9oQBgNKxj5aV6xRWMa5Ev+2dR0RmK1af3RNH
NG8sRLsJuGIbu+5akXu9jyQhe4t7Cj1z0YyjV1GUlMTT6So4WWqi0qi+HMd1lKFJ
7ZF3YWoEigpcZdUtjoOydg+qY3nstJmQ4xPZ2OCYeqaBRD3xzwEJ34FAP2gLMOVa
PY53gd6EQnhrCAeokc9ysFE9qpD6AMY+iU6RKiRntoNof2S6fsyC16GhtV58oSiy
I8+YQdk2wQSLSLoo26tQl0zNhRR54BazZk44voNjuVncFxbnS/ilAfJLR8oww8Z8
IjCyd22pipeKVkHuxVlX/NAK6lHbpTL/TWtzB/Pv+87vEW9fyXkfYiCSJat7bDks
zPbxdTOlLnj0aXvwYSMfSqyFAfYC8sHSdDXj3te48Jn3sJ9GkEQAjtGBF6Au/yMe
jagw1iDGLWjb/VDSOApjeIirIQZJ/KV52FQ/4yCiMB2ZKs3GhR9YSOYarmFItPm6
0zjELsq6xxQwnmdrbROTqwRmUsyw0GP7Q0uc+RbwWTUYsEj2QX1j/a/jlka/NadH
naWFM1yPsXIB7+yS5qEy7+knxPbnwZCWGkoxQgaanWoNcQWV5WGwZW8Sc7stCeWm
lZxDLKHeV4nbh9y2MTNZ+bLKKjIrOXRhyS5n+MDsP4u6qa2mYNJXYQ+k5VfTKKXH
wWZO+Doig/cfupLofHgpyHBFG05w4uccwo+uecphRIZh4vJ6GxOKPdmqY/a6js7+
fkcjPB4TN0Z2Y5L62awJ4kVhXdgpG21qtlO4HvaojOJCMDrU3djBVrCkcOOvHNAs
2d1Y4TwXW8mkICdK4sz4Ng+/uJlCnh5Phl42UK+BkAt1PgMKD9DV3qzyKeDElIy+
71Dyo1ZAsPu0XE9/j+LnG4NDhh/7RpyyVyHEVWgEt6PN6TqhbKXZUdjYM39JRx8J
pij+seG93CxQ6F+Wjbabw9B6qXHwJRkkLybt/bZL2PFFoEoassp3rmL42lhGW9up
bBvh0bp22FNTLdjzFd84dh1g3Lwm5GvXtg6y4n027XLkUsPn5ek4vUBja3+etgJP
xh6ATB6Yhlgynifn52sOOZxrOczQVfVw4bWsicCc16+3qrCXyn7CgmYq+5szg1TC
haO/X6ehcq31vf61p2wa9KyZrOqdxpjDMgvnUCqC5vDSgPtzfyM2eLdVP232jXN6
5DYE5cJkzL+D3is2yhdZ/sNlsiUoNtgGf58llFhW+BuJU+bwChGDbiMEGGrhdGdZ
BNUqBoE6MpbdoCazJoGkJxLLriRSHh41MqlBwyeoW8WsiYwvT8VLgJK2h43ePkSX
/srJXicPXgdGJAj7YTaVeSRynEDydAI6eQOOf8rdbJSdCPHdnHuxlvo0yg+X1F9t
l24FDqos5U7YQs+P6iWlziUAG8VJH1nyicBvdjgaG/XOfcmUTMqZgHNUVz7ey080
QitG03molHupfWxwjCqzYSaGj120zQjqLJU+jFupGgjbZRQ1RY4uVBeFTgWI8Mby
eI9P+2r1TbPkU1c/dMe0RvGw4ap+x9VGZVhCr0tx14B0p5MEeo277NlU1QmAhBSp
v62ou5ig4Sw1Lz8YgQLaovtFzxO77j2omT5482qH7n9cXAoXHhicKN884lvMF3Sz
Wi7Bdn/lFdwCv4PuYW3t6bcva1vioPj3NuWzovK/gZOMAcoKKoG1hdRK4zFkAIGP
FTPJR5cTQo5AQsXmHCi5KWrOlEHbfTw+h3PdYWJRPSNqbimKKQje3V5VrHUcurlJ
nbbwtdpE4yFDtmPYIB4TiTrBtLyZHsljJ8shmwckDsnhQ2ZKd4HmVYwDBS+4vOpp
2poCjb/0tp9qdcNds3q9hOMCjr9JkuUnrEQ8JwHap/3QwlD3MwWWRt98dWITZobV
H/TO95cRDAv3qDM20Q6qQvHJ2dDI6H5ueTZtY/l6hgV74QezXc5iqSl5SL9eVOrj
8yPXwQVOs97atAxTkfBIHBvzWKZcxDtGHXSTMe3g06AeMLSzaY37mP/kX1mVHS1T
n7TRJG9Wu6v2nvK/Eh3CKidVK6oMtocz+7D85kNU96B5FyA3OhG4mwN/enwiC3eE
mfzxMV436IaMJ4nqCr1WmpE0mnBzeE26nzx0BoisSbKpXIPVKAgyjPAtD1ns8M2g
bbtT6ZkBl1WXbAzQUGXhXjuXN6hK5MAnmi+9+19tUaw8qV2BFFleT8QC0L9gIVaY
RVYV6sfdpX65K/1X8wuwqLGN8LyK18iVsw+aelU9RxnpgZxkGvuHwAKDuGJOgTUi
4nlVSWSpaNnZaGPXb/7ipnp1M9FLSnhPdoRubTQJvveHswHtLJJG7lbeJ93L6wF2
M87JbhxpseM6Tp+LT4kZgUoll7mlLgzbW/zlKZSFyxrU5oftm91T0ApMVMpE9ndm
Eqcz9//F+CL49sLygTkSunUY4CvFDFuj+Dhe+wBUcOrC8pej57YRK2INaRL77obc
lYT6dipPQdXBexmV7PjYjfJVfC0NNAIfe/wm1woMLvSibU1Z5a8CAUdRopzbKYMc
Xx5YfXybBzJLtQ2moFzimFzH5BdrrIu4W31/9Ol98FCEmdYYYChAqUXnMjwO5L+K
uISIKFpeZIBcauaH522W+DHLhaRR8O/4qRUdQg/boQQTAX1DSwCEztkqpowUhaKG
tEImzI2GPQfEOAk0AGis4EdwiL9tRXumXXPXptLgkGcnnKIoZTf+Yl6HqZZRLoqJ
/G630zGuGk8u1ZueCrHHNjpE8RvgnnBfFmrR3Xmg10HiTzSnzUPOMoysgwSPPpR3
Jo1uy/f83dkrIHcOt2N63coZimVJ3nzcl2ZP2/QBewiP7a67HqUiddCHpasEoR/1
/cBQQLeoeG1SqjyOlaw9AnSy5utB/euGIAEGrtBR7l7aIvhuWn+i4uf4SjM/UTih
ebCYFy3aNVlZ6oFdcE+eUyk2/Kxj839mJhrzw6fZZFqNs24ML4VTbRf0zqiGKzvr
fV2MWMQ8IWj89HT2aZ8ysGj8FQ52EMZzF+q8NTT5MElj2xVreeRL/Hfm4JsoYFCb
JEGFaVFqRfFkq0I0HIu8umlXUPn/O50RJT8CMUEv6w4+a92APFEkY6wS4dg/hgBe
t4xxIfCkh6v9soCfD7XqhnPbyr5K76FOQXwlWHwMSMG7mKyRXxUzgn9jpR6ue7i4
TZuyB5j0XF34orw5cHLyOhw6QRa9MF2aEM4BMrcbA0AbDREZDSfJVwo4W0FNtUVi
khm72S3cccgSceMQrAV8WehvyspycQYc1Onvbe3lVnYOOyMY5fXoaiFFh2ObK2G2
zKPolf491tAjEhhSdSMBcny5aRf6Ap6wqEPr1b+IrvcQ+BwLA83aG5Ag6Fm9byPR
fVUrwe5BYTdEHMY8yh/0EMTas35gxRT6mmGRhFwOTwa+P4oPD3B41p1ZxxBQQ3gi
k2N3vUJUOxWT+V6dN7cOG1NS1HA/DXWBstYIZvTLzkf+uTul+wBMd83cFPKQbuNP
mESbFQSJB0c+sFv6Q6ZXZurxt5VpjqUmo5PErGStKCj9cxGPbYPtADV9GECvFnv5
n3IPEFTFiXtcoMyHLKBHkAYXfXCVzG3XDTRF/k8lhz85l8B93uEjW4IntV4jf2ku
JjVjMQBQCBQJc3F/UU1NYvD/7pIPXH7e+xU3g4tGZPpxfEUFDUCqsivCVKxyoLWn
A5NCDVDOYgEzT57nzRAuq7/f2KdQtm1XOAJF9GXuvpeREAbFeDalO3Fc5F9/GKxX
FSAj+LQyXGypK4ydeOeF5WzzKgjEnW50Z1uf4vFs+8p+nf7bF4fuO13LrqmfMVw7
wOy+gLQcLJfqA4ymf7TsYeEozb9ejzcfNOQTk2+2hYPYcVI61CwFVHA0xyfUcBZq
tc6AYEeRsTrQEU2OTK2ip8NU9K4XAS6JXH40xmyz/kmyOxh5uJyrRuNqruTnVzye
T6BnyMxY6e1Fq4PLijuVcdUW/DKFAgzFfXLZUwBhcc/d3OR2XUVtKPw11TAv2cfw
X4/SrmzUp74E4ydRxtBrhQpks1y+UE1J+pp0/IsTg5o7ufImJPEfWfcAHVi+06bD
HRAY8LeZ1ZDf+6gsIEZA2M8G/qFGOCNo5Jp1vqc5jJ3QX2w90NKFwaCCApBv5inN
m/FotlM4CF4t/65DxCEXYFCVaoEZmm955q24T775HQpar7KLzILKwArm9xXV5822
mXj/w++pc9IXBqG3Ox3Bl9vmHVqXtZ18JmPKU+HOC/p7lGKFHK4FY4Hsf8knuFOm
87fnygjWbFFDeqKDefS3SFqq7tCN6B3xdp5oqxGQjnQH1IOAG94XetZyadrPxgOV
7/39z2dkb37C/RwdjyPJJXgPO46hYeljSPRQCc9cjJ++kzGqrxb2zd4T4DK1xtBa
38g/h+cjb/8MDPE7+guZyFwgRJagnyB5MPSQ9P8t8ymJ8yc2r3e62RsTlUS2GLsn
Ik1KZSlCPOXps+ddw7KZw5sF1q6bzfIDnLDZqIEIZv1+x4THv28uIdjNC+U5SM34
RZ5mt1DovchBrkgKF1qjPsAlesOh+rJbcfzRRZERBUQ/YY193hNKmtdop9/FxuRe
nqz9j9j1mJpa2aVpQ49kOVUZpDDTh6R9Yef9jLrzeqFjMcD0LRhypesrY3EOosUi
0o1Hx1zRZYi6fSV5+KIzuyvExG/RO/UKk8k7Ke9yaRaDxt1mzhMjyYQgr0A23KBO
ut9dgOYxEL11KaXi/IlAZfWvmMCBosc9Ped0ioeCUVZCDNSsXTlru1jfpvRpYKsD
uyJmDzjusVb1J5qYbzIYvNWwKNqb3wBgbSe6/efT7GHOzjpl8CIp4moplrAG+NyJ
dovua05xh1o+I8Ev53hzztoDGOjz+YQ8HXPFmITUs7g4vOWgIFJleldbLqyMxqMB
zfnpnvLiqcIZNd5jE0rfobk/hFSy8DYSHdv5jnKTBA37qd8Fmqe+BvE6f5V5YuQB
XEXsPw4trcq+ZcnU+0/9XZekxb44myGiQxQulOnxbqv438Z9kOSjYYT8UbT2qgHI
9z1OFwdj9qGPw3ykRENzV+IX6Hp7Qhv/mbQ2WVbbCFJQmxQH8GLimTA2ncyqnUUD
bm/90TcuHGmSq/QwYL4y8/EQhs3KwPSYgj3fzd53gUGwypWimJgajNJ5lK7VWWuV
Jn+ldevLWwnv77ifNtanG/5ATRQptz2MjBcneSAKJuzJU7pm/wG3SfTa8MT7w1Sp
jBbgc3G6NsSkwpe+tBKqunFXh1Ij4jQPWZ+dagTy9Lb3/4QH6gcX7kKXDIQoAFTG
vfxumhSvPdcIxlIRxcxg8ZTTUVjt5btlHbCLEEMPuS+NihLqAGy89orZ1cTjrJ0M
CbeVwU/AU2UJ3xX0/qeWtaYA7eMi19JlPWkQfBeOECMgdyJdQdIyAdGEi4FW0CZK
q2K5WHw5coYIwwLJJpLM9UxecHeI3oV9cApWZRT7fSMZQbWYnT9x1WRXBOVmwcQo
uwpUnayUtIUPVwbLcTSATXT1hNtRV9TGtRs4QA50qcmUkJ0VV5ukbMXehGyPvxG7
C6GHFJ5b1tZeO71nYS0KrrDIhIzVFLTY6T6fWlvz0CQR5e7LsWqEieW4FKC8b9b7
ad63FSbXEoI+bgblR0jKQLpMLdIIIMA4+vdPcu5NOKEReKxh/XEjABFkWHmRpkUD
fGkXan6Z8YzjdK4QsFm9irjDmo2rnSDut3kJQuT2M3+If0BwOlnvu28+69gByygt
zIeOLRxpDgRL9A7uJprXZ1VygZ8g2JBDPf8LhgtYNi3X0/ma8xbubsJmitftZ4bB
QpYXjk+tAcRlVrTE4I5qMxdnCbl1WvunIkdoUb57JRibZ9SPh9OAIfA0QR8DqzUz
cPvvTNqXr1S2taOAw/3RTJt3NUSGueiUo9Mt5pLciz3QBLMJlYfLjuBIq9trdMnU
jIXJJRO3h1EFDXX6h0CwpiR9nyaS1bawMdTotTGu5soRzYbzlX+adkVfPAuCSS20
+71IRwGHYy/QySRndli7iZkjsmlfSBpg4cOgo4x0yBaxqjCrIHdoKVoI1KY+/AGG
K8aXwVy1t3ENMJ88JwOy7lOPiBTila13L4C8eiF48a66ab7lnvrEgg6HizWUuaNC
UoeFydZaMOVYRlFzkwE/5QE2R/5oEUwdEIQwaeYObJ4Rvt5jqgFJWwYXWvFNfJV7
mfxp+WYGnkrgJhv2OZUDj3r/xVaA1EWDpfOY8J3VtYAfF0l83aCIT+CB5XzINEyS
9g3IGZ5qBLdzdO1kyppv0HcdE6a6dg5024WIwBboBsG8JCCy2EBrj2Nd299U13KA
48NMyWJfWyip9Nj4MX2ybDSLjBZRY9QNWzsbMLB8YHYgMxP4IhFLqTGdx4NMy+qc
c7gqryZr2A+NHoOYomDj29yrlcXFAE2LtQbMFfa56V/1IY7AH89I/l1x98hZ0uZT
/3jwDtsSeMicpMNF3tz9IO5nUjs182tX8InZKvcqSUlVvnB+hj3lM9kjZuhsXuIE
8EGBm0/p0EjRa7j6r+MkeU86Rg+KuaYy6Afuk0bSiXS/N8fyjLYfH6WeX0/9WDLF
vOguCvRDt7LyBl6HwwV1C8bglYt0pkdKE+NQYMO9sfIa8X4ZM1sStAXz3IiYCZN8
063Z89m1KsOVgQVKzATk4V/0eDj9ltA/aSs4LL0qaX+rKGFsaqRXShasZk7xNEa0
1r2ZeeAsGg5sOumct82ZW0wgXddPpvl4HLbvWTHDJQHimCcQtGD/6ejj3qPuaeA5
kqi0t+kYMz/WW/aoDWtIWxyLcEZtQQp/y8XN5iMnyH5PVL5kv6c75yLnYs1EuKa0
KmQxJQTHFON8Jj5efYQa43ohbTCGlA+UOLXSc0Gsc11z1xnOPJ/DC4cGtge8V2aP
IVhQJuoHe61zP691OSy8Oaajv4t/FLwYJifC+caFXIj/D1GSZzw+EJlNS+6mFjJO
mot+o4oY/lFm4Cokc2mkY3+Z0mlIyGiSrrNbOFf3CAfqYbP1jxAC5J9nBT3BGBU/
+TZJ/QdtVEfO1oOh2Zh6+aifcfhSMmaBrUAKjUtG4ybXQQU7KGrQhQcxund356ha
kGGKdI9vWUtTvmMvSD4YzstfNM4L107FZ1UiQ5mdiZBqYGsK4fVMiwv6bu1RRCaw
I/+E+pyuYDQR4b1gjvfZgC1uKB+GZsOLlSGN/wCLIQCOYuCKIHJnHGN2W90T88JJ
qtOdnVNQyX4qpD92JLo3OgbnWww5+BcBsh2lZ1WJpZO4Z9q0/98U7VOKLX8MP3Wi
4XdWTDCzzOuPR/Mdbps/GnEscdbP5bdQcz7AwfjJLGtB39tYtSszFsOxqOZqjCBc
AfpK7uhRL4068IkPk9sFJWKfvgaBw3M4/6kywaYusu2VZ2qmDE71DdlISkDGWHel
ScYuL44L1P58N6AWV2gLF8v3GQBnJ/3FmL1NNG3VG9Rksa2M4jHdP22JDfCqfy/O
PWM4tZbu30mG6milcykVWdBV6/otUDPKElcbyQRVbDSQz0STpkJ0N26afuy37CyS
JBW1zpQbr5LV4AYWJk59o4hkuRFuCBoOfaU5KzToAWs2I9dBHvUYyJifgIq2/wjI
CPb7lj4APU4sYLBkviIXEbgaWwGQqcr7vYt7FesxekC0GXIcZl2Qm4UCrEF+Rt+O
Pw+VxwVGQDLw0awQ5hdt7hbyMIpVlJxsB7Lmjf+YePy0jQ3l3TJloT6iXP1Y9/WU
d9R/im+mOleTbMau+Pr0M50J2uzEUpjE+5NjcHQBCez7B++byog0As3O6RB/JpB3
nY6F1ZXF8uvRChjY8ReZmscn9ItpzdNwqUKEwkNJfZYQahdNmHFh9DxUdqZFhWQc
ILLKugerj7Mb1Y+cR4tbwAgUAwGbgxIvekuTtW1IFUXUc5T1M6rDtfhMZulGwr4l
sH+WV42L0tMzfhfU35c3FnHe/XUhMormEmPHp6mk7uqseYcc6GqU/j+N8OiEFeak
tt7+XyI3508KKVHaMVGZ6Vo/aOYipBCGqen4PGGqWa5Q0n4CM/hPm/RmcKDD28AG
EKhx1ZfO0ZKUFdptfXT5NrTNadJtZSBOUYBpTbNwy/uGQHfp/z+yB2WvZu/zqwVv
rF3JXUMCHaXELBvAlTehjuW1tDJXVY1BEspa8KB9Ch78VKJWSKv7PB6IQ0tHO1Ia
1uRhTOI78sU/98OeORigdzGptykHxZl08Wq6ZUQCZMsV5zqeM5cC60AERs7AKwh5
OREpEXruvjDHAHiESABXXRskrJMF0JYZEmkZP+caR3lgEOKtQjsVC8+dijYOjfMM
+Jtb4Up1Izd8URqvFg4/+29pq65V2mrxAsOkyVwoVje6yauwOve/ssI0Q/CS0qZA
ZfZzXlELuFOsKZjMiGEvPh7CiAIVp+kPE/2yGPQw5Oszj81mw6R+wK8kRdeC7ePj
rLJ+3ewPzUrUzLVwkiJbuYXeWg/p3kEK0oyVY7Ao35qTCZZ/KTCqRYeZZQgfM/yE
CfYR9Qpgq/7+SmNOya64iHVVmNZB5Y7j0B5Zzv5EnKShaNc9aceUvYc0MWfURqis
ayTC1Ujx+sahClI0BMgBsaHSUoliiXAeRCz8yo0+odxd0FxPIbyMWez1wbIUepZ+
YQNYLlBHszsRKYCiHvAZCrSD6fcxYSSSRHyW+45Ixc3k16v3bVW26+Qv87IrXO5Y
cJ92W0/isl48Bu+BybyUBoXiAghJmqazGLqTlTeeCAhpBrNuLl7yvcSoEE/WSrTe
Bl8IiuHdMFGI1T7BW3dZMud7e6ZfMnrQHHELUYbP/2O0Aj8dR4rGN5Z2RBg0scBA
oCUWqORMR87DC+THtn92MDv2AEay7lNFy3SMugc7eACWLzZXQnjHy/TfoY6iSko3
gfqB5PU2XO1+zIqSIc5dbfjZjUxy5RpdU6rJsNzn3c7uYX5XHrFDJ4IhNb2DUh6Y
u0kyM96cg1+8mavPHSUATWk3zdW18qRoOE6kJn01YSG507n5BdzFi5mZvAaDvLFd
qirOwXUtFpoWsbHuz5dU44fGHk0vUPSCHV/lf+NlWt3VeNxjVNUaMkDTT7WRQzCZ
FpS66bpWYLmQtRxY+jmmq2cIvYS4oeU5QcOiVHVBcf5qyaVzF1fkt7V3LK1FlFQv
/s18FM+fSfOgijcNKBHx7KNE5R5y4cQuIGZ3+rXugS2GCCCMRQ25LDqC+bol+QNV
1Wxml5fmzdn8Zjqw7ytPM9usbXhZY7TT/NZEwi5O81R1yaxZX+g+Znm2EOyN2ESy
jN/5pHKXouxs/DkTiM53a8DOSecqPxDxu+XLdowenGdt5FrUvmYyjoOJyuHdpr+y
igGqtidNOzw0v1d3e2NFJDG0FKn/EObX1w27FzQkcS19UBEcRRbNO6KPCkNLNYG+
MYke6b14+49jW696cmZlj8g1JOrc2x6o/WzCMF/06ABJqmgxv+ZPmO3B/SOrLM3M
rymjnJvaO1FeDXJM63HF4+ThyKtqP6uaJ5rBXfH1lJkfzWL9xTCg+JUchfkTpJK4
3woZzh7jY4HwP99dDh+yGklS3xPXhnl/wGZnBjZjrzV8vMkANw80HOXaMxdPK3PX
02xZ9NaHPGVE6s3KuiwuOIMYOVgmiBk4p7eR+6zpMgHYfzbTKneo/N7mJjuVbPAG
xEJDlH/ehFpkAzAJ6LQ+ajBilWhtrdqyAbW5xO1E4js5C6kBFH0B4Gk8XZRSW6I1
aOBkxqqc3J5G2Uu+vFtQLsb7FkO5MxYYIUkyxdAUhskfdg8HyaroOF04zz3BGbKz
z7qoHkNkhH7IuNL1EldAB6l4HdBiFVB/Dxg7+yi0I6qeI3e0xTTFfHjtnQpizBEd
bLJMi1Q96nEix1GYtsa+Q5n/F5FC783fgN3fXh7c3+UqNhLzCXg4siGqskxnVbW7
lx8aZHVSRRgZolvCQAmQHm3VUEqAlF7jr3TMAeuOWR7E+pF/Rt5iLZWd9iSTHtxt
YJOTEjmKnc9yy6Te+iXLikkDVXgJNpaC8xqve/diZPYnpb2Y3BRae/NlxmHFPrKB
RYwyJT7a6cTClzoM4rbyBIEt9eVIhDhW2NOjHFjwKV7p9BCJX2oA7qRpz1U18ray
GfEnwqIOd3YnWGEFKk4X6DPwEPwBbA8ebmPG+uXsYlIeCfBVFsngOIE1OejQoHtw
mwq7QFR9y6SKQhOgnByQQpR/dh/TN8pfFmmRUq+5Ou1eDgYFkA2rSqKMdDp0GczP
`pragma protect end_protected
