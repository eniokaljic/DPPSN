// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ULfv13OyItKl8jXE8luiNd/4t8V947uqOCGkLQJRY+MIm51QyUeyPJq4jBDAEP0f
Og/pOhlGG+43MWmWz52isfFOimBoibH0pgc8YZVgUGl9kWBTrqocRnzM1HcllBMD
OvnA2zH9EWzRTzhfwXDLV4d2MLpct5HtmHppMOywHE8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28800)
tE4Yhvq9Gmj+7War6fZ6qUJDS/2ZeUbFzFDwMr0bE4Rhwi4f2PCCSxffgwi+zlRr
jlyJCP+Kr9LY05S1oesiNAcAUCFV3a7HQcSKu69DqqZ3+YmTcRBMFP55Yn4Vug3T
3siPdKJlFMl5mdRdA9CIRbI63OxztW037vLixPQKenLobn+nZvWQAdEA7P7ZtbR7
YjdfTQSQXiPM6Jhv74rMWh2Yx5dnL9M7FM6Mw7pkkqhEUCcgSOTeB4Oc4eM2nIJk
nX/em5E7gWMJ9qYC9TbCbempykiJGOwsako2JztMYmd+Pu40nd7DI6AGFJucTUBh
bsLeQz+0nCnjPSPBr+fI/5p1FijujA7BXLPxdwnTMH/Tx3KwOfe0dYTiHdhq+6GZ
j9njg+TbeWi3Fna4Rm0HQto+C9eTohdgDMXmW9aOXsuNw3E2QArFA7/iRaFKj9bg
m1SbjgsqqcNzOqtAQtoMzuCY4jp9HVVf2Dz+L4UHnPYWyL2ip5H9G4dENS0FxPG9
clRdwGQMzh3Bg5C8BGU6CltNe40RH1LUsAyYu1k7wi1/Y7LsnH92kgNGGwpkLwM9
3Qb0OdNEyTSKHN3n+0TVmRoyOZKlXW+Jf8iXo6/a3CKkkPnVbF1OFDGGsJ0R87g9
UqUOMOO91AiUOVSM5E7fFijS3BDFTqfLkLd14y6E6SMmlHoIDF4QSXy2pYBVQUEJ
J7jHcYOAW9bjfglc/Ic9xhqnvaTVEJq+OlcOn50HJcfNnyVlM4W4JvRlCUEV74Ez
IG0AYItzKzg42bR0RixM05756/gBIjfFrepFnyStrFPsemy/0QlshhQ9wrf0WZCz
e1jO8emPsz2fjcR0otVlJzeyBpak8oXwZsVGkscFHyALSscxCP62wsCJfOsoyRjs
kG7WCMD9aEwZwYfjUgx2iBCXnZIS7OjmHMPJ/VCQDsgkIEqcOks9aBL6sLn/AfjE
j8X3d48TuvFaX0Z+SXeU0/wwJHciNiTImvshlcV3q2ZgWUoS46c4V7hJmEdxfoHN
4/QA68Y8aaOCXgtrQ4zIoYgxnvkbUontHtnqhgjByIMsas8UUuNBFSM+xzG8oPrb
TVHsrontk00H6Gp4s0tbMQ8kJbSmpJmxcHv2qqjTJ9nKrDSZcPK0mn8XIqKQTJle
zrsh//arwHVZEGsUUE4EYsAAoGftz8QE3p/B9HufMidZdQYCsFWFaZy//WChTahX
3jN8qnSZ5QIfoVVeAEeG+i5NJSMPQEz0wU3EZ9cu59Xh3Ug+apS7KEvEd6faLJqP
UZkeuW/bG2B2qVNak78q7kFtbiLO6Doac72vl6s+O4fBlXMgVg2bt9JmqLlVlL4z
GB1+3bkkVmeUvYPgijlO8B2pVqKBo5qjbb8mXL6L5KM/3o9Oscz0p2Kn9nYPBzb0
G2cXz2iptrDYgZiFhfHm7FidlNGp6v68d8Z+JaBsdpjHLxcs3YjkjX/2C4rFfXza
Ub8/vt5WSSomvEv8gOs16QyRPESZoZyHA0OkA5QTOQEPaBJzeSbPX6uLNAUlWNCm
E7yYLCWsYecCuXzw8fNlRiroEPSR2+KMbjIyrnB0u9wkqRIBaQi7rxwvNwc0i8vK
1R2jASuDFZ83eRcUrvXFGzIOpofv3TWM+5FvApTTj+wjTm3JCq7hRd2k5goEQaXE
s1vVMxMUjMNsDfIcLWLdYgjmK9QBBYjx1IEGIebhGi79Q+UmfTtJdoGcjtZXUVam
pc0QHWPon1TIBvP3G1O2z6R3oS9aQczaaFA1qG9tv/wmzzOiIT4hqosQ+O/VHr+N
WE5oOUhwokJG4icm4lAAwFFBIDBVacVJSq04lzSOYxn1fIT76+chLipx+zarufWR
zQB09z7/EQIlev9M+ySxJ6GJ99whvSBUpRkgk2Q6Qg/iJSCpvC7g2/kGNExDRgMe
yA/zdbRqG9Qq1AqYBW49cu4pbMrZe3ntd5PWZ6L3G3wTPr4hVPBBnTiaAcvkv2HQ
z8E02XQyJTWe9xJ4X2TpRqZ3R3PRSaqVw63e7eK0AtxhalfUh8CiemnciUKFDQOS
Mqjt14/J3cuAFAPxshyhwWf2f8XVe102pw7mqQSgph+a5K3ApR0O9N3q2Gkhafzl
c3c8HAAxIu4SLA4/cNYbHcnIHo+NSFn6yz3DM4wgLhiHthFLxH8YpLK9GfsI3u3U
dPEYOlP36QdJ7x2i+Fa95Ibb5yjJTAhtfC4JayMP1SGnw4K31reaGaemJ13x7XlC
YcSjrLQXkxSTredlWHSVTAvHgNgG0lHeMCIzlGfrk/uNR9QeK6hmLT+D7jGRcrdN
E+g19CSfMTePITv21zz7E6istkIEW5Sg4e6lI934QPDUdUUvOUokpeqCdcqZAALl
0yABccwVuit9aF6MNGXEkWcYFP9EXlv/SYskKgt4VScW+1yqU7/9sVBbNzMOk5Ax
0J9HrvrEahg4XeRdVllni3SoxbR9irYBr0vj0KaMqjLemS9qC7bi4EIQQ2hL20l4
BlzFIiYo2ES5aRgAKS1ko4JylmPpXEsFhhqwDkR1Ox1HDf5+wlwfYSEcSwkAEPjI
4ZMgghrWVad8hrzYqsUuPWRsDMfCWd8m6Q6ZfiUPdXupsSOoVa/AIjjNu2y2xSMw
qUOLFqB88QBN8hxWFgcU4PZNf5TWyOD6NJUFjvesgReZlINq1qS3zK9nbWEFzft2
v002CNP5qwH5yuHse/tpI09JnowiV/mAmjnb2kLGfxXBsJZIMDM93zenVZRrjGKS
pox7/XsVSt553TbhbsfDpN39kmNNmiP7a30uoaP0wsdsS6KZVHlkD6XDScL/31V1
Z0Od8FSehxa/IrCvsNhilymytSuP8B6N82YVDdIZe9aFNo6mHmBM3Z2Yd6R/By6k
d0+QL+F6Kjn2v0jdvF/YrEbUrZhn1Tr1Nc/1kVLirZKSkC32guPa7j/mv7lDkkqx
I8qfEQSFWHAWbQXj5TzbFBzJTxBvjnlJXVn0nG39nxDsWyLeuAmZNBsm3MAjrpSK
kKGN3EUwh3wficH3SIm01xbLZMa5P9sOJy4EtXDPgfrhaa4yUhbNNB/XJ8QBjPNP
5oVK7oSPQ92367As9O+gYFYaIRS4rZ/7PV+ObRlDg0c3bYIjunXqN1utHeObTZhR
FOQZFutkwlqF2svMBSwRLywuQfYFfPsrN2F1SfMTb8Gd6QD1y+JoYAsByQ4q+2TS
gZD8bg3SV0568lQGyANUrG/U3Lu+rxrFCP5T/UY1sHqsbAc3Da4dMWLmxzBSaT9A
m2d1i6MCCEM1+YhHS6Suda2AqlgyyflhILeF1XJEuBbnF/p77yW70tAlWaMmx43X
uNfAALXoi4csCQccYkOosZcdckRlIK2YlfhPct0iQhowS/xZjDFVitQ4RqSVKsAe
nYjQHl/LPZgOHXqrX8r15FydYZKTUWS/dRCH10rnA/ji205JIWQeRt+fose5vL1u
XIZQU78cEZ9oo3UfAPhmEhUi31FBJt38Kz79zy1IzKlhZgAubqSLik4vU5iqByrT
MWfxUpDE2HBhMtr+16uAFpWquKQ206zaQC9mUDLnECap3Jno4ODkart6J6b6uPve
DjWcjxbdU9+wlJ2o4zFwStp2zJiXiuJDNjMx+6QsVJchW3+/l+2KYmGyIIFT17iG
0skURgKlh4ErImCdPs12XMDON1Rede3UZ2UHVDoojsKKG50NDSk6fnu7WbR0bnUi
52164zoiRQreZ/rJGjz/tA1+kq32tUzbRflJZkEqEFKmZZPzv4oSuYCv+qYAs5q8
ntrWbf6Do0W54NM6PH6ILBY8A8leiuwQADbcPCrLNoMbU6KpJ0Xw9CSUDP5s2GhM
a8huTdWd77Iw/x8acWhqKnUv8jRMZx7Qkg4EwIoysY0GKxEVo5+erwb3nEaSqEIc
6Qmyw0STSgauzZYW7uBQ4gUFbvVZFBwT3M0/3cp7oykoVgyE5Ilqb/pfHSKWLVDD
HOp0mohiyCjXeHzDyzhN05OA84oA84pOoxQhTjaVtK1YiHnBPFipMNyFe9RkVOrX
PdMaVnwCrtNoRG/sVeoqaPmfyXaK2ZbcAhKCb2DPR/BGJnxW5Xmu/3zcTE9yyGgG
B/H8zInVBMQG1JM6v4vfuNjqukPGNivAvBW61gQH1/QniELnMclMdHNP4lTZeUbb
yGqCqaJ6IMnyO5jXzKX4YB/59PUSOGqTFtQj5dtBZq1gVAbEwUKk5GlS73mR0XQA
0+etGlOMrkH0GFZ80eX8Ekk8nwxjf/Aki04QAyGCZcr/G/iF624RApvhBkbI9r3L
GvSLdxW/2cUvNexe7gS+tK00j5bf2axsIm+ktH2P5nQBf+ZBM3R/5EfoCiVOgczf
6JrCKI6yH6+L9ZRk+/PQt2Mg2vk0VJVd5JTJXEofAt5jTUExpO275rR9KKoT5mrW
/OF9TXNQ9U76yvIGs5ZJuDmwqq12h+xySnpK4Mb2X97c5cOOCLI98bXbax9dTvFP
NE/N8N0maLDjzozpeAxpaP9pPEf+1wdHKvwtm+BfJHeuta/EBdZ65hgdDVFfJhYA
907ezsMUHRPsZ+JBwomGdwRcybLrCaYD7wa+bvoTKpx9MmP7VPfUk4pBTPKDu9id
ZEhwhxeFOs06OCWKOTSEtMB4M8TFPMjJ1XZn4+B60js1Lwer11Ou6eZSblzFxpV4
zqV9E7JmI4H7eCw1/kagJ+F63KXW3YtwFNzsyv8kV5CyssyPxyg5JzT1NI9almDg
3zv2dLfVU/qwJ0PNrpn+cb4hMkaQqiaE8O6BFSxHsJsg0OySp7rGaXawjkDhFwbA
GJ44ns3g57VHcE/3WheeCo+Z4ZWH/c5SFy++69ziP4nEkWy1x/JovzvvM+ZELXYq
nNP8lROl4SX1t2IO1htj5IUaNLeiwp4gAe4MsVXjPIyJ7Ntc6LX3KNHph8BRY/+1
g1IPXYmDzejhIlhQAToZuoPXtTFgepiRO1hJu6kJT9Npp/XU96vHz44//VAtN1o3
5v0KOBpWFp9c92yKbiSdcJLJevIRvQI21cvwrqRUIsTzQFURbdGjYGQzSIwD2yYJ
ve0w1fWndIq3tUBPK3coEDIAbrRHSj7yQhGPvmuyeNsAbuKPyi8XX+M7/isLryn/
XFucllu6u/xg4m79C/EpjLBpNLpdgjI7hMFtOcWNM98hkZlSmWwxwKTVVxYriSth
QoJShRK3/li5tJ6/4YwXOfl42OJwBh0ICXg2v6IjUPmUXL2NCuhWTrGNtnUvWcfk
v3x/ZH2lNfe/1hzbECTEuB7s4ia9kw5pPPjzOv5IsaUUB83Y8LlTTTndMUXYXq8I
431PYla+VTw/NY1ms6s4vGUYXH8koMVQ//iijpxZb38Sy6XviAsAPKrcwX+8fs+6
65A6Qz8O1chbEzbHxJYp4fYqmee0usbvum/35JvvlfOtW2amUgPQQUHbpt9fKHYK
IaXEvZNQJN5L6DIYTrIK6PZyHbJZ2EEiAEdbv3m9pHZIglTAg7C3nVDB20Auhoew
jtRfmngHCLzACBeoc3Hmn+/BIw9EymOPBPYbBYg4TwNH5uIW7GgtTn76jxVA8zvn
njVEbW3t1eOAyq5CXgqw0dTOg+301kUA+rpcJN2+FgbmsdsG0CQCH7D3mBdd0Y+V
EmjLU/3dwBCvMg7n59bAahkdnM+AmYh3eBdL4PniYSlQlXoTvT0L6rftTenfwLLz
m9unL1o5fpQpYUwkvfH4Y9A9scxlZUiDUeaR9eJS2cCNSgpFHr5zQ6Im8hKJdyM7
CxR3kwnZ9zBBsp41tiuJBlvOeEuJf5uh4k8Pf/xWSfITNJIIiYSPinL8X2hGJcT9
BUdjd8uABoXy6KcxVHlIpYbyp23qeuxVTYIZeq0Cj80a+Uc+rj3v6xMmVDXB8Cvc
L/K063XE+XkPzWApFgHbK17z7a3n18i5kA+uj1vy2eGjaUef+x3AEHH+btPTYfmY
VFoYXDw/aQixQLkE9tcBVlXP42inSmLDFjxni3ENsaUS+qzmKkNzxvzQlqZ68+nB
Bzh13+kaMkaR+j3vNjYNu3/DdLylm5t9Be5C0UVmDGgW59ypSZAMgcdm3gf9JZEJ
kgE+YrIU1e0ULN1r//bt86mGsYsG+IQHN9hHG6JKQm/szP1KmtfRu2Z2009MTvPW
ZPcLm4Hd3ulKsNhFe76JVN1LyyzsU6huzCfdEj3mAa0I7JVrn1btpvgcd/3Wp7Ur
gCRS8lbgNRxg4Mj3ATKVALt+D0dbTnas0THk+XPnw0ulFg6g+J9N47Tbj/HLunX/
zNTmxYbOvnSOFmtkwkMRDh1SjlRDMZNJQKeEZnzY6d5zQfpTKBeqzOgroX20V1nV
ZaamTqXHG8srgAw4xCU6l5LIhb42WkWUOkz7CfrvVbVtACTKGe2b4aQ8wMkOs1UL
Ks6DRvOhkI9wgFJYcl/+tkLY1U3QuW61o0/P6uj8Ox71pEOAt3HSbf/VxAfbmNiA
4tAyX74yY0uAKbydqjRU/9OC686w878aIXhgyG1nbjTeVHpQlHypQmRp9JBcAEB1
EC64yi97j9LbOhSIvSxgeHZqp3CK/zhvyDTuD1CNZBJLg6CuWdyX1sde/T84fqqJ
/HSQBht/E4xMUE34Gt4CQijQNzN8oBTAf0KAqwXMdj14W2kE55u1hKi6Dg6NiYWS
hmMde4JTa4NfhobBJfjSnxRg7mps/LlVpM2DwApIBw3WipKrKuIBWxuM1YIrQ5WX
Kh/a2HoX0Io8KRhUtuUhyzA98IPG0YPaYki9UscBRmna6K8yGPDBOX1UTKnaYVUJ
h5Ry3emvVUjjbcU1eYXhPDccmaC0M1IR3aHEk1PKsLeFRsCrSaIpDMjpooy6yaAb
BlGuvyPKAsK8qDw+xB/aGb0WdkoDS1RpaiAMN57JiWQVH5m5IeIy6ZgvEq5RcxQ7
KzFMc83Kfleg+h9+nNnPaKwuJNrjBN+Ib1qp5iWqVWBlxUBxcGjiKN6/pinOgY6p
Imeq1YJZjGloKLXbDoPnqw24vg02SUB+TLeQ07J9ZtvoKhCdYYpY3YRr9S3tcz8F
Eu566pH8tScSHULDrsRG8VwPrAE930ZBvdNvSD4Rj8e+cRc8S/FJN97+7YAlIX6G
h+AezLzYJLO1XNMm0zVuLfFJLmMuLgDMZbUKkt+JRtpSNpUge1RlsuWYXuv5GOZe
cYa9i2PWtuNfV4jyjvkCqwGyzjlDWJONYxv25VBJVwtJab8KvxbXOOUL8A3dchQs
ZK5JE4fwaGDWdkvecUitMa81b8Ynfy/u3T5wE5Pf+KEAvciPfN9cY9WvuBudK5Mu
3MF2LS71px9oDzsrNU8i4UtB2CUNqXK5toXCY7Hzsl1RE7M6T/qMjCzovoayFHF+
xrTySHSlSQ7I/jtNLBR8IrGTtXi1rXH9MwND1Lk2PwkXIVAwKVWuVRVwuAYg0yD0
Zv7CKX8gkPhY9EQBsvYNxGARgNkDOm8VywR7Y6V4SgT9UUWfAX5b+/aXknWrDV81
jfhs25tRXkcjYczyYi0dT2dFHfKLXab72o6awXEoIIRpa0gwkOK/YxbLJ+fEkIyY
8a6t/g4yVj9dJ4MjLwpxMirrbrYlt968njgy7NXYRV5H3lcg55DUz5wyYswRbxvX
80iX+iPER2At+TuCxI704aRnqJYUwXdOKVzmZhVhmH65sF76YLstBonMu7eW+3Z1
T+zOzdAUejSqH6lnzBrFzNWBZO+MSqBUQ+bfKC9ENiAuNU3XvoaSXGaBa0lDwrYI
keMbPeJAkEyO4uhxlijchi2QDK+80LjdMnBHUr+Zb2iNZCt8qPsQNOQWPPZSjl6f
8KnMePWZd1z6KVPt+bmRY53Flqxii5/PtSJBMJ/js7imqcGILj+aO8x8y0OG5rWH
P6M3vnR1Eiia1Js7YWY1lcwnvMNvqRDMVuC2MriNeuMRVeHRKRw8TO11ATvceBgA
lv7dH3l4oKghLFb3QAkg3UZpNJTT6UP9deRuLQ0qF7j4lIf6ifZhBT7SkXKulMTb
ZqJoZqkOZywTiV26YJ8aMIuFAjLOHCshbEQD9ZwzbThzMBeIjRCqx4npVHuAw9ep
mbE7Algnot4dB7hZKWIyt7IBanf1xawSpI5FmCb84cUAplHKlCfvERzsI1OZw7cZ
+/KOZffKLBG8w3joYVYHCMlrKAwJoJXf+iebah1Dx13IwBneOANiCUn4s9rfejhc
9RtihMPl3WUfQl2BQRGYWVPCwgAuQwUn5ZCMzr7qEdRhmAKrQPr35+qTeuewkiVd
t29YuQBs9S/AhZXUk1LN/71HGaiZafhLBP9yrLgoITW97vNBlFdB0VOM5kf1NraT
M0F0VPZ1AvlA8o7AR1Fy80Y3TSNzYrA32YIPkZit4PJ5ft/Ho1Dzc4VZNgEB/Z7N
FzmLx5IQ6JzN05IUbQJa9De7QLh14s0AXocSdRb7yQfGxKIQw22FZvruNQydkI53
o9FH6fIBZrxf0e3ntjG0jYKfVTV/nDZeG4rpRtdLpCNYag4/h/uZ/jlGkWP16Xu3
Dlwn+ACN4u77wu+1osJ/epUP2MXti0CU9Ph1CXwQ43vOc8iWjTVqUCvDacfOeleX
shbthk27uc7+lUeBJxnFIPB4GjejWBdKeXqXcHO+HFYKjxubJW6uPz9fDfG4H8rB
UTELUeHrNwJnp8nIP5fXR7+KIXACgcDzpTrXL8R+BLojuCTQcu3U1L/tmgbQ3XPc
XDLGYiHmDh3VGXbVCldWkthx7jumHNzsJhCYC/NqBMiauAzMOpZIu7GuvFEZi037
Tupa3Eatxfy9n2ETtSclnA3RtlBSDj2kwbqm4CZib/2KFf+Fnh41pyLZtUy3B9dq
unKE6Aeij3Zt20DaFmbcvh5yuXniKolAWrTA0cYjFmhjQ6nx0Z09eEoDMW3xwud3
6kQ+qwJ1kP6gAApTfzsLrWdw9plyKJFu9NWjTTMWYtCY0i9OLIQWOdWsgKVKIWsH
JSB67S9DXdrlN06Ds+ZgC4A/HnO7xM1QRzBzlqAqKr937OVMXMCqdIXcBEKWxuRT
+KVUDFdk8OWs07lxgaVUwo/aqnFcbYc4EHe2cwi/pQ7J7TzTC2ySF2OBqLyqOTFG
Ye7sXaGmy7QwZdsH3Y+p0Zel7i8KaNZ07focvrQh0CBhP9MZAbCic7jxl4PrH2GI
bhcfeeak2AHwdsQfiHCsQJ5ETpU1Um6GK0XckJQXmhvaxRb43IxYSfJkQoAVGp0I
Tj7T2o/OiqGaPl2V3mcxBKHuNQmbdh5R1b32vzoj6jXYRI0twym4uuwM+spcWR2X
1tVXVb7Bhc1J8oJ48y6zdGBCyF8zgs9QvHtIUhXjr9/WsQtdi6O3Jgt4g2Ipxaof
O2/EPSY8wVn137g5gc0/0nZ0hsWFS3DBK1rubV+oYz0N3qOsLFT+QgV+jfSJreju
g+RFROtB/6ZN9hswnvhRRXAyYae3DHAMEjAkL3SX9IatIlcjpW60NgcmYC3qZiKT
YUDvyN9D57udZtR5XRiAHEKo2nW3uuKcPWg8EeWGSGTQGVqk6mXYQu7BXCBXv4KJ
FxILu1di+aCzxOj42wDcjemOL18kTTCoxggZieD/VlvWHla+Ts7rrLKMVORacvyA
EscB+PG5NNZzxjT2ejC2KXlnKRHD/YBRww7HhwTwMcbTRdwBAnXWZ2OcfYRhrC9T
FXJyN5K8NTnKQw8lZChRhv6r625OFAay+Y1mnj60uUvQ5bYEC6fe8i4V2J7TPmUg
eRTgcdo9GWOdHplHMiHR5hjVONP2rrrcWIaj/+3OmRKQ36gzsU6hehLHjQqtO60O
01w7EMfV8MYEheNThk+BoelaV5hS0hVmQvBDkNi6eymg6AoH165XrljlQ05LPN1Q
Wryx7TLpwF5bQRmGBioJRWeu07YT+B/4BsTBU4VXbEG/M5GS25Gmt/7GZTdt/xAA
0GpiW8sqKvKDHfN4HL3XmtPnPJQFIRF/eCNjhgSWN8Cl2yHGZs/raDVSADzoTi/u
4BzeqD6HAmhQ+3er8vsYF63qG+Vr2v0wB2vnzV0c5/x6x/r3YNmiyzKWAgxA6fSe
+J4gYK+dMdJZc/nEikJOHzj1cl+1wDxJwoMHeqU6O8M79rS3WLNdC7Nr9rXMpjaD
ZviyHs2sHixZLDuqGjhFb2oBXqRrsGy9qQqPqdh7cgnyy3k7t+tOiAUo71/HfQkb
jhbHT5nMl3zAYnjqKammq4wBFVJG1wrnbXPuGGohDlI7fZ345qSfy5d4xDZecOqn
5dwZHZWd6JI3eLwbg/ebpLjYVwQi2BfHYueOjtq4IhOI1urQJ6sP43+ekVpfya1a
VhxX+CPniEwznZyUazI6N4pTSk2/6gfaL5VcgENM9gT4FUNET/rx2EFaPF2c3kGS
IIzzsSH7O7Up9KCXgt1FhNMSx57pCwDmpU2V5Lf4hXmHvEbUj7U1mTmc7iJNG6P/
TRyjkyNtoc5wBH3peg2PQdu/Y9D9YcV8SBikK1FJVLCeVLbaJW3a4kl+lDyZiXsU
GNR71l+8q82mgHlmFw9UGnsilVhKNK67alOQyYnPQk/8x+EI3TDrEewYft6WIfCc
KUsj8lzo7EUs7BPO+RVM6GoqQKCDQMqGKdV10cEEq92wj1t2asT3OpsGkVSzo5H+
OhuT1NQPQcItTAOJ6Ei50gOIglaSgKPCW/rEWu8ZNdVR01QlGj3aqJbQbgEB3IcC
shYYZNBap4jjstWCkkSUz0SU9HNcApbfIxsYkkGNdnoh44s2Bc42xsdg2/3zrAR3
PRIZDyJRWgTF6BHqvtvrMFPEZ15elBSUsCdJV9Qh0aMudaXSvhxU8oTcV1lUre+N
QtSUiZ+6zEW4L1w6Y0iGWL6rIQwB9TMTg+ud/aHbktQyx6XhrQJLTw9T3SwUImxQ
1MmXM6cY/DtSP6c0kvpj1XNsxAjKrHGkniALvPOeU8Chq7qLV6cx1/WKOvsXqYhv
YyiT1x+u806UMDRqT7AcwUciK3oi6EgqZ/3pjXafhk8YEO7pzfAvX4ymdSPLSe1k
xtU7exEyavuzm72hzGf6wkz6Hcp8w/gqR4pqhTBOeX33ZbPHnEFAuw9wPhO+AL/W
o8O8VKobYM69fOKlQHXQs0fsoyEHzKqwc8qr9OmjqgPx7iJ5bFRiygwqKKQ4Pcp5
qHUZeYx7zND5XgZkyRyewLtnik2plLtG7S+oPAF15OEzOlHD0AMCOAN95kkq/xdW
wFpjSUWx74898WbJ9jqgXxC2Qn1ibxF94FMvtLMB9CgMN9XmQnUwxfNM4xhshWSZ
byzgT4sJJnGdsgZboikACdb8mySyXJSP2sJMYQpNP8DsH7bMdJtBu7Jstx1sK3bB
+feNeoa4PcNK7ITlwumyu+b8Xiv46CY6pisrvFv8grBZLTvCoXAWaCnEZkhtalZi
SWyi7X9yGx87ffQ+X4PdxewMEcotd/nUnPbP1Oyyz/6FfcdHXwF2dyuXDkzNz58B
pFryyrojhM4Z8SirvwqiIKnGiYrtXYwo1woDd5u57fgrI47StrtGHa3aGeFzU9h4
bsDlOYlXQEuHR4c/94o60ubT6WT3Q6juXVFhn7WHDkc3EPnBL+ZGz13Ix3IGczlP
nBqHDumxV0f/SUhQHD6y1vOG95SDqp/qHU7DbM/FCNLKdK36M+NQvDcsZ/mpCpUx
e+BT1eT1iO9kXRoQ2g7E1ml0dw8asUMvwAX/F8I6iRxoEf0MM4nN+saUaB/rf6Rz
Dr3Z3aICdGSau1Hcbqg7ycAIQZ3emP8BHe8kRZpmAPoi7OCJPF5LxM55f2yPeIpT
GNX+3m3d9l6AGGc2Ax5Pd4Itp2NZlTppL5cbQfpfXzRR5QjTIPdfrmAg8ef5HUjt
tbQJGI+bmmZZGY3/hbxr7Bw1a3ieZQzN4WYnaEFRcbRdK9MyECxbQOYTemlSa0Q8
SgyIxTfC+yz1LTKVe2SJqxBt8fCETKeLowE98vOTS0bISNJt9gjaaoVIioBUUPl5
4Z1iFJUUkWfte795lBeitsHTjzraO9cVM9kZj56vc8IfTJAwU594uIaFjk0PGL7J
3n7pdwtBWVAAgN7E8hkwqwbPhrsMoB+ztGk2OVui0Aej+uMRyF2Ljry8gRhVdHmU
2mf9OXBFut1sA7oGA0e1jBa816p5xrXebDZ7A2CgGF+qutOel/823enCJB/Gvxo+
fF4SWClE9fnC3N+3ARerX6/dQMDur/oW0bUEvKuwdjLmJW3eIQDnRX/f7KyJTQaR
r4YwDVUh2/kk/b4mRvWfqpmpkHoBpnskveGS+McHd/Y4M3HWQC3NAjHeB4ZTmDVK
ZrwTbYv0NklIzv8cg9QlQyLNZ2Dp9X9SlnKxkNI3hLQW8g7+h5EpMBYELWx7MwW+
tQGSdyh6cH4UvYTCW+d6dWELyzgJKn6OUaztRfu/TfMn9tGugWn2t9y5Z4uENfrJ
JLQh1DMArF8HpR8B2wrwjJ+ee84DpRyLJV+2JzrYxezKAiNf1oB/9ArRy3ussLM3
mf2eyI4/GpLL8W9xJ4KQ3BrfelarXtB7Zpo9FgOTXo/qFgCWPhu6DxQnxyFd59FW
EFUNoeKqd5ZhwyQ7+Sn+euqm3QlsmPmWVQnIWJQfF/T24eUE/2MKcEe1KGb8wYGe
vIth6/50wDhz/v+UochIfrBl+PGE74QC0u7GydiWIAO7eC/a8CKyXVjRO2zs5c14
kH1BEUO/iwZaLp+mcN1I+aS/9KuetmNGo+OvRI1CRY2dycf5fN0gY278xznp1QMz
7kQ8LoMwyfijwOTBFSMjoev+871JCn5YI1OU/j6EKzaE//xQMQyJNoUPIJJmPVVa
BzEwJfb+v2jHWyhdzOj+CeWPefdbDpKlxQ8G8S0Nn43wQsgxzRA5OxhnWvTLiIm3
a4rd1aRhPVzlt87EZZbqADo5us4pi4eA+MnuEqlO2E2mO5YdTLCPzM2aZSRHAS6q
0UeCMaCnjSF+HRpNNa2ykUiBhZVczp+bYQDRci6RHUt8ahtqmQkVK32aoTSJUULd
Xku6nHKkzWpHeWtGJ+MALdfrZIQT8MRR11UTcZlXAZ0KPHJKDLvPZ8CPQgl0wTZQ
fKU7MoDyS4Ke0TXvNt11U4YWktTpJ0X5oHuEoGF0auGK+EdYP+ZZCGnmWG98S984
yt8xZ9Z0t4w0aiXGZoYYBQgMCTXx9owbqGunwgk+dQWbVybrNb3l6ftzoyCcbHyv
ZjTkVNac1X8u4eYXwfYc2L+A7ITBNcsrhillpSn+4i9OmvImPRLTaOmskZdRJy9r
cgP/fMJHRq6S4jUQG21ZCAHD7pqWPTw8NFqiMCXwRSGhMOU4HPg21k4FDNn29QRJ
od16OgMH41OeFP31nANt4GpEDppD4Pvn/YeWO/K/JLqXnbjxHxhODHb5m/mzVflR
0lzTfYwItlZSy3Nn6VqKY2GQA5jZsFYPNqEOlRnUzdkjrlCHL9RCPl2c0HLH7jsf
hZVqdm2yGveBD9xo+uMdkS3GKrEImRnFkb19H2y+mu/M9pzUE+565LYKK8w3NH/9
S/GrtGswSxIMVFzSDW+hJCYyl7qehWbNcNRe8NNvn7JyCTwqvgTyU8u1FtUd4YTc
4YSfsi/ajvSE5ZIAM1uPRLsZGq0qNPWcGaS3y3nLxYSMPIM2BbXzCVEgZcqKkUIE
dHyytquBbKSFbu0uXqkNKcR3hMNgxfnLGrkTLz72fOV+9CQp4i000c9S5oXSGo0s
jpfq6zb+/15tdZcXDGxY+HcwpqI5zmijtDEWrOVEFCYhD7aO57nBL2VUHSgk+sEI
pKNHEjrMT5fFefBsvzVQTxZ11sNsilL0jEQ+etvkz32N0QGj3LUuYb2lOrmkUXQR
PlP67CZqDgWQ+m8OBgz0NkjPzrO9OwXk5y7KRdOSFrc7Qpfkl8BWsAVO0r0osOq2
rAnRlBwWC4ZZy6pP3LOS4Eu9QeJx6dwNNWNiZGgsDBx+0HXch2atfOJ0jZUb1HiL
vlvKL8kVVTiFEKAkO54OFAv5apfCw8GdAJV9n1kvYIetg0qW8ruBzBoYOl2ocZZ+
gucAAYQrEjrHgFPbg4sCmuqf8pzgLqL8mNHELg6TiJjOYp9ey/nxdnnATR8wIyPe
0F1R7WElKoMEwNB+Uusy9lbVcE/RLGf2KGt8uP7mbnna+AoajqnbH47Px8jqU6N+
ITNh6hBlxUrQE3Yai267TPOXnEchk8Wta5QKlY1cnC2pFV6saOcgZjipOHykI6gy
/XWohSsjxqOHbx8y01pkLyUt7stxs5416PuG+xp1gB4/YiJxTfDjP7j36tZgILXd
3vipmrjubrzM/wNPdDZoPYrnOOVflkBLIPe8vY312++ci+sfBZXdqIqpZjdh9UIS
q6FuJyZr9dYb4RgCm9INPeiU/LbxJpm9MJvRYsV8NRI3mSeq80m6hCcXxvZmdX4C
ov3yQdX8BVClvD5zANiwFQ+NbicUu9P7ZznWBKw3qjSI3R+GFeXLuOHQfOKgGwbc
ckgJKiUTB2+imoUYFDqPU/rTxo5wfR4FifdOy6Blbd5twnkaEIcW6dO5eakieaEy
vYYuOIXpb8Qp++CVhFx20G/8vXVhjpZ3gIiAZGK6PDe7p56xF7E6BeDbMRlEeoIV
4M7GdIwvhXCe6gMizuaJ0/+zEJNFv1lrJh2nZd93EbNOQeOK8nO93OeNUSt0x7hW
zeI40HSq/ZHa89f+E0OUGw6v+HIhDg5XiHW9H075HeoWcuPw4fW0PnQtT4lY8sIU
lzLmnsvdGQAkBZ6rv1jgcOTT7MlczIRU1eyIHEcR1lI/AFUZ6CX1VwXInQtw8WCX
xm/ndwKgXIogZCKHH+9BOi/WdU7A0z0AF4EIkc44EVpaQD8aJz8sB58jOAHY6Nfk
qLHFq2/Lk6WfVB/8Imq5joFMGC6dgp8rXmgfLDPusxmmD7zIi5lRrsEznMwBg6Mp
IFSAYVf9ozVkzXRg60ab+iaZLAd1HSf03lE+hfkO4g5lLZOeMCZ2bM3K9tfnRgvc
rehRT3qJojpVd+hoHcPjLLc52OFJmB3+BXVdgw980Eotd0QKVT+zB1gnZsqMC1sF
0UdNiONAYtKKeS1F+nhcf2oDO71vi16NMV3RpO7TDKvBM7bmM/9174zFeDRaOhWj
RcFNXOh9nnxlukrWjbttQCotyaL8ErV0s9JGRA8dZ9qPkwFZVoI0YFshKpcs+/9M
bvOpRPxhSKD0h78dFeHpxOBolyV8yasZ608rV8CxjesIem6hsg5LYwNE6f5iy91t
RIkBroxGyiIy4kPxIUjR4qlxSO7XAaGHCMir7fSLw0/MXNQb8nwdjXHaxLXyZguD
hH4HuvYbO6irRceR0je7EQW03rGrOzQMUHRynkwJ8TkmiRHLT2jQxZbsj7mrUQEz
lS/Eg5RsC47V7vAOFIuF7IbsS55KLng4AF8puX48NfMRC5FMMJ9bZdsl+d9rep9U
8V//+nF40WRu6WrClHmNbSglqLywmN4Mk4rJaHG3mtdXmyyxUnMDLyCaUSFvhMIT
g9qVk5tZzBHekdXxOfKemZTVTkJwtfoY2qnF1gMl0083OWYu56AP7mEDhjLYsOS7
1ixnXZC3i5efUl6/HRcOB14PoiEP0hmKap8sWF5YjqWYDzwOKjZy+TTA65RKblHL
UqybIgPlyCMphqeIPC7cheqwoAMBkj4NV4kp4f9vSz1DOfhrM5hQYvOXYuefyYfn
PaOb8ozVciVL+99ASUhf0xqCBH0tWoKnD2bFPB2mc4QVKymPzI6yS76N2bs6rlcq
Kmy2PR+kRwM6MdHd4HZKq0p5bLB1Xf8BO3IUn/wpQUtXZ4RXlfjG2mp8DyssCMig
ro+om08ufCN2Z4O0SoLbXRtUDOzsqQDaqWsy29Z+tjhstyLq8RVRvnlz7pRh61St
x7Zpfbn9j9O+eg6Ns+fPpKEWC1QOcjQthoRAVC83LSsXKVnq1BPNO9j6whOpo7Yk
X9zvJghF5iLdD8Xk4x5EjB1VklSUx0Q5oejfF95DeRFzoAdOFGrhXHLxoW+g1gDX
SwmnFPQ+92XrOVgBtAhjsBnC2mfl+V1+8EbDfNJvpoqkd7SBRXOC3DfNQhCSQSdC
ZVcAuAo4cIJhcL1nDq/YfCgl82oCvVeZoFitLaRV+l2Nzb2wft/Qv/NTo0SEQ1kc
nFN9+SK4Nht/K3UuczwPf6zR6SLe7mn573HP5uPdmv4pwcEU4vQMsuy3+itaILFS
Odzj6dVT8UmWA15FXQqFqJrAiYdGTQtkzZui+c91QbkR8txdWtxxeckvF0SuXoj1
cjn+7s35aO7YByCCWG409doA34Q2Ls1gDVKMeAFWntAhPFRlWACvacrvqx8quZm9
wApmKIGd7rvZ7p6ZiVMenCBb7Bm6YpjIJBUF8Zq8BZd7EAE3gFs+kl6lqbH86puu
eEPDnAJiB6X/HwIrANbhHhAqTcPJq6Ny3j5KucPYAJJi4Y1VzPFh9QepdCbVDY2P
+NIqBTYjMmmhv0EnXbeg2ntb+30h9KrwGnX4nimwVBRgShe7Ye55nmKWHLzQ58Ts
hoZ8D/pB41+czY8gcE0wZxMHHWTVSAk22p7lpSfYnbBFJxCcb2CHO5afgN+uq57L
v8srQ2HORR73y/K87I6eWpmDw9+3EbfLfEFGUyHZDrUjdV26qvk2yZMnJPRHZTVN
exnIEvC04XMDtmcnGJb8MTvep2lLliDCNDCcnALixQvWKIdeyKzVpP8TynDhFhvY
z3jwm9EzlSScqNibKdWOK6LgDNGRpXzsCE5Xxx2WBWUwmKenEsRO6+y1njChOyKI
4upg41QYMBge3Qnc9QCUlshImnTO+LV5JohwYRa5DrNzy/0GXn8oUNgtZbmC/2TV
xKKKPdfLsh53XU+viH1IMznHOdslVKPM+agSg9Vkh/XnPO4O8HSZ1bcU6W04l815
dNuw8hKGCQ513qYMMWSteEsENzlyEXteQ1FrnxpWKnuu2mjXYsA6J21BP/ooLHCK
kj66HqfNRc5Xx1tkchQBQyn2MK6JroDqeMdR9uVgwOtJ5jUo/O3lhqldeZM4MGXC
1NAB/EMxzgRuC+J8EuDgfvbB46wEWQ82Yjut9KeX/yQgwlnLde18CkXVYLOU7e+a
wMFK2dFvsxFcE8sil56hhTQ+kkCm01s5FvPUg2n8r8LfWh5r7bVu4JdBeGPFDzW2
6CoD4ms/K7mSitW4C/s9AmCkOYUErZAEjYEKBVfnfMhFGbyABux2gjUhcezfGObJ
HP0Onh2SCt9HdyRxKPGjdsafLk2aO9TeqOaf3vJ5zPidT/BMLk+ywyxqiXMwHOFv
LivyEzpPEohNMNFOsvsRlfUwOa4DGSVumE0UF/CllNndUjwj1RngXV8vL+Klgby5
IdfQcDZJ91DL/kzRAujrMh6FsNjOXUdhTemWFI6vC0znugOyomcamoCPPUQm7fmF
hymGID1UxTnbqTRENe6+Z/h5V9H4ifh7HkC72uTgmxHBdPE/ydlgss2PlQ4UBNHg
4LMM5WWQXbu+VK6clovYl8HnivJwYkDcVon1Ns+gikOwfQ5GsGBYYVLOJnJice7n
TxmKX661gqV3KMcduWWc+bgWBPcY61cCkH+oI/lWOnrmzGnC/wJ3ywXRu68N83xA
v5V+JcGPoN5DU1gbTSeZEu5Mg+iijtPUzerua04yqceT8IshvGe6cEy/yGWzcjCX
4dlPv1+rvBZAor8RcI3TSP0E9HHE/EvGER3PQkEPoVc+0QlxWzUdABINpB00kj+1
zueez043EDmHVJZg6zwbIcHz2CT9UHKISeCJ45UzTKw75XaYrc1s2ZdXQ7lBmoid
n7e8FL7etesLtkREXX2wKrF8IUXpLSNRi+ZmlKm40Bu2QY868711Tu+ZVyHqW9uf
ZlJy/HppOWae1YECgtlYegcuoJxNjY/iysm8GTxuHMjQRA9ovy5T9uWt4Nepk5nj
ayZJUmeagwOcHQR3p3b8JlIiSrxc3jUa1U+KjVddVLDcRbiOT7cvC/Kb3/jP8X80
wgS3kziYFybQOebfzLO+LB9wSmwMKx6J+dlxp/X/3huL2hFdnChX0vC4SMHDd6hc
odN8/HqHiDo+3ufiD/J6mlSgQ7Yf1Ql2p/3YUDG8OIaOTiXsH+Xv8s0y6cgkMXKR
Pi+FuIoguyNnGS9BHc3re+sAG6/0ag3C8OM9w15XLN5WA1+0y4MEz+Y+480AfM4h
TG592elaT1cjLusSnVDQKwMeN9KPlgvXf261ZYPco46qkOUXNfAn3O/k0joHo50N
H+dQfcBr0ugIyQgTQQ8Jsit3pmQNWlXSfEKR2yz0/bXif8PwzBnb+p6N0WVdAVSe
4DSzVl98FgbAhU9qaE4M4O4AwkgfT90GBhlexfTAfEreRunFtB0VEVPD3sMpNwKk
os/FJNEXhixOMkFX1gahIhqoRliRK5EVoRn5UXMCKPCefbYj9CaVYsmCJ78/FrrP
m+O2J0JFPFQt2vWMCnvtp3Woin3z3OrVfkVUVDdC5fdzrUyp32ubp4mlp339KO/6
ziUusGzZt6fal8+4j+RqKSZkk8wrXESL8hKj17jhITpCaNUbpRxxeNKjOddThIWJ
VVvcRHAfP5PyVDCDkwkgkxebJDhCl+CfJjc1cJx7clebSwTnhAT1FCTmmyVbCGIj
jHnSlsXtGvU7EANaCgolV1bcmO5A0Puq//hKRo1n35lm8qPDzSOaEZzhkRe2yrrY
8G3PUnv/BaAReTPao9n4CQ+zpFGIxPt3pAzbBu7xoAw/aGO5Kh+Di121pZ6hSbmL
dHPwUcZ23Dy+e1y2hIVFYPXCDDVJIqZ7Gjcv0xC0dhhSgl/67+mkM3sSZU4yXKrG
N7Q68Nn/aU8kOuFYgfA1CsmDPYyKIf8Mqlt7Es35MRwfkUiVEpIUSSITyFqagUgc
qIekLnI5Ay6+iuLNm5Cwz9mqzz4ytMlcbfc42l3u8bRgeZAiro7X0UMVeEPOvrDu
Y9Wi34JuxqGQPnnE+49x1VkOBaR5sbx0a8cju43ErCyaLks9oF3270gk1sT+Gr2y
prBLsQP1G78IW9Ud17RlmP+A0MNzAcbMt9WJxBRjx+eaUFJaU9a2pX+uQerdUH1S
2pWrRKnquO5f98fHnCFrhZTkahrP+VHwoeyeLlNdGKnz7rPL1WSLZMEtrl4XWh+9
S1jKHsALSCXyGnOMr2EyXBJXpAQvOv2HbH2OGQWzrrI/4twNDoEVwFB8hE0z2Bko
OezxJnCRshtqraL+QmmIRmefk87647/olUca35miGz8RdMuUsT52EXk95EtTCJyP
Fphwy784Xqj4VCDXIAneDzlaxAdJsLu0vMivdKaHfXuZwis5vNpVDqcdfV3Yatwu
vw2xOOu9mtPEZ3Qp3+26ENOg+92YShJ9WFiph4cWBDea3UxVDs8ynCj2aqw0suyy
5bUB1+jvkZ83JqQimjdFBy42Up3WSOuFgaTs4FXM1mtVZWA6JlJq6Cf14rBIOU79
6YS7yDvfUnie9sEl7bb2sr7XolkrUJ/jTwcg+ThLtmMvde9insvRh4uSJYJdU3Kt
iKjnSlLC9nD9G+sGqlr0freOf2UaGCbbhOOZ2ur3ZiLYiRAr7Fcn5jP7HgSIVAYK
gpNuwsEbpWdFpv9aflo2EDLZ30y18JeKjzXTGAg7K9FkW9QLcRBL95pldCaNqoyk
YbVTwtoJ1IxrmQdwqsxBPWm7vTDJ2BUOizzj+ULhlTRAKFJJ692QNAJOIMuUFWuB
/DpBBvAz84Q1pggkWwECjjR7ws4Z0CSnLvavE4obhmd4Evz92mRLG+a6V9q/WdLa
VbXS9+Mn3McF7LuC4tHBlcOC/m5I/9j8OmBzle0y5cIogP6luDSTNMbiU7jZhgBm
s8y9BSsrWCH6jnrF0+c9/jGA1RldfESyZODjOJv85F4OHGRZyuLdGRJ1AV5d6FQN
FNjK1UPlgFBuESxP7OGsAExngGZT0Ay5tqBzVcnGQy+0CAh/sTsKKqXn0H1fj6Wo
Tdxz85Rdd7iVOAdcsZmx5SiuwXRwfWAfOEPhGZxxIdi7vMGJpI0Pf1VedKJud3YV
1xa6rbG3onyDxBfvEFpXic89db8tIjCuTtlaqj36kbVm2MPyvxAmPntHYZPmRJac
5e9sU1YjZ+osC24ir8q7DuUFoW1lEP6EMhPkqRSv/wtUhYZMY66j9XsTh5TdtTMn
tSrfbt1unkbbgvild4hcsd5mRohg6fqdn5kfm3A32IQKGhCxpAwIr3TZp8Y/fb5n
PmDRP67Ugfqh61+3Ruk3ai7DBRCKq0DPqn4VyfvNRf4wEzZapbqMXmM8EHEcMAPd
Wk40WVm1BvuWNrIHTerwN/3MiSQ5jMUuoYOENNW9MPT+pIB1SGfAmP3xApbtd68H
+q5UhYtCE7UWTcpdtFEN5AtMezAweWIABfuqF7ZHADJFOf3Yp20/SQrd6Qxfr604
KU3Kl3JbhN6cWyul7pyABc1FOEBHnenf9B5kCGO75LHUPh8ORu3ruYi8x8zur4AH
SsxH/hDB4AFIXrPOuBzrDyuin3yFWUthcLPoPxg5V5qvctjVCtQD1uCutXX/Jys1
WtsFOLw8EQ/e2iMyiL28O4CZPfx6ou6vUgwHiOfq36Z/0bjOePJDE/ktW9cU9nkD
EhFRBCRKtGxEerPqD+pxQb3XVDPtLBuiTpKl9U+bSef/dUYEHMu0LpA7WoDVK+Ts
KsIu+pij9DjeGiqOdoqMEQ4A3itQ5c+emL4NBevrZY1VyUHTkvlp2T1vZEtfyuFL
8LdGYq3S4hiyglkrn+1wf0oG7kdrnh55uVZXO9WHFHJy/Q8cPyy7mYqiNQHtwJXX
NNao3FauXUh8L1SXR8Y0RjCiyseZ2Dqz7SLhXFzb3yH5hP00TjkMKLt6oY/qBQFq
XL9tZTVBjixOj+0j+QYE1aBjpCtSBfI28AnyntQuQXbnDXFAqWgMc1Hu5RBnXZuX
f2mxnMnqDwCywC3R/c/f+XUVZpceQCkQvQ+CdrnEkvjOncb1qLkMhlV+C/OzO6KA
IYuI2V2P/X5HBbmKECZG32uG5Ff+7NhKYzuVrXkt13aWJy+RSzXd3WBfgX/Q5+La
PnGY4h4Z5jNwsLm8Haz2EzxbB+XJLsNVWDY3ygvt68Y3NTj58zYLiH8ChJjhsotT
bVysaQVDc6SpLc84M+4FmiJMA3xlKmffNj9BEMtVZZ5kLZheeNNVABsCFnaLenW5
wpCkbcAzfvycx71P2TTlyyGM10HocaU9y/idAbcN/Y0QNsncGpnlLEdS/qM6mQt4
YkGfs9YSiSGx53JlA3eG2usL1a1/lN9VsSU1c2e8Baal+cU3BGHvaiOyi6fPgSUT
urZO2iohTPQnA7t6zZQYBj65wYYlrna+P31QxmsGc0BnRoHGRJBhxXNVq4Ox3v2L
CgLYR1eeprWCPV8NKZ21NIx/sfyWQHQ6NObcacUP7H7Rzv4JjlmqP4X3OdzOzimj
Kdaza9mISLj/VAXhFLwjDMnAsr2RJSVGJIEiYUHKYIdseorSJ+o2mDd3zpQdc+k9
Uk+f2SywgDErMnHyJbGv+nhoDGyka9A7465EJt6i9eTMU9JoHpqht07EE2z/aUhG
MUf69Q/hbu/zFN8VsbW1pTujRxny5+bO8rgH0fzZ+bMerEhLxI8bJETYi9KPHp7M
h2DxTGyR2EW0Cg6xV3gIo1peCOQJNdB+Maw8DDLFtGFzrv+bdUpZQqf+l8ifEJqk
PgDzUcrJbOe3cH/wXJgxpX5dpH2ri8RX59fWVB5gPPFAGOxigUjgxM3KdkXAobqm
xXskG/H33YacOTmqTD1+6Wah4/BGVc3mhO3vQHaC7E925Zle7QS8juMi6rvr8p5M
KxXqfNd6fQ8rhuli+K4PiMLaemPs+eKYMAS1HRZdR5DDr60IhFQt/Z3VM5BtbCPY
nP/PM32azM/7Uzhug97XJs1xRAswcEc9h2qzPzK3/oDRwRs+V/uYx0VBOpwGlgvi
mn3Su71aiGMPLfHI3C10xa6V1LovkwPQ2ksDFJTonjjyInB4pqIH7e2JqnFsRdrr
4dx7pSPHgWoI2fvKAFb3Q+Yp0JwFiH3kuSNn9ayb2VG+ZtInp59qhpOqkLFCqBhr
2GlyVTYpMHOUifuSlg3pvg0MmUKYWeM6JU8xWeRM03E/C/t/v/qELb4AuhYr4DMI
b5cFYmIOkQ1rui57ryMLzHbK7MkkmzkK2lYPc+K8rtCvO2eOTlkPjJMjqdOIyYYI
KsuWemx7PLSFhnDaTr9wAWxm1ExKJKHqw3diKc7wzFOXCRZV1fl64tt/sUxVkTNf
m2F0AnFS//AzIXLHIb7JNLnhac6AYHzbLTPMEVqey/T1GdyuXCXzKttethcPxiuL
8riLsaezEpGBNTs0EqvMFFgeqdvCxTkHwa5HDNhGFyqTPFEBafY30SbSKdkAfDFd
cFoqBKsWSbbuvO9pK9CVPokBLl+IijgcCQdVE4XpFo8Tdflmo0nkqp8Q97JyIfEk
dvVoVDjnRU3MwB2qZRiHFb6R97p4IiPntbp05HbJ3YXu4It8V7PugCgaQ82XpCK0
lxSPC9GsqlCrY5Hded7DrIRhYUb5hbXmvbV1oZYU7f2aZBQV92U36nSYr3YPMfAY
2oGTWXJMchY1piILAVD+hg6IgqFDgIkZD++IU+zcccGbASy30iDm3vRpk2cSjsxh
tJCjpzAiqbaHcpnieVamG4Qf3mzHmzeHEmpuPIDieolAVNZv5Jgub+zjp7oZPXTh
AaklfSBYaIkHEB4Jr1oNap4A2Nt22qOkcqfrTBMfKzgvxVmKMi2Yuk+SDJWj2yUL
kKMil8etXyNe9OPkAiVYbtaojqcPAkOGcrITLjDiNPdWVOXA4RcDHN+hXMvSrM6W
6jInvAQ4HBaM54uOuFK7b2JtKE3XuBoqtfWLYGWV+D6Mu8yAx3KoMHBr1i+Vmndc
JiIAPDDVlHg1lo0jenLSPatBKOaRfMCs0D9XpDBXlUOkdB+lDx/uW3PH531tM3B6
mtSOx8xIW3I6gcdO4/j7W42OcwZ2QdOtBIMRtpEKbhxz4uA8rgs5zdvUHVCKHD02
AN6B8QEBcA3Rh+L7cGoeMb6VhQAVPLZXjz865prIhUH9633AzZASv+BDEU4Y3SDH
AE0WAJhMtJh4EKoPTquhxVTPzLl6MTHxyG4r0+cyrXehG/0QTNj89wcl9Wc4sqQB
A9CWU0bqg90jHKxdn/XiP9TAKWRc2TR+F6uePxTAaVmweI235InaKhWWHCuHT2a8
u5YGY1Yks9z7DKnfvHLDJrPpsNarV5nIrpVCoIxBjgV68t8YA4spF6MZGByuZbp0
mXISh5nb2DUOrpQBorjHEbv4zxeMSQfB2FC2fhzWAKQn/sg/L8KE9Vvn6IUD7HIs
rD2TB0gyF2kICs0H7x4yqs3re4xK9gpVnpAFRQwQAhgKi7SfLP0Kv2ApaJxHXcpf
noOR1CIYCiUmKDAMKMZylL3QAZ737L1WekfaC7Z4J3BI99keIEKvV2mnXTrAHi5C
dHUjzhReyn5zf1XzAe/Gwnv5U/Yu+6nGMJ08EVVgBq2aFNm4nFy0x9h0Eigsr3GQ
jGKzwQnhzFFZuXWB50ybaqtgXuJiu7jWGIun4q6EeSyBAJLbB/mHSD3ZpwGkTHAF
jlV497oQ8NlP170sTEXB9+6qNgV6wzSyktgQmjPfbwTK8BbSS43I2fDhQ3b/b8dp
ZEQ2yjNNyda95HyWcQONwkHT6Exym48xOJfVHOWkoLon+jv6HYvFHy7coWmCLERY
NACGEw3leg4tsdgvkPRBwYc/lljrdDdQo27k3rh44jzvDsoaFjA51p7FhX2iIHIi
5cAHwO+faTGnaAxnOXc5eSZn3yp3YVBqXtMcd74gFi9g5QtZU492P/GajxfuQOFv
3OV2sSi6nsUUoPbyglI3b3AFS1ZaCugRch49HUvk043S1O0yfCOBP9kjyfUo1Xp6
3YJNTvYw+oZRkj78kvrrjjdhMikfsVm1dtqK3pXDaNYp/QrA/xZTcJIUIMh5XibB
SbhbpJobYPO3Z78LEW4degjTw4lU3F9rj+6f64Lp4iqrO9NoARBTBUbI4tmeaSG7
jFb+ftnUfj0AcAXmCK7M6mfJOb9MGu2Rf4TBbsyhHbh3UIKwRh+EOse+8Xf5xKnF
V6R+8I5VT4s8Qju+/9lV8OOf4YiThlxZpqgXmoq6e/HCYOW2SLsbLzRQTYuvoJHD
UQh1j841Nrhg5PNlwEen1Q0NYMazK7aIRKqOCWcupiHQRtjrHytQiFUDfFfP+Gum
FA0gmSOGF62BohnXuKF/MYbBLrbujcbeGxLiuYMTHbwPjsTnGqLC9pKWf1txd2Pn
+lJEbdYCrAvile4s9iv7pPdvT/K78rEQVEllnn6jeg2UXXO7UNIHE9lUefGafi+e
QjLaGWTlamEHGbKVJzz/tGhiFGaemq+yuh9IS5FESanipZeJbPAEMyZbFU8q/vlD
J2TmfYg37klJyP5KHmA6buVQXdsKAlZhk8LGjJKzqNOiekMQV4gVRWOJw5XHIj2G
v2xbOaxJ1NbFwUprgcPIEC2EiWAgMaIOTL7xn17J6QltAk2Ag9HZosN3aOVcvPtO
oSVKn1zmZmGLikGwtVwKBer/iDqN0VehRgytkciBH7sQ4MWifHtiDSQ0/96jtxoY
JhqNaLK+0plJm4UdXjN3F1tjqn4Ms0VjMWEw9iNAIDr+5GJSutxPMGYPS4qJZRM4
xo55sJIG/fl6vS4dAq2Ubfoi4VHxUUQy2DWG2CH/4tPtgTpJVD+FH1dikrtplqyO
sahxy+QS+aK4uLDKgnodAkD8sJNetIXC5//b3rFuXN6iiky+1PNGlvHmEkAF/jZ1
Fj7oU8G5ZZYe5gKaQR78Pr2g6XRMMk5PN9petiGCht5ADQRtEq7JSCfuDCz4H77b
Ad4QYAedSJFyaHVeHqTQBgl5ydP//IclvqWdfjHSPEdtZu8TWap+celIx7Qgwqg5
Wph5/EBPnDPgNfQdFW2JroASRx3ul4nNaht/Kkp+87iWgn6AsBg2ex4ZEcBonrEz
baDSG1hyHFULP+xXuBUr01M21IWBUxb84dR/sPLlvbTf53BfU1hPqEa27sDnDaEd
kZRX3JByQgiuyb/ZTurNPBf10RkRTu5hTrAGiSASy+U2LRvOlMHrYjA5ToEAR1b1
kJDFHPgonXVOWKbAkm5rdbOVc9S9h+TsIQitrDE7AiRYkakEvgBGYP/6yD7waM7a
sbcHAivufW2qIjyfSioCstg1b48KIauAdBcRfNEwF/Z8BghnVcY/PaDoKMpWJ5Rc
kkJK4Jq5SK+syyKA+HHoNrGAs4d1WAKSDYPe6MHh4t6k0tejUksB+lr9hdRrFnZy
sA1L0MM+MfzHSYjw8kz5W/GGyLRmmsy30O3CJtocUhWr96JvYDPDYnKwfa8F0Y9b
oRmHB77rnueOfiQSNH9ppnMstjL9UotWwADLjE4dANaLmSiivIBTOdvfF3IhSAGt
RmoMWWKJ94g72D81EbgMrwCQw/FHRcbANo4NhfqM7lIVVocaKcRqGzlVZ8c4rdnt
OtW3RXmu8V/5wD4lzKl5pv2OsHPi63b11HARuSiBP1CNQ7hbByOpUaKaoFpklxoL
wSnBPQryTCni5Yodt6MVQGxq8y3gdcOpVnt3xJU+R+FGaGOhbXDbD0TbDHQkZUmk
/X1gEdLCDqLikHgWpR/pjcvEd4BlnHIxPQ8oY20Int/3f0umGruGX2ztRM0qtN2p
Li37E86mGaEKlvkzKp3yABBl/2naJASL8FSyVsSIQ4pG7Ou+StDmEuLWzKXRbeDj
F9PHXOE6dTmaiuWmpU0A/Qgmd6Cqqp5yKq08mCrlV3oprHxXb2P06MO8jEamgkQo
7im2Oy9PsSE5njt813jI5v/BFaqETNFds7cOFs/sxhBlAWht3cjaefvnElC0Hhf3
BrE8plI4FdfiFZq1QryEznm/mz9/d5zYNHep4T77ggA2eSpFYMsKv7WxrwOz4uyy
D9mVvW4UtksRhyqCZOArZO8WBjqnVgqF5KqfAJEG02440Yn935+y1WohFc1rxpKT
K4pBC3zCWLV4LU+BVfDTXe9//dJPeTrA/YCA2r4OyEO6rTjqG+5NgrcPz0otcMbI
dBjj5doejGjxozIgcnhMFzbqmalCBGQrH1t4JdopqwOWU/ZEWgCescEiYjZhS1ZG
qV97yOUGMca2QF3hiUPM1kuGjzCUW1UtXdcSpsGUqEj7Pnq5xpGYQiU3CSGjrtAM
FlYGh0W7QCT2wh5Os96j3ErERsi16aMVQfsoKoYpVYHTKN5vshjuXNJxMfWrWZr7
GTqYsT0wig+C7308bXQtC4QFFsMN8fHdERnJ+JyqhzU6CzweGMoM2Ze2CqHssa8s
yJiAPOfRbNthGDfnuIO5K3K4BTR+DV8PRLUNZwyTsH8XlsrgGZxv3DF7Iqb0AdgP
k34ebDX9Kx422F7uGjlcNSHN68qfEivOrEA2EHBEdRg04fgLte5rwXH3meIjpXGR
ppi4+dRr94FeiCHeT8aaF3nDBryBgGlpXBwq2gPIGiGQCLUxKxPb4w9uHA7sJMd+
3UUw6wz4n3tA2Gytc0jMO5NGoDWC+cuW2jdeDZN/ZfOuMoGDa42Irc7JYiCJkjMu
Pz1kZ9byBpKd1wy+9eM0WMTwliYBV1a2lt3CSeGzu0pccorKRvmMqjZr/ynYG6EV
eD7rrJmNIO4xivX8KmvFopgfMMHT/8mXjOdnuttdWCPEnsM9l9NnVDq5CjGmwi/Y
GBa8WzcUAg2mmOJVAti66+AjEzS1sKADyYr77aj4hXVWh5+FiSVRkSR92zE4jRTe
lu67o8plEyZuUZUgxNvQ/lMmgRZ4hkVd7jmCkxq7Iifbj4prtBR8pJzLVPLGomXz
H0wQYEh8XLJ3Q6F6XSqBYEUnJcXdoTmxYPadfYBYjuXSDbM6OmWU/pkT7bDERVrr
Jaad0RoU3g2nsxcJzt1vvP9JbqrXY9fCQP/8tc7rNeJbKqrLiQptqfBM7/5xHXPE
59Y+iy4VkzVBtm2RTgfmGyIN5Pui+cVr+dhmTqsWIugdSJsKyTRsAGJMrgSbCQGh
/awdhlBa+QE4CnHKUHva4+fuKe44rLNGcoL0qNWv1NLn4Xx3eHYN/kA1zNP38Uxv
aVl4EE1eLST+yWvpt3G7Ux+/naTBwLQRXVlGoKFe8BQDUlnk2YwOAHQKJLu2170j
Ms7WyE5ntlydT2+jiHfNjGyoUJ5qxVgHerfdBzNw959RWUbUyNpjkBp+iy6oNzZA
aAqyOOFaN2L08NwnbXANl/60+S1atG9Vui3gYlikK5JtO0Wtvdr0OMvRx13Ve7zy
yItr2LnHmD0BFJ7D9xLWsL18xyfSojaNaf/tCf3Y0iDpzQ2Q+KMXxhvSjJy8PEgf
Y0HoeH6/6sZPYjrOchrc7DhdZVZxBZAzymqT278FsoG0zTftXLqa7nSG2trhp4cj
q3sHNSSOhcYF3yXVp4g9j6IMnqI2gkXlrSUY5ruNbzTFcMEBZhG0mhN01FzHorAV
05e7LHU/EZ725Go1BufAsAmDlABzgq0ZoJd7xpkDiVqCnEP1Alc7Jbny0BgFhezV
2O+OGlpMEg+4wJEIXxt34NQCrBxjyJ9IV5qnQ/c6RnAmQt22S0jJNBx7oJnB4qgN
4HA9Rn1Bnq2pmuKDgJpqMYiQ9HB6UHRDBWLKdY4UOApGcWGEkT+4AtyL5h8OdDez
c5XoHcj0UgEMUIiYK2vPRqdWYMUi0aZ7UF9HBY348ZBko+bjMhiWCSsmSUxM8MQ9
4+2TINACHMkE0BgFoBpp0Ypp/cIK8VX3oaIzNyH0bttF0u9wlqYpdFI4BUhiVc71
mchJTrgcRG0Er5Q72LMhm/jnwkFRBr51I1C5yNDG7QsFlyYPM43FVUyoQYQRB8Br
3iblioGj2UMbe3hsXFKopR0iNMuLWCerMZZO3XYIb5icRB7X4y+6VmHySuk13zMo
ZAEbZ749rl6gStxo7iuIeG5FUKo7RwyBYyRBK2DvsXBFMwCxrebqdo0RqYNTNun/
TKIirn2MtDu+fgZeJM/te9WC+AiZxiAZn2aYgoZ5irzLwMVIs+0xF9WUc4LOTBtL
+KyYBBmisMW+MVDzipEv+8/CYlME7Y5SWC8kakjzyA9HPut6Ai230dgjWqUmq1bD
74WeX44JraI3SZyS0NoZpGFzOsW9o1NOhgZACrOWx4GGWFbQOwLav5g5BaaOmfB0
eIfMcLR3xB4mLBxoN5T2axrZr62JUTQpTXpYwYVF2X/noKN8qmRW98Mt5SRgjhcQ
gOYBNvqUa1R46xAc83dRVr8duO3X/CanUeNPPUnUxrFERKzH7Mady3wh1DK0oTYm
HRvz8a4PTEKeQsyzUeZoiam0OpjboZ4YHasSFkpxquwK0X8yRj1WeAewkxgKRUpj
h8mQclQEv/akzOMUz1s4KPvn+FKw+a/X+4of4/Benbo5Dmd6S2GxT87uy64rkQOx
JJooyJggJ0qNCjyuXvq1a6voGwOvbfQdPZ3cp7IS5CnBU5/HgyaKjUZTfOUlCO+B
lVaKAE7+9ksuKbo41W/St84iyZsq7cwo/Lzn8RQVLT8XJvgM3R1eId/Z/zYSjVM4
mMDp0FR/eNGd7+qeJlRaA1IxTZqvgv8NBMpTsOuIi7sYZgWF8fH64bI8BSRhDcGD
8LI72n4BgstCXjA/RVMMxG8qArNHwXKe1Z8BR1ciSIivtmTv00KG+fkroTqCzRtc
pboFXo4eK81ZMXxqkGnvMGppwsSAOJW8vU7Alj4Jih+ZM6K51Et6QTzKgJfr/F6i
tMgC8VcoNrRBchwP36/5PVMI0BJMvsRDyrvs5CX8xPTrFlFKZ4QsKaxM2zL/2iga
9jOtPoAd+OsuO8l6ID7AMpDQREhHIH2NwJB1WP0XjZBaBgTbACax0Q59AibpvavO
i6k5+djjnyB82+sWk2ZzdBM4zyNt3DacBnxmJrVfQdCbG2vRTgeRM/inqsNEbZxw
Z83GYKrnU4izGvbRkIZgGx6/ylRCsDTLV3gk/An0y4IkO+BjoyGFoiJ2wY4TWsaK
/nQ57pA4KB5CD/byukdpDcCv6c37FrSZextdqz8EY+qHq1wJVoXUzPqwDHW0G4Nv
g/oujFDn04nAFq+f95RBjBobA2BJXAMroTMp8TK0gtI033m4nuf6GMu6KtyscgtG
TiyQB3LlXH/vrahAb/9dsjQFTCgdNMXzduO9oLPWZi7xiebl9biPoAfFTju4+wwq
5qjgMhnMOrrrqCdBTfCkKpUlShitvimQK1sbMhrxvVCwdStPQFyPXnZsPEGHcltm
xyHLk6gC2/Zvbe/aX94SGLjVl3KtK8HkickLL4JLegEZKca5BWvm1YHbJx57oDIJ
quc1bRUIU1kBtVDA69zGsXgqeRivTVasoc0lbjIco82Upw9EU7CjuRmruKSueIoL
1LqCRsM7nljWq+r+wgtDkUP2EMcIziM9XH2jREy1HJa3wDLJVqhINE5tnqJl66o0
vnWn7VObtgGnsge76ia6U+MhNG31E96SRkwN+aFpU5mqw5lfkeBYvKSmf72zOb54
vBpUEeNI+EqBBHe0ssbxIQOjEhhJkb601peO6flmroYuoOpOpqSmzx0gR/2uWTO/
OyxHoIYQNyyIcn1/VSjxLYRO4Tna6vOF7WFM0TR1qf11tMhmokRt7agMdE50C8El
NuZg7uVPPrisuGwmyEG973Quc20abcenSnlxFC+8mlD9CY4gl+9IAMXnNOGDacN4
NFJDivQJ5GC3u5ebPJ98WUCTZif2arKaBt/x+6OP6HIdGAEnvknr3sVQALBdXSkx
Stu//AWED878KYNrMyuHIm+kOsQqZBHlvze34GKr2W2jdOuj6W7Zofs1+3nqiqnD
NE1bR6wbVXG+0KJkFTMJu5a4tHV5n1QUJl2z6eDkurTFHTOjKpy+HM/oMyvuOCV9
V2daLylLtHkEYSuvUeXfrnKzWbaQ0+d4Ac7Jc239oF97+gzHZ5Ngsw1mIdqKPEyb
zBe2yzYDS5OwI6iZ1BWEqhHJ2bQy0P539fCpeQqv3KYO5+cgLFYNhn2imlT4Sasn
BN543venPKlPRX2XoXyZP5kz3YXOcLyXF6CJjoroqDEvjkylyIzKYL7lOx4vTIqw
kP27j3nmqECvOQGiVykzqAqXJ66IVvYeboQjtgCSdaU2R5jn2EBi19QRUsJ+fLBx
okPSejWtszEwirhSkaueYeeP77/C1ySOE+C8/zyT8qe8D5/A5ahwLsXCjbA3n2UW
51RazNMzQuDJyaT667+2JWmOExDDKCrHUHK1tgnusNcdmB15841ysv6NqM4Ibngp
fodHr8O9FTIa3TcoyFdNAOGpLf2QmgFIgEp+4dinv+9TDY9hj+Ft+Cemk330uz4i
1ge5ZaxFtJERpPwSP6Hy9R7HwtLN+hSwnBOwmTsE1oM2TN5EJuppS6xBpyJGKrnV
TXgR3wNrl0nGqaBoXwKEgI8jjG88Zf8Yb8rr6rI3EItDst9B5zyTcsujce7WVeha
GuPB4Vqu8HgBiKVJDnfEuNdkVra14NdH2tD0SbiScOnnVpAI9nRpsQl6CE205kGj
1BCqX7ULGIGSZmvZKohF741LNSLJjA9DY5mdbLRbgfTjWLF1AYRZtR2Fg/+DvRgW
ZX7Xq8qJQXb/Rar1+Uo5Q7Vn565FwDfR9P9nAEiPZ3u6N+111c+TNgoZQ7bYXHJG
LThMzWWuYAKGFKJclRx3Ni5NGumuSbQaelVYzrK+luE0Vrn2XQ0CLaSco1xg5NXG
xKYT07M/CZkIb2/yPqWTk/U5IZTgwN19W0Jo9OXoePzWAo4p5NWwVUcZCZClY67G
/+TmLV+QfvuDdmWpFfPpjOqlbXY6AJYxCmU7TCIRuqQJZccoNSwUNfDYxnFIks5+
QNzhlLc5hrHYXhsOoI0VJM40brsD5E2ZjMbPGGRNGSTceUyARAFeVPL682k0/66T
VO4ERCH3b2VholaKhe+m+mOuI6LE4vdTTsFqw97EzASVI2IQTnjlW8xHNW1NyUjn
CcUiA/TEpWm5uI6QhBSSCY0r0lAKqloCD1lc8rar+bsxwMwWo9FfimwdkHg9Bf9+
FjqtJprOLIa2pkDGTb5DVimd3D/ZY4ATjOrgJ83fKeSmlnVU6Z3JjLwF7kc3/RBM
fVqwA6NnjeS6qd79uyfAAJYPUIsL8GKZWS5P9tXEwXzUUUg0sAP2e0xlsVxebHaN
S0JcC6hAlLIG5js1BkPHdd4EdFKpDkKtCKjIMtB4qPZisAZD+CX9abTkBO1aU2FG
tKC5DAYzRcZ3SQQdAV13uWABcc8OndJdwBDvcr6sa7GUaZbnp8JWHF2OGxjwQLCx
jH3DVFoGQuQR2FM0Ld0n7V5itvk7MCLMEifUf9QBcHHrlAHjYU0SzoqAtmNbNNLI
FL/9i71S8esIqWyPLjraCoKjFb5eYxsWtzuvNWRUBi6ifX8lzzwVhq562BZSX+tg
+haHGBAX8mXKgdTeFFyOO43mA8D7WnGpY/NHYYHRURkbGK9kqh6ZD0MUX0B3rbfH
5iu+bgQbbyXZIWA8I/MebBrhtByUc6hb4eFHpZAlfnoHxPW1ZGdLRs8CrzDET9+0
aDNiDZ1L5DRbkJLXqvVI24aBbSY7+lA4t7NSmyKBZTGBccg6fA4pYybz0mdg0KTM
DW0Pq7Is/8QVUaCEQC+qfXMQ5UOUagebFIPk63KpnVViBU+bPl/kLdudLT07oeof
v0amrO4TFv6RHCTCBHF3eZicfIoC7XJvMRFib5WXhuOEU7PD+pHm8uKMDuYO9eQJ
IRp0mHkYDkdfWdkxabUv7d9sylxPxoB5D3puhWFAErXNSGPBf3sRfVEkhvFEgY5d
duvYv3Qmo+KSCVXh8NVZVgjXYRUNj+2OfYQsjCNgAOr0j8MS4ysiryV/ZtjRto0R
pyz757nZoPL0JadsNiFVe6qe60SB9BabmCJVmbIlz09CUN0fsy36dRm87cPCxbWq
2YqZeqfaS7eXacg0LJlWaoDSYBCJiOEBJzl3GEtfET+SPZ3aIGuTS8brD4QmwWCW
kRrItpi8LMCEIPJjRj+pHdkaonH74oBwJp+Tnnvh1e/PxtjAHsKkAPZvDB5w7s1E
34e+1581klpeYtttelwrPWWZ+yfIH9OqlQ0SjHBqB1ktBA9YPxCZ3fIMzX/hAZNb
m0P1PgMVwO5eFtoU5t1KAMVCIwoKXIg6429aQBjCXuT5BvhhHv93de/UuJUq+miB
GUkg4anYfplpRqJJ4FHqKn5BgMJQZGi37uMOC3V+LfOEeqSRnvA1o0jG7dJDw4xO
UMXHmnSlHiaQuv05XY1sYmU8CHzjHllczJRnhFwY8+zYBS4sRiym91h1D6yRrG6E
KJDh1w7nL+oHzeKF239l56Dfl84p19KdGUMMc8OKo+Fl/bNm7g2MnyHT6O7DxyLI
XGCYwPaWAvxgTR7ARYUZ18XgKLqgBI40K6hhCl6sjanhBFMKlknzVgoquFD+4aPY
6Ag2BvsddM/A1Pac9COoUvRl6SJ8XabMOOC4IHrQRULQY93p1/7NHDJGE/rV0ol6
u7yE5n6jUAPzJIgqyezn8U3oTmSsYbXHwyAQJRUj1wsP60WI1M8ieylNNFlkOGiV
iKjSeTzE2pF/pCAgz/xA44li9RvROKFmnbiq0GmBOzADbDuJhugebjQS1bIT3m2p
dWp8scOy8leJbyOCoyEAy0HigRTctl8lCIIPS+UXc23Dy9Vq//jzXvXJhqG2hQI+
kdaHXQqHZFBO7gZ8QkjbwXT/EeJvOlew49B1hGSnH/bwpz2mxgkRm2JjVHabwtFy
4D/5yP8dL9Mocvoh+xoJVFkZmjNK4VZ0JWCTZv3Ppr5jSyqrMgkNP7O+aQ2wb90D
feq89MmP3P/ghj9YkAa66i0W7vBMmwAgi9RoQFb9RWqnyHO5gC/JmT+GG6sK647S
o4fCVlIWP2OtOBDyJNOa+FXJCV8kaN8cvv/0RQtDqRVFMpJMzGh2xkj2elHksjVv
cN9B0o13Vcd5WlxOqPKVv+m4Abu1h7qJ9QOkxax2qzl3ukD8eUDmPVrCH3M/tVTw
Vyy9WkwrV9FhO6sHxVXaWiRKISqM0Qw5edKLpY0GYB/TuiHJKHWalaiopTlauxrF
x5cp3pODBdDUvJkO4qfoOT3heLUbVnvKs6xVfg3Mi+d2oMCaxc8fQIX3qaZUZPeE
l1r0gDk9GZPK5nOvBLYZ33bJbtM1K0ZsZqfxSEIptthYuzsjJ1VBkRKVDpqilSFP
20TtWvvY3rMHsLhaTVBBQARKQvMQAt30k6jk+baJW/fOITB3noJ0ow25RQYDeGep
ESdl/tudhP4MPZNILg3QWRdeIC+imjrrw/UyxOZKbgGu1wOJkWGRWEb+jvwxey6F
M+P3hEqhd3iDOOVhGw5DR42YdqDLMIRnsx17mN5xm4OMTIagm9Z8G1aUPa8jmoEC
iMsDzKkFpr6teq3Dem0rS+XItWHrVax4QM1mQ+5B6E+41x4sGCpEqFc/n0+/T0og
czWpJpSG0J4zBJR6D6pgCdpY9jmCDJHsKugDSBCwczeYWEHGAy1fDdJraG8rR/yC
Dub2ZIKXPZmW9fc17AS/j2aALxaMGHJSrSDst7sme41bhCYmyI9uEa04r6le5X/d
sagGsdFO+XGNRQJd9sQmfj+dL49uptA3XDEGKRND0atlyDQNG0Qv/6LoLxdM/3j8
Z5agP2MoodiA5Tt4kVk7gpnMLhDzds3oqY9A3+83KTC2CmsTLifPmSpbQ0ikQIv2
HikufG72NEdiRytt1/d5BIuTjsTVp0zsjX3EaES7KWAIriil/sSj9GJRmxDmctWu
H6buyhRjDnyMDIlK0Kk+RIGE6ZIrELNpBJVADKO6y7VeTzSDk/DLtX/b2ZUlxMs+
xgghT3Unp+gHqZERztI/S0cHGdM2sxPVzw+qJQ8/Ed3oSYmvdWggKelmJKTS8ih/
Kz0Nnco4M1iGF+C8L/eXP7Aozeo+mdg2Xg/RBW1aFAPicTwSfG1YaupJE1ctU1++
g7xKcnTwrVV9rgGMKmvt2sYOCQ18e7eDGX4OZt+dPeKGQrG41Y/gZ4IWonfVTF4z
kOF8LueCHM2PVZOseenbLFRGUfy12VJZ2i9t9zosQHrFP02MvJrcY/8nMiVgm5l/
Lv2qm4U7RrEd6xx7Tbqmy9E0lo+uhWG83a5vG+p1Jy5SqlfwJVF4ZGlr41/pjr5K
XWjT5y8Gs/bmjvQKQUzPhcly4nIj3bmdCCUl105igVlxTIiL8FtxtfMjZMq1hGeZ
SwacdAkt1Iea+QLJsXUytMasirp8uEo4f42ovETRfjoWA7ecYobAifwL5EpDaTD5
/rv8QHvPY3hpI5796yLj6j2GVFUpQgryLk0DmxcoALh38K4S46djbfD+4Ez3X5GW
ECgZdXrklnwngrI1eYzdou5UHo8orGmJVMKmW48CBDxu9Hr/WvUOo3XMRgjixWRf
ltx6lvj2Knf8ccdAgzzLl1Wbbt3JY7L23+XqPZKbMZNkvmyWdTYAYYYt0R27iy/B
bQo2fs5ok7XM9Juh4jGKw+JlDrzsgxGKKrE0Ahx2Ml7FkQTvjEcmzQgu4rAW7mUc
/+zRgmpYSSvJv1kdN85zpugPZaY2qJfz5IoSfJtJ1tH+tSBJNfXN7oa0o+x69pIR
8IfkSZf/L3P2wg3YOW+IeQBS0ZsaQY642A/WV86DVCQdMd39ZvDQMjoUmcpqDedc
58BQU35XSweJOKfoW91Q36Sgk76lwwNyA/GKAGY/U7DQXfYMY/0etD+y37kDYZwz
2wBMhmuX5xTZaEhiPAw5Zo0uWpBkxI0G/95D8xR9oxfoCdv2DaE2MtI1q2QiDFl5
2sWN+6Hhyxp2WnjpE3z6tkusnW7ufHnFghy3fXWfF3j2+k7Xujm6NcvrfaJwPWAq
sHwA7SRtmvcGdoBQuYUHtQNaChMKwaHeR/pBbDTgCFJZel95h2Baqa1+X6rBZ3vH
Mfzr1R+J07ZyoDnvnw2M93dIAphvsNVpBUc6K3pOP8IL/qG99i5Yk7gpUhwkrBPt
HifJ/z/9RnO9qkwZ124MTWLJEY4BVacwluOkKzuYeogxaR9HhLaGP8D2yLv+3kt7
7sXTFVfYI0YuyQ/nOWLRyR6KprZJeUHF9pxLAQpAEtZRz118GWm7XSpDwwEOMiUb
v32hdIwTBJbJxE2/IRuMZjJkq77DuqU0/i3F/DGRttNCGZ+rISSmKt7oSNadXk1F
4T++GwMvuI9OXuGVIXdcj+CKrTZ2ZfHJQiq8XZJB0VKYkaL/AnUZCJ1Bw/X8Dqxc
jAUhHaXe8fxoKODnt7HxCoij/ptQBc6ijNplWEpWulCcMNcRU/LGSJxjQIpO8KVr
3f4/INvGVVklFdxYHsYKZraFNHzu3efEIEO32wsf5bzmF5PaDIUCqWw40hyu7z8c
v3POOhnrB7BLSn5l4PVkDpzRqCFhLg1A83r0LpbRXpujSzf2Vs586q72QVQdQ9yJ
WA1wPrZK33U8ULGHsruYzS5naxhY0j6jvicVoyIJHk9INsoPy9Aui1qk+DubssxD
nVyY1V7wlklrVaXdDIVW9vmTrLEk3LLeGBp0VDJH1O89AuRFKnr+RF2S9LuV3zCl
fUU+CQhQAwNII8M7sJqVrgxRBsQb5Kgy3RC44VhuLsiKn19e2qqalJCbQ7VB8j4c
qWU9CDTuZ5n5myylrkJDL9cZbLOHB6SMgh9zKFzHDjdtn06QtBBw3U3MpOsH4wov
mah7EAEC/xN6fOphL1mJ/i0fnMMUQLqC3wgciGR+/0xJYOBKGHQzczMvpAR35SYL
yrBrjniKKwRPz0mC2LVn7qcZKSYSIjHAOghxBx6kd1g6CYpWcKWi6EYR2Adg3o67
7ON3h566u5ggAm96V3KWS9OytIS+vqi5lYELU0UehSNtzAZrC2B8AHw/SskYO9tA
donimR8zTrn+hTW+cVrMbzjdxcdWP0/nunjaZ8RnNJtLIxg4bEjM0UnuNuoKag/z
njzfrw0ONZXTE+nMucWacLKXHYeH9Y63zsEhhJMaAdWqHvDzw883foNrEiWFDkyy
IOEXq0X91liyY+2wyG52d+gW3Drq/CsWLnVkjghUMPoBCTNGvXZ9Sw+lPM6h4yQ+
LE0lqbb9iy0qPiLGYb0NimgRKV2tbuNB6dh2d9gafsIAWtlR60dQ4yRuZx2/iSUE
kTmfSM53P1xViQ7WvWjcFVUmHjXv/YQ+B6O3qNFxirLv5SuQ+rHe6xUCJS+KJ1eZ
j1evvnfEYm6riHxZQmcVJYFGPPwfJVkBnR9U04kPZnLxJ5tbeCMCwxurtKF6oknj
qT4tI+zEWg4lkA9yuBKs2cciGJnn4jgQjTXZZl8u9i3Z/UFZVrTpZNj5JXWgmdSd
1/k7VkcLnkX1NHaYFwhh0GNpOp7JbzIq6q86Ksgv6+wEOTbq/ScGcE57zFafJoAn
HYKBIRIRtp6ao7SFGVtDR1vkDCRiK7FsU4I5KaMf5ZmoWfKtFaZ3qteQtCdkdq2G
jckde0hA6qO4/luReAr4Baflsl/MAzhkD5AU0widCBqI3aIS1umbJBR7mpGiUQib
yvHzf6S5lQ2uxXN70I43ykPhtcNfgin54/mxWg0ahcool534CNpaK4Do4EN2vtOZ
ucFhEkXdkkP9y4kO19cYQISOrIUzSwf8VI7v4F1n0MzakRWyKqv2cQDClaVnx0YM
e67x4JQe+R+qxitNRfDqrq73RTZUDzj3VTVa+L7cquSJfApOsemRBT9Fp3PvWGXW
c6d75iRSRbCF/EA58YuCBq+gVdZSDeG9wz3YfwBLw5B4Tu7TsZYoxsCQMxRhqgOf
w6OFxpe59RkunpY0kGNFrqNeyOTfSxQTRBTAAOhKa7In4o06pkrLWyc2nL+ZzQ1M
1R5J3zG8ybz1CXe3qapYmbvTA1jtYCKkkTg0YccT3It727PkfE4hP+G52gVgwht0
doEzRxDGBn2kSB8uU6Bx2kHLXNbJKE7/ivVQwsRZk5k4CiJLVbXfjNP3dyh+F+/I
njfViXBq+/eLN+2mDKB/9yaq5T38s7Cq4y0YqJ5jbFl5px4eFs5mb4CnwczSatoc
7M9UfhlantjQ1FTQQsYZHGahGdOtlq96jxdI03OS24Hzef3DWiAADSBWmxShJ15y
Cz5U7AnW5f7L8t3lYB4ZEW+/3vqQpKD5JR9ts08yjISmdRUN/gAc5figEzfLIYgT
ZbW7+JbVMXrGjVd/2wGRy9McXO+wqH2eKTjRd8IyzRlaS5Db135aUV8OAH4UaNNJ
c1K5ysGrBtMyOdRkbIpRuZYqyJiyjWnjcJmsaDNT5a0ZIqO6AULh3EIv501kqveL
iHPueFVrVP4T1L4G61uR9iLFv4/thBHnpkN9yeXlaZ3aZnG4RnTMsOJdwkf4taVb
wZ2SJZvuMsU9/0xEfpWK96xvhNgeu4pB0uGeG+D24acUICHFztWe6q0S/9vx9Fju
1nSicx7A9SfPKDTLJ7J7mW+rVgHljXqp5m6XQyB8s3KynmZIHa8UNHaeEwhv4oz3
j1d2FskcwxT9YpQHSVl/rshyGNCEfV3DdyvJd3Av5WcOJTnH4SHYtjEtouZjSaPM
8YPjC9KnzFS5kqzAeRSMk0tqCjY/3dCqgsHTAjLumYNT+dU3LDBGwwIIQzGBir49
Wri3jskPiindio0z1DYKCascEAajnhD1wlzStccqtv2OO/G3BSEKoRLeV5CzEXR1
7uJxeSPHSVhp6yYahNITFDOQ6s7yfLTkjfDAEnSVByDpr5LihUA11CEaVr68qO29
2ad9XVBLIdzU4V71vy8RnqfCCmTuF2wXl24Tp8UUEGewPrZTBTfFMJt7wHnyjdHi
x9ZzziD2sdQSPMeZxJ/6zf2XAj1F480XFknNZojBCa51OpFobGjOHweVrfFZAxRu
HsTsajDuswmqMpsPDlpqmTLCMvGK8ugl6RN8cdI6Jk9GW0x/rYg+kRHrCgnpru+i
eth01b0e5wXS0quuPj2A30fMiEg+7kMbNVnFVG3o5EWk5CCqlo1AW34LGYoTbOfF
5Fzxl1y4J6tNM4lemUcpf0IyCy8E/weEk2nLUZYmOQtdyicjr4z429KnbzaeEztY
x5YdGaqFqoVRrdn+sdZXGqsu7/9L59tb3ejyDOONvSLf4CnlqBeMW5UbBqrNP9+j
TTmxFT5AlldUDKwwxZPfEQ/PDz1xc8yGoXJmjkknJedi4Q+UCTR0bU/oSh1f3vY6
qQNPELHogQKQloY4TXIPOlbzpH5tiVRA92qLwmlOSEdKf6xxyMxazRzvukxeBhP0
qBwl9scC0ZtsxjrNYO6e70bGRN13PxGs7IV9wFXXjOsXFZ/USvQgDMocgt+peXY+
`pragma protect end_protected
