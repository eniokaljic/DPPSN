// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:50:45 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
de2FKsCR5BrwWXUccjon20IXTpl0QC0S1t+ohod9wuVx0EP/j4jh3w/7TPQwD60o
R+EniBaerkpLKNPGZ9rKT6rjjXlcmNTjNXprwO1qr6hXM5U5gNZp0ZNU26QX4JXp
OeeroNYtguDwQmhXxB1x6IbI+VpumijTNIhs8QGAOMM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
gf4vTY/H1bBH0X+i0oN4Z1OeL439N/TTHuOvbK4+g9HiZr8FhoDDW20CCspEB4It
UUniIq10CrJRBtyWQaG2FtyGM4Urk7XGQiJaNCt9Q8cm/TDDaNUGQ7vqIgvuDVou
pngPVvh+ZXM2R3hvvHB8FL3c6XJxmCS34QKTKdg4xDftT09ny94u0JZslBZt8hkE
GLoxVl5TqmMRaR0nX5pZAfLCPMUCiOvcUrHMBQjXqHzE9v0RjAdMKXBTzKC94g8P
w4rBVF9P9k2nZpNRU8fE+ei3tHfNSnyGqP2spAB69wPnlV0J5nwsKvJ2mI4RQgJD
gezG8A5/sBFJ9jZNdy52ekNT4x+PozrPS/xbIpF9XCRb7f4ecJYcuWQMmytu3zId
uZIXASqCkgjb/zNatOyJ4cjwXGnCjNFJB3PWKpdb44VEz+k1p+nh9FkPeiwucfui
h2R+IlWZiv2jkNFei7ioEUv3HiZpg3TUBiMf7RwxNb5O/N/LSsf4UUelLfdYIAG0
TeXNYHKIo2GEyGG1ZDi8vam5GHT/U61KiQHq8mT4N8Fbuv3FiQVFSBBzOPgWogWZ
P+v6v1QFIERCaeyC2RiYOp4z/e2jYEjY0oLwt2svDZ+BEdV+AKsv39gaX9sTyQ7W
ZMM7jrcDsbhV5Rs5sc93nP9CCG+Daz/kJBvka2FqCxU9dmzOPWeVhTdA8tg2bNya
6dg/cDSDUp3KFYElFVYzc9xc+YYD6J0dYsnH86UQLmfHQ1TrlaKMeb8+eP8JdhVu
46ch4dy2O3i8gWl8JAzkGnc5NESFcQN0/Z3RfMTG6T4CfEXrxtuM1i0n9ELRTpqt
F7zXVVFd6IikrvOlBDT8vDhJk3QiY7n8DEPYfmmHF61FKpVTmox0/u07LljvBBB0
vF9PuktMsjrLHEDO8nqy2UcC/MyusFo4N0q1CPBeD8fDcRThbZNh89YEEONDalKV
2Ck8p9YJS/DwVKKDxixoM6g0ZylubqJqJr/zz9ZI2H1LWOWq29yKivWJ7RGJUBSc
3bWIc2AXB3QOG1vh/9+pGwLfO3yjYg23YfZMu47XI9ga3kC+NLqhghQ+rkfXYeU9
fElI4+9AUuTtIcSiBwq3r88XtcdNBuLKkKSaV3Yue0lyxrLZAQUf2fr2HzKLKi4U
QSsgbTpv+aLwDWMiGC/I0BqVjFNbVL9UtQLqNCdg+jv5Jt0q8ryJcuTWbsdLABW/
HZxTRJHrHglYDBilwtllz8SfORLH6HoD1agonhZh7hwziGxMt0HXFPhLphPuDXWl
VLsf1BbgX0d+XtALx088zNDFOukc8wkeKvRMIL/04RXv4sAVRoYPXmiU3PiZ0RVy
k7fucUNlwRhTOYMX9ltfG38E+k/kwAo1FBG/ZPe/0S4F+hXxJRcKFRMsCvFIJreM
wIetopYuUoAtBYq591pXRT4qkEPTMCgvcCymVefJEtSk6if1bw6NvLWXBezhRhp3
2N9cMi8zLTUHepWiHpgwXbm3UXzH537RGt7yvfWbWsv85qU8lSoHvv+S8x3GQ6+J
y9HlnEmmHJLcdr3+aSUvmtWSIIPMd3SCU8uPxCqUaTVnEbcooHP3v4hWHb7myzFs
huWyUoD5v4d7qncChjfqCiZv1KOU4hr/tE3eHtnEf0sm+zFjMn/N0fTALSzz9SVX
MQkhdT+MbaG0ZnQZpaoE83tOsmlo92XMCO9ENUp5Duu3sF0fy9lstUkEeot+HNuz
Xp/bLEBc2E+8tgi/Ied9CRHR3GfM2PE7Ql1GUmZ3cTLcRXhJd2Hs9qJSY2aBanQt
PLrfc/dCBAhpPWG8UkOEsEPoj6YutN1Q7GYuxzgAVjZRxfwuXzRtW9c4lwRGrf74
PJ6tiZhkRolx5e21Q/8usPn5S5aKLujYo4oBqiCADM33/wFaODNaey/mMoxHh2Hd
OcnEZRYZItXkXcMyxgB8O926+f+jU1KBiZEFasGvHnrq6PSZIlz0ACcC4riAI/me
COkyC0QuqltCf4ZRbBUq0Bcf9fwkedSxnv6YAuCUkNOML2/yV65aEj0WGKxSjUeA
qNPirPqxXzDQm+Jlj7I1G/3TlLJYOiComX0WKan9iD9s6K6O26YZrRehQuDYu04b
LCpOA+V7h+N5EwMPVNpbR5uS8jlerJd/tnpq5sDYGOtOUF9OU4H4bT9XWVvC39QU
4aeHEUt68vzxfWfOLyheLIbUj5LiRpsA8GiEDyoCuuyXCo49ul4aJL8fh5yKLgSm
HAQZlxG9qLY/6eXDg763dMMaCo05REsrvsKRi0H02mMNr2UmoDZB1icrGd7g1w7x
fTmny0mGl61NwEqcgwVfGa7XY7GjvWb9E+pB2MhobCD0UEaxVjpDSA6NO2b0nFT0
5r2GkOKiqlkme7OevrW0eK8I3cREQaJXDpJx2+GmnprVnTglE6Tekr4+O8dZwUGM
twKkDBdtFqg5J76TqRGPUt/dQUHcax0u1pdmNidQYSsxi/xcmwg+VMOqAz5exvDl
owrYU1HrQ1MbVM/YMTHoMYB9dEgKbe/qxzMZUIl72+Wv0jStFYixW3UNHM86sKPT
pr48NV1oZ5vdCSpts9okV1R5xhD1eCN2+9P0IUHrbiugK68l+x9Xhf7w4weqhknh
haALKUt4gZeayQ64goWs/qk4czUHV2kY+0402h2yiV73/VuBAFO/EjX3bAdqsUXg
KrhWdVHLVwomDXVbJO7AlrJabyCBAWQc2Bml56r+0oMeCmvoCwL9s2x2N6d3Fkil
+hvOOfoh9Pokp6qmYW45NKrx7hDnC0W7GbwQ1dzs7nC9DhR8+JzgR5Lq3cniBTLp
H3gt0/tdJ+uvDvTK5+JihlRoXOq5BKIIYrVywJ2J5Rd8TNjJBYmlKAgOCuPEn2vu
b5LZq1eSURA8lydaSYJJJdILkPEt5mNz/U8Hyktzo20YARm0bPiENQ1MvJzugzWT
bE4kfcFxet8jz8DOmSPuFYcf0sULnjSVTsiO9OMXC9Hnl1wlw5PQTso9N1aVcIe/
jnw9mqMB27kIQ8ZUpGUfLqTAftLYa+dCnvGd7+Dsfu2UvLckpwJ9snGVshVo6zWc
zQF+zqLQtaIk4kIW4uNCtmRgiRgHGCu6dShS2Apsn3SEejxaRq4L6jT2GxMG91nJ
WccH0KVBQvu+JzpscV6ugkmn65mlOPF3N4hmfhvAl9Ohe4ljwLObpG1LOAAk4A4n
gdf794rAbPYrICbLegeSUMufG9h9Zt+tXyVPbZcHLETGGoiTm1ZJ8z+YjE2TSUGF
NFIViC3docRmbD7JSB5nG9M0aMuUbIsxRPhzxJBx+bDb0jEifDHKHGwblueC78g7
zPcQZC0EDeZbHNe6PyIreF1dgvFaypz/687JOxlSPv8bs5me71F71nAhQXmvVIB8
NxNF3dy29cyiD6EH8yQT69BAd6N2h/HCLiyR5QKlWnXqmuFl+MZMO7Xjyp27Qlz4
9Cs59j5pK97aasXTipq1HGLjo8w3tymD1q6JXst7tRdQrxxLwlFLWgiZLFAhM1F9
kkTsXv0lbKV2bf+tG6upEstAuuFy7aX0M/YOzl5cbYBNemq92Xtbvow7fHiDyJD6
Ae0TzeRovoebIrQhs6w+N2YFxR/gVzWWoSSY8D3XVp6BTr2tO6T2iipt9T7iZyri
u/jD+xHcdFhoZLhDI99S3cxbqSUI7dixuYm1HbNuOzoqXk2JD4HzE60dV0zlcT2O
v5kY9r79ak9k+kT2wMNq8S7cHZV/P8kON5yTj4mpYWGQUET7Fh9RbZwo45svNm2q
RKtoRL7GHDTew4Zng2gh0maFG15KK5ZihAw/HLYYrRnKd+PAn4tMTYlPsgmTO/3U
KIG4SIFLvYEwwNqqBpBpGEa1cOtrTX6WaXgoh3Xtgu+NC9nHc+N0m3IB9WtLhVtR
XVZ/atgQN3dRgcS1oNI/rBbra+gA29VAY0iDEllEV6Tk4E9v1DePBl5TLkeBGkyM
xk+1UviPSr32JmK2b4H12SFFmmt+SbIHK3cg3s/2NE0mXwn317xmM1joYPmANW8J
ky1wXxfNv+6gLcvgnyjngLkln90Kgf6uZnZnvf5jpcotaydrU7rdF5P4g7U4Wv5B
c+Zmj1ZC4UQXu+BUeV3v1LJqNecYg1+4wdYEwsmzDhtEXWgtbXfFAOcmhVZ8xP/E
uwOcO1K/qC+sqOETS27mzIgrTOj1uOYAs0OAfRQgx+PYuTcKNXmFL+BDVog5D+xT
0o5NlSwHKDDejNEal2cIruImdDJ6xxbRzMAFyFEKJj/o2KF3WX5qwzZWxvgO7DKI
RHY3B0qARbU/+vRF15/aBGO83dtQoK80dMf8qaWTz7HPO85zjec1FPOv1ywfntaH
TuyclHZuWEBW/oxMX9aES0v5eXsoA9e+z1QubXYDRutOmdUWOE1TLkKY6NHN2Lh8
A6/wOGeQBSEZott48Zo9l9l5YCoE329o9RAY9QOagrPmxI9qRpx6Fv2Map9EhJM9
LBV2wFr9WZvk1iffotntrACHhsdxqngktD4ZpE8ifDMbj8JuGsNPg1M83YNEBQ7b
x/lIKMs9jLjdWwoZ04Opn2fn1l+o7o83iDJlh29m/+X4YPgPNAlDNzxeU09Hgl2Z
JevBChqH+eceq7UrR6OOEskT0i6lIgWbQePpAJzW5mHUhjS/pMy2NhDu3cTJDNEG
jtACnztI+Qm7D8WRi9j3GKfvglvAA5L7GirEnY51AHpSZ2qX5KvApgIDMqXHxHw8
1GQMLQp1deHbydKBfA26eYuEP8e+UFN4L4hQ1WSCnC9PTo0j3Q2vq7aJCTo0+ZYN
j+EiupqGapgJO33vX4ic7+K28EdthJcFVGzken3IO6tXJtHbLMv1iLJNX/9et6W6
cXVSkQj9YKIYK2guRYBans2daJ1Ye9LiwVan0DPfSjR10WhQV9tL2O5Ylw2yGFqj
E0KlkCp8cb4Gt1bA85LevULkG6vqFqRVM0cuz2XnrPlA9SbSvjhaxrujtEoVxYil
qxtRpuMmGFEpgY+BoCkowpSe7rzA39epbmwDK2PTIl6E0SzEoQGUUe1O/dXBzw7H
P3fOGlF2ERKoq+GjPHEoPJ7U1je431//9Z4AGbswxKiBRgokru+urb5wud3ZFoCE
y2gcb2khFekz7zZsyz6mwEYvhf1nzgOdbDDkZWfcxTqRpqEoEFVNN+zEKqrDMdDh
7TRLCmGSkBlKLnKlETjdcoiA7ev7eGpYK775i0B4u+ZXxJ4p+P9dWX3EgQ48GPWq
jFY7tcyDt/57qzQSH/DltCGQwWgjy6v7db0fQAPZOLUn+VJGa4Q7unoS9hySetjo
xrj9RFRJYj9x0mdIbKLjHMVbVuSyIeLzXKo+vcQ9LN09eER6xjOT8xjnhwH+KfD+
np3LzWR96mY+W/e9ULoR/TCCKKVWlVs0y/V5Csi/mVSLVe64+W4UY16FDLgyHu1+
qL+D4jU/hsTwcAulkpFrPC7PUqrRD6HjLqDwDiT3A80LpHaVcoTKmd9+RL2fAhYB
JQYpCNcglwV/2okiCXYt3JVgKHK2ZkO1J7kOmgLd1CHTf9XefeIEVndKtJWdmU05
tbSEMZl3gXI8l9ZGq7Q6gLsGPu8m6+XZMJk2xTENq3IONs1BD91MNfPVFwoVJcKn
2N7AxUkwlZ7oAZQiRrdPPBfQmUM8NyieBLQeplTg2V+ZS42ZhkuFXiipU7fu8exN
oWsFqOjrPjV7SFTSYNpgV/5w7GE7J1jIb88x+SGIsyBqIc0D2PJyTCHasDgUloyQ
Pr33Mm2Ivwt8OMGGoZXpRmFgDmZDr2zN4nYfAHE44j05eSo6HrU+BbOaHnY8Ibc+
j4TySp6/E0wNcJoOSJQw7P3PgaLynxt769u7EmwHu0Opif60vULkEi8DUCDjVRsZ
IxyEsgzh11TTDarZBjCLCgVf05QKVAiUrS97h2SW+SCmNzCEFAUTYa0GQqfGOi5j
IvA0p8VLfoX9ywjLmb+88V6HDBCjB1o+9KdUf7+lkND10vQYRAAHRtFLyT5a4ROm
njVUP7MQYymy/zpponS48D4HRAIpwct3xJqQjb0iGumCtEFKvwZRqPsPbhRith9y
Pk6lMJdQuXHavLJag1Cc41fOfIH7tjO8u/AJgRTNKbk3GSb1JOHGiKBcYfREy606
rqNu+Bb1ZgAeuBalhGw0OnT2/9FoiMW2M/G0QYYk/Jq9WCOnATX14rq/QwoHzJrW
mB6baOGpCExbjZNj/s19mXh67HbptIoYBJCxKcLIDKPV6cV7vBt+yE8Sksy+Eu9p
TnExBDYBr2iKZOxHbVQmfbe/Lz5CparzECOkqrc4ol3epBsHENCLLcSxSvUYI42C
+sr0u+qrtqwk0DpFDiuhaRFDxZJ55t7APkl+tplIjD9AF9KE9JoIOjWb0uDNBwma
I7Uo2pDj6VjkMmeXMUGcXTblyp1lf0TZhWoN9oK8gSzcMCY8oadqd+sHwSLuClO8
P6zV3eVWLPAJlCHtY0p3HNHMGGhzT0ad67p5+7dYtp1I6B77Pve1p7NZZWfoUD3f
nE4IUNX5w42M09yyyzSa8XmsJstSDhZre4pBA2gnnDTJe3DrEoRQwYT9W3lwoNFl
J2jGQ7q/kxa/w1pMZHEOO3mATQaE3my0WX/XOxZ/YzZAzFhupB8OFJ9QNn5b0DHZ
43nRDSuTe+7N1MSU7nVo9MU168Zb7LJn05taXRlURdTyB0qNNY+7CdwzxKswrYnV
HVYjHhhuVS/VFvXYMSeu9BJukt/AMi20Kk6EjyvP3waMeKTcjM24Vj9BmuqLPKxP
vNP7sHXdSucCMnT9WaAqDNr0VllBYZSUmLBbIgGjRmvkKjxqLmb9IVTMIf4LjGjZ
4Kl6y8xkhNlsysX3BNHUo9zC5O8SC6IzcZ8plQE8iS7C9DCx9IzGB1a/GadHlqRF
8nANCgbjoX+rRm6C9asphSWfMBx3o5EqAq0T6FIzd2xwJ8NhdyRRofbhKwFofQzK
3JVgks1MBxZtM2+vxz6bQjFZnmfxTBB8V48kEY811TvrSOn+RDUwgCd+/32fbXEA
1GLXzQqYj8zg8VgS2BYZjjo2gyWKgc7XCeAY4wQ/6yPzRAXePHP6G1hkE6Sc4QRg
EtHD6khwZ7Hjj5eBoXWsVVDjRJFA5hcuxlWnyw11R0bFD84yl998zPaNgFhcY45B
+8RCTdWrWWEI27gpx4kkTlpuDhD9h/1qyFTvvrMj5tuPzqk0XWae925jQ/QcB0hq
w82EcBB2iHi3tJ3zWcP4GIQ37aMmr0sCuGTQHvLk6ImIU2lwHs201UVhNqdGaH3h
hV6UF0OeDuZloUARwpovHmBJg4PAyYOmfqsaTLSC0DGBxiLAI4DB+FgWWTEHTqPP
wJfOuk58W1Co6ypOSfoUwSqZAXFTUad46MqAGjqB3OmGUNw7PRv25LfXhATMej5F
5oU977GvGF6baYwLud0gt79hAiCWSSeafDnw7M/XhEw0ZKcquRJR3bajsxI/oKAa
VwHRE/5H02M/8Ypjr9xCiKQS92ytjlMZCsKARcfAn7y9qeY5bF9WgizL4GhNMfIY
cbucTvPmhtPxIIuSopB4AEN6UZDAhKb1D8aQvI+UcoOsQQk0GtR/pmAEyft+f2/N
134m+qlEIhNhLQJedXC8ChCroG0EISCfiwuFp+HRXm9NujuZTzkkV+UUo6P3KgPw
tq1D9/WRFU2c8qW3TkB92oPpPTN3VEYEE5yWjZewWW0=
`pragma protect end_protected
