// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:35 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NPqDdhiBBCe88jnR31JOj/8y/bX2Hw07Z14BAXL94DLUoO9Rf0QlzCv2e5h/eob5
QdiDu9z71Cu/2Bf4Mq12qOhH2qYvQB92Boox19FEFtVQuIpqHK44T2I7UnmmF4AA
3M9X9GV5CzdiBUWUbeLdrNPX5qH6m0+IelzTY5rS2oI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 324336)
EynGpw04wHqNcdQ4kaxK5sjsbyjKvnGvM1PAoPqYNo6A4VbqtEIbgQZ/tdTV3Cwh
jHFa8xcpFv3XyBw7y5QHpMsvm5qQvc68OaLxU1zx7VPk6ATqX6xXJgdv+zx8MnJ+
MAqgtkRb5wjIPQk3+SGaXAOlc87egn8onnfWb0FkhhStytAt8VS0CBjvELx4/mc9
Ki6IrNe0IDHDDKle7zW2NafmkLr2vdS7SrTrsOmabkZdk1XwdEQJ+eL4CmJJoqfm
1a3pcedvUiMOBpqPAqhENFD3pyhNyIDwf+H+yMg9KjMK+t1xR6snuZeLEsVjIZ79
puA4BPgMorHm2CKXL0VJK5IFe3WBlIxcM+TjAXGbB2J2nrtQJLgAARf8gPBq0pYu
/AY/sqnebswtLV/LE6YGNMqtHGqqywJB2XwnT5AOpnRdLZcLFo3R+fCYnLRfFrkF
xkMTR0d4iuTizxvuDXC9nTPQQptXpfqO/ibOfflH7LW1vvqpiq+GgLPf8G3rx0rK
04wp0Fbrce8GLeYc0C8H0N5DwIqaKMymrTOokFXaHwmgqZkUVgMfX+TIhNHhvfsU
KdRt8G3WYV73ZL3cycsPqJhG3s87qZEZMMKn/suj86lCKdFoGgbTv4fEs/4xQTLm
FUwMsdG8D52+/pWTjkuDN1ZbYVtVXvVKwFGZz3Vnkv5GLCpIBK+EnbvVR7U1B/TP
bgcoYTHJHhZbgkIES3haQkR4Ijoep+6OpqlszhU9QbdOc8/hzsLwjyAIlhD256Pb
x3IaHVi4k7fFcvlBAm1++oQhRSNFX2sAVXif1b0P8jtNcu4H2lJlFNvvHTv3Q0Se
jgKGDY9DZpRr3G1s6iRBz8X5dZe0XeBT+p08P7KO72Q+3g1p4dC6N1PijDGMkrDR
4uILyKs3j1Yrl3vzpF7MTNo+i0z49vehUCmUwzIlQ4myBWtK/FPPtkQvzPIWJXsp
ei7z2XuBNSVwyk7ZSZ+MIw3xL2NFUWfP3PEz7f5hGqSw18Xhlc3d8ayGjXgFPXGC
5HlM1GHgSifmBslSiSnGPlvhJzFRVMhBYN+URwVV03VGTM5YSeT2+knF9PEUXyoW
gvbv61cG1GrnvV5pHrReItKiJpYP1XrQAe5lX4fcOmZLn/WJleMk06Lzn1EFi89r
uQWVP/W2bLcXc8r+aRLCjkDDhE4ib5cn2qlv5LwqhW27uvtCpqwryHTJKYWNboDp
3qag/sPcE15cBnhXUlAO7Q+B0qZ0nXzZXONkiVnVPRh1wPAZGN7J0thKQ1uPPlah
gkTd4kCpWdM1XqNNxtKwNoH67IUOhLPygICC8Ejp3EltwCEz7RN6Yo4OhLM+5D/f
sHeG31kqvKKtKX405LbyyQWlyyz+yJse+fux8qZwaAzYBtLTNNMQvK32qdf8AKOx
csNuMAgFYjrbgQ6nGsSksmXo42R8MbZSBS//mapt7GtRlfZHmkKDleQUd+AfRPhQ
lkwXIWAoOIPoZbfCrKkgIRZUIi7fm8OOFJoQvSiPEo34Ao/5gtIMKSFDOD5OXjpj
lvq/O1uvxJLu4qozqF18FYgC/aUXlZhKA+3hFeqauL8kwnwVLlKvznNCgBmMY0WX
xiwyXheREg5sq3gQdzEMsvDwQj8Ub7gRiBy0S8xoSswwyUfZTrDnuH+DFb0Tg/Kl
1LocyBTGsCzJKW34Uf9kPmSJhw4GyT+AU4xLTe7Y+bWgahVIeEUkNtszZiy6uDTD
omIRoNtdIOTzOQFwh7AhJBcfKUjGoeDBZxxo2/Dj8jGwPFJkuZosxNpFwDb6i7ch
+gxXwJ6UcJtj5B6Vpd/QDxrXvr6JFRGsM/9unMmTNKoV0cmdOQidKw10k/5TmmPb
5lvqXiZf4Ctttuv7U6TP58zLy9E28e7MfQdn10RjUHpQ6xCi1Kqz/KvBHCJz7+oG
ioujBILcvpi1CVDWZI5CjprfB+OfwejAePAQYA5HAQIcuiwOguudzp5s6PFblGUB
y4ZNCKhNLVqNRvUmUx/2aTYE85MdYzffIeyzJb3bQR1olPNPKIt+ZUj7FvKrN46e
iVR3xI6vx5gF/BGma/U4wfkFaJhiiexT7xEC0vclwLDlSrxii/XIW9wwJ34H53+W
tjaGMXKjPHLL6iM/ZU/2Hid2HKaxiF4mbZZtx1GvtD+AbyClYGjF4jnvnaSSMJy+
UJLaGihFq/aohD9X2JF52/CEqtfwtvaTF5niIPWFIdpynCPkQRDaNSQ17hZy0X59
JlrFRAXNS+9VtUN687J05cBEPmuIn0ZnkLdmMMaUeQiE/61lWXObpt8ji/VzFAeG
YhO8mw3B2xa16oqoCyDZHJ9MgU1UFfkdIf5TLzmd7co1c2xUsvMhvbLUoMrnGlDF
7dKPjg/0G6gsfhuLCoGKlOe2AxK/btMk4TM/AcxgVWs5KGLigdcVwvK27n60foTf
UH1TQkOVTVk7iosjZnmSikMaGJ9s+UPkAK6thSbFsIGxCNBVyDcLAILZUosSnwFw
LmZLqN3bGcPY4SyEhrxNaiQs9O+FmASA1sSaIP5/H+qWI8v+Ys50eykJI4ZuYkuA
A8S79Xw/498TmvfqTp/SiImRqouz+gsTNkzJphuo78Qw62tY57d8CqNvfLxa6NTd
3DWRsHPWQOgF7TqSqsmlTc140Zit2yvAeX1Xo+Su47o0h8nOWFHnfyCP7MY7CT83
sTc0/Hb5x7Dna3Td38xIl03Aqg5GrjiOlYz4glkIKHPOWLd93D4VaEmyEN6cnif5
TXVdoThpI712Oka/SY5JJ3pqvLIWVOo3EaCZv0J7on4Xv0VKLDOGFegkPMeWxH6S
qSq5ZhLWnuYIEqHRrGBF1c/ZqHz+vmYyz4ezkymYpv7BaH0wCz5lqNrUJhzVGtnd
8aibWjsY9mQXWs3k3RAIXS1jt5EjaGilkOGrEoABysVz+GtrkGxpn+FZcKKiPUaR
li+axJj10eeIzW2Bt6lItsm5+o22Tp+Yknv1o3l6JNT1V5dj5XFSbtJuchz6AlAO
VgeanZbzrkMdze75k+Clivzec00pIPyddKdJ2iqk0FtNBQ5WJ+/G+Z/KQmrDVUoN
kxJGqP2+tu2C+291XAqjVlPSXnkd2Bg4iR1w9YQqgcWCmd2355lbpkaQ/TW7jMv+
dwSmGLjEsH6YPICRrtQkSfcrnP59I6M1/nLoNWqTfARN5p6Mgr4SQ4eUEuwRFgaJ
SVL/8FPq0pZz7/7fWpfQuT4Dpc40b36RN6HEmcbCj4M6kptCA8trbNqnGcT846At
JfbAy2bSsycS2HzT56zxsg9v0FuCyMXwldVlwHVzFdB79Jram/6c8b2Xts4oz61C
wLyuPJlrTlG2ohqwtvFLA0xWSVkjc/96sRd4qrNBavs+Ee8s65mYuNDlhroEOTWu
bWUzTWVAmqdsYEcOW0u/DQnxeBjdcJRLkkjfuTsOofl29q5wMTwF2RfYnmoU7Ghj
hHZ6voeO+TzirB/dY23uFUjIz588dVDUzivKehvOKyiGMHF5mFdTsoCXGlY9h7en
n8M6lr399NSHPpIEfDGxeIegcvSvLmdq+AYA+wW47o96otbmWNL6FShuuGol+HY8
uYyzMg8ZCNQYU+ZmcFP1OMG5WP0QpUfARFZSyVa4cj+5iYDcFF9tfZo02edEpsaA
2ys8gVUb4LlgVp+xBOoaspuh6D3eXrwyPoUJCYypNc4RW/loTLnDM4MJxjkZohWq
1vR38KoUpb4Q/TCBLg+m5O1i2rfI1C3mHmUnIS7+xOVS82MFmDfdhNofSkmBz188
JF3XBPCLo6iWAXT+P0EF0U0uu4UPxXhCCBAvuN/rycC1ntA0zaOj1I7zLsGqT3Mm
YmqthAJdN+lkoenIo4s7MCGpaeHCqr6rrB3kyO/gOTL329perPwPgS/Nw9qj0LR+
bpt1TuiCXCYjjw/Sqv7R9FRaF2lIJN6wJQS0f9NY4i/GAJwmhaZk7117qT6IrIWz
puM7jzR7nj5H3lGSfMW3Gbfg8e0Qis21BHQI2/Mu0Ems6d8hdYBUpam9tTHvyAPp
4l2g3JfkAxq56J6k+ADI3kwJwXI6Jn5iKTVStExM0aIxtzcwU4gMX+cwu8PJTJd4
zmzKCHE7Hc7NqAsAC5K1HED2K0Qu8Y1O4a0bYq+ErEM62oFVZyElG2vDjRVQW/we
i7dbMsjgtaPFNtIVIeff/hjuOAIelknBXvZz6GK4EwW6FBUYgBvnElUVlcfSdTMZ
WsEV5r3LrMDYNeAI+B9cTrcfjX6ArDi1mRKAnesQNzjxpfs1O6/1amf8PGvHpyzw
njUeQTexpgrh9ABK3FkARa41oWGr8k/pctVaJEdXtKMNeZbc1wWwOTxg2ZQNkF8w
rkTqbpJgCgZh49MxBwRW9KKRlyydwVaVWqsr5O1kJvRsNTfAGW5pJW5+Ltuw14ag
cCfxiP51aggGZoA7s9vrF1kHTsPYLheKAhQctQ9mvzfxgL9PAFKf1AGkjBZkDkax
nTt5q3MSf5B8DaWJ+biCc5HIxDdm/V3iDNWFZ8ZFK6L/utDjJPwFTzqHgPQ+75r/
LsqPXNwbS3KZ5pOvrNfd7BEF1upAz0+TkZDX5kSSpEm9n3AaFQC7NjDpSXdI30fa
cPes/YI52CWDhGCzJGLjnsCnFfInXDBNRtplIOp/6wu8njsprPs3ssJ4dTN8rEo3
Ho+i+aIDDN7D6BMDRpe/A4/jqCX1nkUKzEAecUhz8Q/kKaahkb5VZ/18WB9SF114
xJqajKjycAyP4vtPtRwxu1U1/8v2a+nb6zLIOsZDmLEQAAgXlf40XA48dErynEal
gSW9oLSR5Z9pktIg+WKGJyPRPizYNbSpVVDNTmC/RBxHbKyQMTYQySj3ZSh5vI/s
2t06C3x7UkLyji7sEWlDms2cPao07SyKwgPELZ4V4AcO0WK/zTwgb5ORm0JIh8+a
ppPT6LpM301QjsKVojtBbiVFx+puE2TELfAlvDwfHri+dPzEttFRRErZHrJPyy+Q
Y+qKO+8YwJxj1eW2QyG/w0FytRJZtmcpTLVYXFocvbV0otg+8hUtjz+OqMNdfmNu
bH7K2vnQLfUHdS70Wuq0j+HvZtqU0VxZ/OgfLCETGjZW+KplVN8U9nnGLN6upPt1
rN4Vf0S2xdJbtqZGUVT/zAoorQoaToTLqiQDsTwOcySScWQ1tiVD3i4aqWw+CCiu
G2LN0whfJaePHgFQKDyz4DVlUzsM2dhKhjHXdZsrmUVKB9z+JBr/V7klwCIEDMaq
7ZcaoaUG0B+L+j1AMl/Kgw0SmquvZoZEmdRgxppEBBKxdYSU3SOZJM5jCqtPbCfi
Y8w1d9eOicnEj3BNfI3a193MFV6+Xna/cnLnkCSq7/lwOcDcN7dhZvhJTphLM43u
QMAHzKb8cjV0ZIyM2yJhHI46NUjiFe57g+OUZBLAFduaSwUzk8kJVP9gNOynJL+F
FkMiLgQ9XSc0XIalNk5SlrQ1YczWIFbI8pV3WGY0eFzNWPh6SId5GcW5O31/WDwO
x0ltkqKgSCAO1nTLMR91ob+ZM289pwV39b2sbpcB8rkJ26WLVnb9YybzFqGXJqp5
EWOk/qXy3skam7DxnfqWJ5XGBgEXURZ/vifBkwq4a+9Lp3V3tmRRW9D6FewVdFIQ
QYOFf0jGva6jojnDOQ6AbP4vbp2MbL57pDnxuRKu+a6WtdScvVmVgKp4+m4fpbPI
J9YOPMhiSZEMAxReawabbJyHEwgt+Zd1vm/Km5xpQGUEbt3c9cXAzP1qAtaIQhU4
zKexUjLICsmPnMwmPNybjpkHiTm6L9vGqIGKFIZwfYmTesrZo9w+L+NoDkgYwXgW
L6AxXMWTnmo4b4sNTyNhoINplMQLua0VRPYnSl0XRbgY+NPf/xia5c/E6wgnSiZF
/ADID3tqALHoZjcpKo8BscJc1NYPzciHCj+Bklh7wdDfT7GJJmN7NxSFttlNMwQJ
PysgDlFc4OjVDRmRgodtPgJFuHR9bnMgLkUp1mPFZTy4YnqMBjBv83qOs+a++H5K
SB7oKmri6TWnNq4I67T76o8zrf4Nom9vtShgZr2mwj2ObbRal5uE00/zWNBp+SNI
5QF96IE3e4Az2KHHRMzZ9wow6ysDF/N7khZw9dv8ISPRc0FwSzcCYWHHCcxMHtTc
0Ayb0KkXIhgsLRPOu6tOio9cIFiMYmk9ULYOlGKJlTTL/4TuO+6WHmORkdDqLg38
BIIN1r/mmUYZZ9z7hVd3uYptj2l8ISmXVR8eFxk9qzcQXZFMkL/79S+M90/0wVT7
RcXbTrJKXd5/AOY/vb9h4tAQ+GwPm5DVKe++3qJIVWEV9CI/B5tlFtKTOAZ1xBZs
2liS59ik8H3Gx6iwJVyMYlU0LtIAf+3Q/ZPCA7NTevYOYb4LCwAknE8FXk3zbsnx
T5Pswn0xaPOTtd/j72KUlrvecLSJouUpKWvcJuVgPj4a+TbVt+Q7l2VKoewr+Sqi
PmRztuQZHtmrSIpygWrdId5WqFksRoQNwt2kP3P3nVL83JluSxbwPyqVnhoRFE/P
Ojs1nIKNZeE+tM4THax9xeZR98FEN3UtN7Qy28Y42tU/dE/Fw5lJy/E1b5n2AeUJ
hFXyJHhR97KxUH3oWA47zbf4mW2E4d5cVOfR8eracPz20oICVmU1EgP9NOkLB3r5
OXG4SIAuG+b7qLLux5FiFBJNrpJgBnxYsWWWDoass2YMsQ9ZQJ/2sEQ1vYrAC5t5
GfJZHScGzNVmWthwyS9Pei+qtyZ4nx7UMMC10ZWwYJvMUB0ihs2O8a3eyXJbNC2j
8YK7OMWSCJJWlXCkyRtKnn53cMfA9iQSTYCzjtXONYBxFj7+tNcUam6UrMNmeWA8
3k2FgZ/rG5l5XM6Fq+XaWSfPYFKmb2bf9TW7a8sfk4xBrdYpDBFz1aHSz6aVpToT
BN6+lDUw7UMqr66NZHUa0ccqxaPVyy5592llopFC+ZNSsqKX7qoUaxyUJwBC/2hJ
77QtCfvB5dDgkUrI1+vXJvIF/SMZ/sppNynXpVULMAhTZmtrXz2wLxd0uTcyWVMD
c/yHc3yGT7qr/YGz2FxgKBTDi1JaEP5EhTu6tooxcGjI62NcguYcYNqBc7fsjYCm
XwNGmVOzh7BUwEaPWxeAZpTjPFpW+BRiuTpGTjk5ay/6Q0hK3F9S29tFmSDqQ2he
0HEcwM9kl4hIsdaBdH0wewqFh+YTxcZgz49dE3/tKI3JltCc37JMDTN/HAy4xbde
9mz+J4ywK/inZsJBP/CrXWlKm5WJnGdvlCqhSlcx8lmUAOIXj0j7z5BYWVSmjtAE
9aY8NaPFjCKGUNAysNis0nDidX1+uLJFPNslrG8fxGNUZmqSkjVY2kqfgyS+D5h5
gB5cXWDTaAVcrgDMRoxVxzJEGj+SinWzH+RwwcFOx/1qt2zMxMq451MyRpg6eMr1
lVJgDrbP/LZ83A2oofO+isviY4Jgr8cp/Oy4LqAHQwc1t+7fh4S4cSTWH/pGcIAq
tUN8Dq+eZtHHwSIAXLJ7zRBF9Loon19iQVpuj8kolAe/5k7d2C4xmfB277rpDBPt
EXhLQxoQKvRMGAD8uDjO6aIguTDmFapFKFF9KJMPoX2zFZuJT62LsJvVwhsNCGnP
CJP2TCBmyIf1eQhIQUaHlr/aHHojaaeKgmOVCdQP5eA3F/trOnoItxBiP0xJn1ol
FhvMlySpMkGMmDlfNGQCyxEANpzUgZ296gbGP9guhq+oDDBnivBna1549Jcul/xW
0YW6pwZqKDDUyOGNVVsCONcymiMCF8lPZ35nTer760E3gB/yJ5vc0HUhMLw2rgJE
hOgjD+rKHr76rwJSSzcDzFxF0qTYxnOD3YNUjakPaF0lo5r0DxoC+GTrq1lxJicQ
BcMirOxmQRbHYzyL+lrOoM1TOv8mTd5dZJPlBUryYJ4Di/VdLXGH7R2uucSXoIhh
gajf4xHgPwAEpcair4sxR6YGOo+8myCIsWQiudLTnLSWYSBb+4VzkKpi53oXLIIU
5I9oR1NEYGHpXKVWBTpE0iRSjpa4vptLYCkdHx1sXLCv6OIXtX1/ptPpHWx1/M9K
EiD828bubTKM+IIHB+fA3I0YT+X9a7f236jnqv3fXLd7k60JvpHdxMl7NbkE05qE
8lSHdZGSNLKyqLjvDk8pGXdImQaZ1gL5d3ioj/SYeGf9fB/utBTDCzq3OYCltaWP
sWJdB0pKym4lskQWXjgNr+9ppmCVHkOMMb43qx7Uc4Tu4tUkWYq1oKTCBGzdQpPZ
qLPTPxuLRdl9gJ4BTYFKh7TGVRmwefsNk2CICVf7flzkia2CVylipcSG66ypQFdw
znHYVF4x3Iuoz8rpt/75yf3evALU3mnqkONJfvg+KdTlnlEhVnq6qJ+gS+yzmvAy
WctWs4e99E4bEyoqBzWAVpZUbXxpPnrZRGOuDHnO1dqYE8cgGKO2MTbvF2mBkxHr
cXfCWDZzhEUg7oITocWQLTxTfrinSLEjzEEhQVGYQu0sKeYSmM0LQ210lFlyUvuN
VJyBdQsD9y7OZT9sbxX6Q4jeBJAsnjnNFC3I4NDlRrwFKL3qrpHipnRSR/6/uFx9
Vu7hkftgkDHMYnk1guiRKfWLShOkc+6UlkcZ0nJf5rF0Dj4qm5+0MsDaJ5TZ0Q+6
/0SPo/qSHJgmpcpsSBglgbzNCWjA0Z6ilUj6geyrJufXR/Ylnvpkpib7s8GGtpOk
+MG3F8ThTEIyR+MZNaH0gUXRnfWJvJXje3Cqh+BCpeojTG7f08gz8T6ETiHRV1WK
lb9xRZuGOdObMo16j046Ig36OHUdCwH3JhxmPq4MCNzKQYVquhFXfWelq197hHz4
2Zoj6Ln5srFNzwFr/7L1Ok5Qkq8zrPfZEFLl5wnYo6LT4hqXuzzVZbpey9UnAISb
wu3CHioBKEY4sUl5dJWiMynKU2iboC3RH4WId4pzUICiMPG5DPVk29YyUACfDW3g
khU1MsOVKMUeNQcVxKcKk+1HTAAG9VgtR1ogr5zP7j8uLoGsT3KWA39itD0Slbv2
blP3mAqVdkDph9yfGo6hjImX5mUz4MeZ1UlvkHmnhWRHHLOeXl5dLtBRbD0Wx/Fu
ZP/boVjyli5pBWmDzXaUVKX5ervEhPlQh96yjOOYm+/vrjN8ftSgqDmAMVibhr6P
208q/G9TTexrfSk/NezQ74iG6HjA/dEo7dFXo0oA+GYXn2sdvJufrZH2zBfgXq7f
1h9pHV7Kc7q0LwAkkxrcBsKxfWgUCsskFIwyBi5DQDV934rgGkYsiy6JX+88PD4b
QkRQXoD+zS/oUS3ywGYGO785c5wsvuQOni9L/8vNdf1shzSQQWx8vaK69o9wQJVb
MHBVeGkXaRkgfvtnlsDiQQgcmmYeGSDIG55IvtORUJNhyBqi+XLVM896SgmZj+5+
eLIOzGkK1E0TjI38jPmP6JHQ/ojJKR/KTIFTWrc1nrOizO8RMFpWf8U/cV3RvV+q
t+A5n/3znjsXgc6ru8wUvLKGiOZvjRpmgkZjy4LBWYu997DUwXkc6u/u1XMoKlzt
ONzEE7JZ/qvVTIx+QXr+3nICjv0gKQGVTvNWpLFXnNIpw2fvw/Oqsrb7qW1LVaXM
9LMqfp7BwKg/rbYJuX6Ny3ZAsC/ldGZhqrQCNcNZ2SWOynh6a5mqQ1cMUDtVyUk4
95Os3+5tp1QSqDZvO5dmcTP16/JvP/x0PuVVBwWXfWj4ODmDoq7g3BJWl/SyrV7R
UYpJJH/FhjbM0TqsYANua11LB2L1Cg2+/AIAo7p2uO4genF86xr8th2KZEII/48P
j0oXKCgjQ/mx+N/wE5S/bocP8xWaMk4vQAoZAMvmF3Q53RzW7fXLZRr/ZlCXJ3kJ
QBrCmh1vxFnEOFm404Evz/4OZoiReIgByc6vx1nTXbBCBzVLVYFnXDmmIyuusY/a
kVmezMWkVPgZXaHYRkGtmC8vj+bcs6u4achqtD1EbMySa2fMmexukQ0ht+qS2Dd1
ZF0TCQ5bzWiAgCYvhM85XBstZ6p3SIEpgz9mT+7vXE+2Eix3zaxrTeFwQlKEWbLR
RcAwljkvIn6bPFsJ/9+dRTTM9XLNRevhb5iCAXtfmUSdECvpawPqDanmdWOFFPW5
wabFv1DYwxjmgnt+76fvoxmg/re69Xe1BfAtLg1YAWWFfAjY37fpint5Khg93iUG
abwdF03gFOsnuS9f6h6LWTekf0r4i6NAqpPiEdSsozN3KGUlccCfxdJbmkWaJdUb
zPnUOcsBTY0kQ5fDANSJzgHo578KOx8/T3ao0ysQIWXI6W+noCN2xt73WqvxYcYg
T3obyCElFyFN2wGq1fNt6MfHG63mN5K52iu3T60/yCroL5tw4FHoc3a54G5RyJB0
HgksK6shlam8gIAokpG0jLdFcbX7eLK4h8LDn5xAsi1o1kzRzIpS6w/MFwI0Fwbi
dUPKLqYpnR0zG6MmYyvIGbVzhEQfAyUWC/OPYMAfjfC0L7Q/jRnB0DZPkAvNW3r4
gYZO3RCQ+GopqXsCPPRYjgqvQUtHUTV2vWM4jieLmh4++eQuQLdeHqDo/xsEgZjw
9S+cPMPCILF6n2npRTJYXZTJGLyw3cAE55UE1LxWnan+awUuua5o/pE4kMCoSO1y
L7EEmIcy6mfvVq+oV7PJGg9meFOBluD3mxTD2xmANn7qs6KLptPEmHoPN2erpKKh
cUDmHlgGbik9SlmZ5oEFj9kYKcEvADwbIOqbVmOU9M54wImqNWkjEtWXIvSxFP4d
08PjynAPrGUm4IblewcItrOjcuxYnSatkQAQoJZ/c4twopwu+N+OURCUemKX7gx7
sQyBU9y3JKBP09qDB3uKE3h65MqFerSUbPmgBvko33cYP0kKVzHlMvw9CzyvMwzg
1aXaJv+SHIJqCc/ailaYbq14Sl0RFbz/b9ZVwwrIkSGZD8b/g8iIHQSFVdOJIoov
6JIMvmLvLLxlfMksDxGcMwxfTJIAnPHRSU1msDwAGPXt5aoMDl1HNYg3hwHifo5O
lf9jfaAs1QyTFKpInVGu8j10VwcTIA3xtH7nDvmL4mADZ3TInkzRGSxJhDqL8qPW
k1Csddg+GaxUKmc4kKOIp/t/cygWNHEw6OLHOr0FFsPas3GjTCZyjPRm17J47q36
kp15SV496d8QD1RqkmT+9gb9eqOIyk4RtHxHSor+5E3gk08DIHS23IKvPuCRaZMT
UHHPTdp0Vhyw7alk76CJd+i/P51WtNNIH5rv2VB9u2cDzfqihxMFTxq2NLi4652k
lv0emhTBT4v5QQg65vSV+f3yZzLI+Jk0FeuOnkKN0GkSaab5ZqwgE2y5voXan8du
tPgl8zrLN/7lWWgWOAv3Y8fnOWr0wgjIk4hDq+UuCu/AIr6W1MBnxQTBCdgFszbU
ERRVpYTBC5ztJ2szgQtXVpkbhxVjNnlsWefiAiYnxzNyuxA8fdUoUIZPd1kqL3cw
G0JHlVtg0WERbdTwTVt30+HboZ9Q4GXARU5YSm7yXd/MOHyKTT03VNBVekSvskoq
ePRWFCM5k0J48NAIcURuE3AcpWSkiBid7lSdzisKAfZXwKXrCS8tTbq1I33YPnuP
w+CdiYfeWbys4Gc1cURKXuYYzM3MoCOanYc8XYSaZ6QfJrnGy4hWp54LptwDOnf3
I09jd43hOUYk2OUMS44S5ZbOf+qESHylPWACbc+/ZawJZ1bnV3S2nhQVE/7PqkCz
vSF+3ksqvwODSVSnIV/PqEdr5D5at7phnQoE0Wj95OkJTo+HIWWFet42NxEnuvgT
Jy8RZ+wRjErMl6u+k8vf8VOvV8mRHFxJ0pG71A6lx/4pRcMv9Xr1NNmM0adc/HNE
GatXQfmh69GopSPAEjYPQDF5lw8w1RRTy4xVxuJ3f5F5KDa8uLrjDxqnn45k2LAg
hdMGL3bwAmFJvbbnWLTqdQlO9/rZ6EDc08eu+gvqNxzyNiwuRaSklohLE2ZSRf4Q
OtiHqk0D5y4rhDTbcoW9BFC6zasTU6i2Hq5WsLV/ZVKeoc4n5el7kVRBo3m0oMCw
tL7xz/+u2C36VeNEEGQuGSvoluvviK2O7YfYwtZfyA8u92xGWRhmLWP+5ZeWw1U8
ZMuEFQ4fyQFqwB75I+uCL919XsnlateDwOkBVAZgSashA65gxSXwL5tC+7KojdZJ
gbjbF6YtTuiVU9/d3s3Ik8jpRP/djZOzn8H7F3kdoGFZ19T82jR2d3l+DIG7SiX0
kOGBpKMLXpFCDSQRZaQxaYWuajE9sfxMwciHtcJqCfxRUuRrZ+YA3MQtxE0Aqk/e
NOBaxjfxifpoCpQQ6wGZhlXEFU4SVaoQbuQ5m3YMRe3HzpmeUOA2VfRbrPcH8oaQ
OGi1IoMAybSW2ZX25voMRGgjtQnKrAiOUMftE65n78OuZkfYjxbFPYlaGkp6XRxB
sKxoqI97FipBmNF/TfpH6NMBIMXYekx0NWFK81c4LBynF2dqTurtGthexuNhnFpK
fyY9rGkWTRDGauZHmfMQvbpmS1jL4hHcGCH4/8V0VeDr/SoCSqLmrn8D/v4vXFsH
FkBIhU9fgX5R1PAMDWv0AzNTDyIS/rKwpxLp8SEwcc3Iovhtv+LUvCXJ1PxTwxZ5
z3jlAzBsAMueX3g1BhsAsTxCXKaqH4b12D20DRnALKf4zXtLvhjPZnMqcpw6opev
+wgh/jY3TOIal1S/WGsc4q2+qW3fVWQhCNh0VDP3PhQM3/H7CttieJMo++DZeoDG
r6l20A0RmZny8PnCTQcA+YrbCC0Lkv9kVu373pcmyZFUOELKfSHoy2OmZCSRhky/
OKHPXFP3jOf8KwCAzerfPAAn5StisEIjAJZoaMdm7TYy5YDlBYmBsrouHFNuR6uD
Hfsxky8P2k61CXMwoYXEz2xAsZbGE+gJrgkQYopUR1qYh7fIDmIo61Y2pmy/+piI
CpAUHmflQECCTf/Qdm0bFQ/DC4WLaNtM6eIkAKugRSBil8UxLFKLNBNO8p9ltFZD
SHnH8Ow1jqE4guG+jzyKXkZKEpYRJAHkgIPc9o38RuHiS8y2+IQxnm/lXRct3WrM
5deo+pHIuJn7nKNwYiGWmPpxfh2Xsus/ibo/bKHiQFbObYJnmzBbQvWkxuv93qJY
fY/gbw1pcYjbzsCJ4iVy/EmNrILsz79T2QZn0c7RnKZEZrby6sEAFR3Ga5qiFPN9
peMU4I5POKbcZe5xMQ+98JN3j8tm7SOcvgGp3Uqv5iwyVjxPOEyl1jfcYo/nV6OY
hBEO4nIrK3WXpRek5/1vWPEJKj/bWKB9PoQUpUNXYNlRPMWhkhRRFa4hnj17on00
tDgo8rXrSqxoe8v9MoYCl96mAo/Rk4WDq5LlTqG9My2fLuYIGeQ97bP0bc7NecUk
2NsXWJECtm8FaezQQCyWWUpfmfnBE1G+C+/DbiBnGdH+I4o/LuXoReUPZWgao+oq
NuumlZQJg59/Xvlo/5eWXsqg+/zQSXIehTyoYrsjnW439wWjx54CuLhyGoMgDTXU
7sB+O8RMWbO8a9Yl45WQsHkd2R10Kd7HKK1p+yBDI2nj+qriuIAhSFSMjZ0Pucw+
4h1E7cPw/9DE+UHQ9pyGe1qW2EIU1ZVpay6ok3fMbJh8Pv1zhjKArqXT4YFWtBCK
sp48fVuii2JR/+I9D0vQL+cHSXL/3fwbk/XNeq9plRDyL8ytk9rx2m8TJcca9H9l
EPf/y1Dlx81H5RrJUaEwUsgXorpDiUieMyTtz7t6BHfnEBlwC9n2+pT2bNuu6eoW
Gz3VAZcQVEgTWkCfcajr3flv2oRVT0NoF2pzxzk+xzBQcEFDC5xsMX/l3Qlzfpdm
HK1j8QPIVc+mfZ4GGdx+jIWBV/GqkQAul++icnVHKiVEXmu4cV9Nm11yGixzGoWx
J1K14lQi0JhVkRoc/c1qWYVlvEBrUaPDE+yGoDtwP02xMEywTbx2a/NSRqg7UmNV
YGszAc3x450Pl2hrjWLWKJCu3TtoTYN/d+8Ii+g+ISwzCwA0zsfnHx/JQ6gFtWr6
zkDXFQdsVtc5RxjbpZSPnNnvhIEOvBzBBYxygTu8tojsT5PuKzsB3nu2YHOKHVPO
W5AEZrHm0xFCJeNZ23ps9njB5T4Wl5pYsarB1DkaPLESRpEucP4MfsBVZQjvDGqJ
0ePEYx4MPs/fvK/bKB7U0Ewube3qq6uqXP6Qu02B5iXIwwwCeQVpTSp039cuDBPC
CXguRTbxJt2vELzzubAxrafTIVyjIC/lDNYBVCYH3xbxU2mLoOVMuwcdhQoUP5zA
ro/vRWt8wKYQYm6Z3pzpVMCIVMsGJPAoJIpdxCtDHkRW4TSqO3h5mtyy6A+BZKhI
PVBXXxBDRlibnGWVeYk07eecMoXVrMPNNp7QzlXCv8pGZJEa3FfENwtLP7WLh+qb
ZwaeDuOdltfErH2uzKFpzhStIMDhuHCvIdoGatOKKAtt4jU4Fx2mxR4Z3yNanncf
0nV5aHFZGDbKRTNLr5Ddz8FuuMfqwXQpk5pzsQ3OU6+8D9I4rreUtWODQck8l7lC
esGBndQa6Kmh2Va58urMy8RmkC0Y+nEZ4Oagw/Nln96SPLhyNxuYcsO+s6APd8qL
pH0LZ61H4xrrBLTXthJrp+XjZQjIZF/VJW8bVKp4pInrT8vVDyXVzqB+3s5FJkUO
LxYhlLKgnDAGxKrmNdWqEmV9HcV/HdA7y1Bphzjw3Z++BtvdLZF08GCTBHDYz1Yr
wlYxxTi5D6KT8lzYu1zqaC5NayFZDNUt62Fak3x+qz+I98CHYaVab0Z/l1k+O1GA
/n3r2c0+jZlrPRPOcyflnKfDwfVDJu5AhurfptG0zVWQWZnwuKokNS8bRFBqHEYq
LE0+niNDsmhSYemiJ3dohK9iIUVCWYwynMP5XV/UGpoaKiSAYMDgaxh9nEqWrmVa
TmlP9cq7AhVyDm8zKgO5WcopX8NoKA3cbmFTd74E26K8mNDEwpNX8r4WVKsdYGDe
ePihubVDVSHQAl+qgn8pNDcEP8+36hjjWRlM0tYxwfA+K61O6jaQsOK+/nocE4M5
kuEHGLX7qt4GtSrLzETDFpuLvh4UcO9idij75sEYPty9qHzkEfsVp/0B+fxIQvTg
abGjf0t7qtwv07+6bqPAaeVsA08EBLYM700Cz1u3bBA3PA/aBDZsGRKTKl2w4dGg
fuYJEumw8yZfmnisVmqPYIcJtStpVPX5wqOtOtbyOV5TvvKtOxXa4fJs5Y96gzsd
u0m+lSnYeW4TWodGo+2XfCsNzJdFH8VZkSdkUOQaq1tjOcPV0gTBryXg+fxwgWq2
gRajUGuVtHZ25vCePwY2erurOTioe3KRZ/IcXVm26ktPd4MZpeB1nUJY2Q96sHFU
2fuRo3gsshuAi5VFvBp4n5GzIrYhGgbW0jaHZPwKO9y1GpQlDDIS7PL8yEFvmxoX
4w4zqzqUBpP5ECan+g45thFWgUA7peqFVxnLwntGxW7lpQvKk6kv7LiMJJUs3B4F
PqxWCOBnhVduCzLDuEuMkWweRU6Xn1rT/avno2JY+kvql6pRI8PuX94ZNUJ1tppR
J+2O7IHJxS959UZ85SB+ZQHok7H3McrYUUJcZb67CxfIa0npSDt5vy78OTbqij4r
kI11ThygezkCWLyXbuy0ZXMI4VCB9xBz5ovemX6BOYfD69g0/zcdgHYPyy25y1Su
5klm7+B8WZAkSx8u759xKaiWe7ZjMTAJm2tbOle9jz4sql6fbVbQtkZGd66e9Gy+
Rqfrpd2DDhJZcvJjI3bzNtffGR8hUJenmZBhgk2UkmBgyIIT83dFXLAEUz3Yzjbc
KLDtR3XLa4JHkHUYuRyU+YBQneduS2zvIjFDXPA5XEqydrJFPxhB8WsIqEbu51Z3
xOE8kyzddTMif+44l5LgQ9WAchf7FzXEm74uv3/nJWXkv4IMDMqt+1/ZoateT351
UWX+ydX/KqZkuh/FgRrDfSh7e+9cBdiHYiLFSnIjajbNUw2qUibdkxnuzGTh1qHQ
R0Ch6+TWdhEA/LGnqOTzQ1ngfE2H3AGQFbjzDS1FmFPKVIdbxrvwsbKNP5eqt3Gz
/5LphxJTLQCZ8Dw612b5GXwnX/HxWLAFAuLA/AhIVaJgGUp6jW+V94m71dAgyvpJ
SmBt8DaFyRiJwiMk2dmpNvT7hr/J3x6nc0V0Mja9SgByWC1ygRmr6+wln4NRUL42
qG1eR4cQR+9Yg8UW3r712eyIvQve5VBNL/kDZ7HGaNz+6hzMq/BXyRifSheJ8rnN
0CAklCD3slCff+HBbGIwghUYMA+9tzSeUDtRcMwehYLngE1X3h8FvPnhRJS693Zp
+71C5eqxOYbR9mUOtvTKyU6JLig5MDlQbJ3vuPpG1Bj7C3H6/3IShaLhipr5AjVq
bEsR2NCgaMgHmY67K+8gC5qefrtTzA23m60e5elAu/qgz+a+KJ1Y5bJvLxraXRR0
QD3h6VzCs0Z8A3dSQ3m/42ljVraGQH8SvJI1RyXyjIga2Wo9JpSxHzPDrAcXeDmu
4gweoyB+cCHKASZuMtjyV002caSEWyXQca1EfqcAuKM9ymkI20iqC9d4maoMD0TF
CukA9TJ/o19cHWgTAu9KGh6FADBB8iOonRjAihSX+qECng62J3GtHuJo/ptTKZJh
tkLcgRT66wmtdAcEo/gckBIt2kEQBYj94JqfIws4ddIsPcOpDSpJ9k8T56mKBlEw
mmRTEABmPiRbZSQKZTuQj9h0TVNGXq2WV2r2kC1njYqv+QcbKDMVeMLbhqjqkb7d
QOtBvIP2U+KWNbk5S1v16mmTY2lOWOFiPFo4IT7HuH1aQ9ojPAFWaZr01cPO8BuA
gqRKU06keXWeLYFBSAgjT382qWuMHS4KwWfGEGvnSVw6qBMOhT36ar25k6cGQAq3
d8fY6mrFTnsUOmb8r6xfzMuBB8bhWnhlSKdtSV5PIEkaHrzkRD8j7YNxn16SW1Zs
IQ9giVuMn1f4MgSwe4kwSltg+SYo/jiSKQet0EWKVd4iZjLwn/7HP4LdlUmmuvuK
p4IerjHPMCBIP38szmefuKcK9tT8IfO3tou7w1/ItxoDyEwJ2iMRBEdu74fGaUUx
Acrg9CP0LvwAiiohXNGK2WQLxiMgKQOKRF2HaeUm9LsHYFBAB3+naUXZJvrv2/Wd
MgJT6M1+kd52BKPVIXDkGVnpNnuD0vy69FRjl8icVknb+32WdfOM501UPGqKrmcy
LlVl4c+cQlRrqzbffM8V1xDSOifahf55yA5VUcKK15CkNzqR4ALFtYEeeB3vkXdx
kIoD4CxvXw/dzm+oKB47qpD4lkTMNe/3e7jLuzTre98U3FWbHFRLAufQOVZjuCX9
a4rKJKkKkwsUSiI15pcmhg9sEoek6h5xSn8igIdV6glo74v8RbXJX3JrbM77z2nq
hw3z5hjklOoxKHF0TQ5unEWqHXGAzSWFG/7iy30RVj7uLE1Nu8dN7yUkXne73wom
ESKAP5s6PHyOUBVLMKoyX0mMPO27GnB0d9Zv0t04y+lfgaAlrt7pUsxkM1XAlExT
IOSQJB5zj4BcE3wKLvBUeKCLIoXOO4DLG8/ymDXkQbKZW5X8m8wWUfabJKYOtn6y
zX0KfuuMiyP1qQgFywxDUOgjdB5gI9IPQJhBv3VUrQXfVrF0rK7DJgfkVf75UWPl
PF/4hnieA2CioA0eyZiKVmVpJoAmhxnJI7ZLbju9nY4UblNVg60+fIhP7SdFLRC8
Qt8vN0tRA7JOOdgwoRLdazkHjg45F5T8jMdVSruD1n80hffptm7wPKIqROhkp2LV
VV9Nszgh4yISqaK/kOuQiAkNg4JVpNaiP2BwiPUdb/vNrXf+gwaW1tdudEGpBlN3
rvwBiAZaouVjoChh3Y56/COlS2diHNqSt/iiYazucNE0fqIxkAo68XCNRKxmfsLz
1f/uPRFsIviQ+/dv+/avVowrzaS4DhRMZdcuNmG785y2NZabKg58FPN1JXUBFuUx
YHAiYRQ2nl6UzNhzVQEfTnyMt9Dl0y5v5JQV80nPJYwSr4+Ci5XAX0EKdZdhjBiZ
divs6DTascJuydPaLpY9OPSEQ1zwkKcjE/7lEj+BdOJqv7ADb+apNpauoMlB978Q
bZ1GXWkgORNw4rl2MV+ph2XhDI/iavA+iCWyHjJzi/Z1kr9t+0ysJDiVAxXWIETY
S1s2rFOBc02UlJj9nslYUcd7bXzxAxA4p/rqW7R6eaFJmKhZFnj5+wy4cHS8Lp2a
Zcti3ykNwsZo4641H2m7UEkB1dEDNci/8GtXTIB5mZak8DON/OLH8FT3JVFlWzsR
oNua1AjsVh9MeSyrACsIzWjrcgDKGuBH9+ufnSIWDz3xsiDKWfi4kASFkWFTZ1Oh
xW6/2fTMT1UaJlXDY31FwjktXmnqGzfmHNn41C7LkxrVMT5QDr8tf2K4zd8/RUE6
s3w12p2ILBjbicXglRNoQtS8gEEUUTGvXdfkZMw8jEFXf2uZ0DJhIhML0LLoa8wo
WVRsJBwq8aMl7NHwrWl8nNg3RJ+4yoYPvw1ZgUKpO23yIFTJoF0RgvX5xHTKzZ83
vGMVUgJ52xf4vKqK89JPZhInKW4lePiiin2w28Fug1+Ji49h31K4tCIanjcR0zp0
mLzK34XlJCT2X10HHehZqgQcjMGu6yYPYlFM0kZDhP8mcTKZy+9fbNoKzUy9gAJI
78h4k/F8LKAqKwlLJ7c2mEIrx7Q2Xi9RNGflIUyJvbU0Lpk2HGCY45dj2BVsif7Y
tbBPcMao3psTxi92EI1uB32sU2qhubaTJE1VQCo+Pge4IyFBXt9tjPrrh7lZ6q6p
4HmIOKHXa2QBLZunCQlRZiJ1sx7IWwd94zmR2dBs5rn1kuT6kJwK9ckJEMQbsCD3
6KvcWSGs1MxLptWf+p9jFFj1PEoO6YSYEKRZc7oJ+O6Gr7jo+/ZFMJ0M+S8ARsKw
IXE29iKiLFheFhOmX5y6eWGsnjccGsphdvSnRy6YNYIqkJWhYkNZ6/we9GTG7AWJ
qtV/cedHkPY+KnHT960MAH8Wt9sduOMMOOtml6SuFpNDQ0inBq1dGCMeJnK/Jiiv
ZATh1PeMBFksSWPaMk+dP5OoPdZwjtQB7P3lZgZbycVz6CzINqjHl7COs/YkJTPp
W+K1vB6HNjlpuN9j8dba+UB8JZNEUwS+KTYlcIjLCFvoHHv/yu5CvUlXlb6OR8gq
1Cc15gaWirWFYlx4AO/XONSzWQ/Fzda4XLjlBr6B7Td7Tt56W1IV2O4jDr3xtyH9
v77d5Q5sgC4tjJ1XewgmOX+xVRu2cK7d+WBSm8DQJFnYjbkA0+FnTRFxTwGSE4g7
eFIYx81Czgds3Lt+GL4dtYnWAeZ7NF/17VB/5A2fowCMOQrE3sLENj5VutEkKK1e
h/6Q99bO6Yfbr4oQ4aXqaMoRN5DicLCenzRnJ4iIN6njJ3TYK1aQKMzE1gLJv2Tl
An1drzzvll3lB13CV2btfL9HIuywTRbil+o53PI2wOkasnJ1QMJB5vIgiSKO9thz
WvMH/i9cYDfUOKdYgeKmJv354INiAGMK0sPw0o4AGqhbLC1bsE+UgU8Xdm9bR5PL
+8GB7cetaBcoZlvIxT5yTOYrOBItIt5dLGvfgvtS3i8mOfm6EESQ2pyPSzDpLIKS
bgufdtqr3jHs4g+UDxCS9kq1yPU/ZdTgst7JxE6Nv4PQdRtyZViBJiVXdqw3qD19
cQw0Gm3Z2okPU4DJhIOQFjSnK1v3vCBNhcEabD4Ycgrtji5sOGO+qLckOtTCbkk5
EuzXaC7itvH02nXIMJMkAiZ+jN7iub1Uc5O5o/Adgc1SU04lNGMqjBrxwPOOAli2
/5rz0XXuXukAG2CN8WMLjiEmLIc59SI+PjWiXeB20zHsoebeUtnlXhGilLs8RgMx
iTTk1b1ezuiZFYl1nWVGgRYJUR/yK6HhDtpL4PgRw08a0QKWnzrTMZHKhWNs+BZL
35t2/OKosUMv46KV1XOvAX/cKesLjMwH4ScvE3aXUzKVNGIiYFHKohmPy7w/mPnq
4ePRExR4iBau7zrWqovfYbwB2p+ZCkR4WbLj+u/m8wpFGntoLsez+uBfCB0nNZ5M
7HX5FGebsnSs//8/8Ugnh8+QMR83rEcyqE2cqL2en1YTKYhRzZCj89S81V8v5EtO
cYLmRrAPid+dtEvMbJFwLmb4RedPt1YjSkcfSQri67r12g9ZLHiIesVj6Lz6PKL6
SOu9F9e6d+7NkaADTRpdb6BfOjaI/xXkGAfpVSiiWUCa3HDqOSVg5QIOXNWYt3Cg
Y4Cph4vjDo5U5Y+VngKZaD/S51FS5A8hP5UdsWEvH5lS/f2+0Xr9pWC5rYOKYR3u
OC6Tw8ZOfau1TqXEdfgt/hBNWqFPDyMw+BkwmdWCDWSPg3M+5/SuZlRaOkfugf/H
13uyddrtbFWTP2sEJjJQw++RV5DlH/KK0yNODfhqgPglTVmLFiYKJN8wJ8IEaYgQ
GFBUtvVoBKkoc0X6V6RBQU5atKPOkJdnq5or05D8Iw3cMtN3KrJj5UrYVq/qnYrW
BBQM7V8DysHkX+kQusFCjTTpq0SXaEM4xQtrwzOaOb1uMnSZigTVFpXCKjCEqEeV
Yvl0RSUlJFCOEVekk8Ar3fuFczYuoFAR0265UpDaXTTYQd4Fpjc4I+hviXy7ePNv
hpHsgfuJkaoVcNWrz5jJm3C4ivTGgplZzY3aCs4FtMffcP8dI69QWEKbSPdRjkAp
G/M7vZbk85uklhmu1vY+PjTsLejlC3Wdr6+QG22WUxqV0LNS8UVqdM/boKuQRV3o
6jGeoj00bs4tVze5Icxcw1pxTr8Z1toM5lCFSTuOdDiuRgsPfhlOmak8D7GMf1Ra
nFTonpQDyWCIlnTZ5mXL3wvvfIDfGgZCLH0g7491NC9FKHSsNruPTBE7qF043Qnb
Gx8xIP9F3/gYF4Z8fpgkEOYzXdJX0Z6zu4SvnqCu/h7XANgomHdUsSgYbjJ/i9cC
dr5/f25p0xSC56muemOvBZvZ0xl8Cz8d2UilwrhLYlsuraDRYGVpFv+9rXU5MWc5
LFdBT1InR2Knik7kYpwiK/G1LRM52M316mshT3PRXO9KjNmKwA1hTIo4VZ9OPYZj
6vwfqxGCeymj2TMIMp3wvPinH4hKi1/HMnTtNqk6kXmWbq4VKDGPSYWXYhKc/mpc
rZqd+NaoStrUtrF7xB5cMoO1pR0VGIfQ8UPudmVy6wyLL7RI0scgXYcm2daUMAcw
F1xhBOI36pnsJFR1xYB9+CrvrSE0WH1CL5cSl97KU5knfrZEJwneODNMnhdJ1q/j
oG9FPlKzpGoZXFasYW5zyKQzzenRIvigE5zm+0jhOs27dsJ5cfVR/sWb5iTMTypa
eWmrXaYd670iqfY96qsbT23JS3NFf6WQsywRewr2Nyi1ivncG7vSsMZoZM0EBhvD
TQiLsMxkxtqg8825VQOS3/70uPByqSlr3LSVaZzzXvETnAlGEcEkVzpGH+AWuBDG
ZcDjFir3U1o5SJZ1+/tF+Ez2wOMu/pLpMDlRjoOLxnMN1lCwhJV66iliS7LcZom5
iSGeSvuYx3hAntVMHxZPJtCk22BE3h3GpGoY6vDqs4bUITY9R6sWrBAz6K3je1FX
dpL0gJXMwHk7UmtTXlk1mFXqZDbNb0NB5Hyg+3Y6SXsxNzxH3dXNgCJ08DtgK07F
TTQ7rxoswVN1P1UDXFgFgVtD8YN9Mn7C7AgHT+JLIQjAA3fn4BX3jaqnkTBeUOmb
4FgJuDzfpugqUFCrOW8RoRmkTT0XAWNEqJ1zxzOfz0x052FFaNAp0kuTDMXrfXvA
mbip0Bc2RJkiUVRFW0m0Vq+Fz8ZQCa5TvmfYCNZIKQMymwdv3ij1P93UwGZ0y1qA
X0erLGD3FWET19DxsbZRnD6T/xylzakgoHL2433xI1Xx62jcDWS5S9stjODa4X3I
WzL43pZ3oS6DW+lR1ceQhiWG/bGo4Af+6UWfwCU2HIhK8vT42CsbkZ4359Ubrz71
2MvPQErIrhEo+98/uoTRhVI94gfCCcZwdUdeQqlKs4KU6pqm9K05N5ekXpIVs+om
wEJkqigZ2kuNPSlxDOqQuDFr7qtqUBoZx00Pghf6z6Xw8ahDJxjDGxEwHg43ohva
KuvXQLPpnLMmRsNPAXV0kb/o+nxjLjrALg32xCoOmCUPGTwhWfdUqd3/qO0uiT0q
u/iLnJlsKpMriX1CNFniVVBAY5RyhVkVvSjDqZR8697qI/bf6uKExO9Qd4AVPRrE
svHIv7GVIA2/Fqw4hbMOR9QbnqRQXw8lfP+uvwS1LYjBdLnNR11US76Bb3LbFyLw
lS0mPdRAJubDFtndCZv6yCoH3pBTpRnBpvom/CAiZDkxoqRtfqsy6reLEzHXBup6
/Ll91zaJzMHC5oilXXYwOY5F3y6NBBQo2+tqcSGlVeTdsh5myrxlpAjmvVB2Utcy
KnQp4eJWnx1JokNUKssqzIA67AzMijt32ora9h57xmAqWqUd9MERkf4gLvrjgsAY
5egNzqE6rPp7fnOhpcXZod74Max2Gi2p2bSg4gzO31t5LdxVxhJI4Vjx6ribKQ6s
St3ddBepOJuFxbuYzBFKOEOoKDamNYh5z0/lkkFVV38/X4EYfGhFHUHc4C2+VQNa
GaH2MHIhrd3fY5TtKA6m0NX4Tn+18dESWfN6lcYj9+Z71s8vMILC/UDBJ3JGd9Fz
bFEnReHi7XMtftGQOqqJpdWhlAy8jpLlhxcrgCOexI7rbBiS8JRrC6r1HtELzR9C
ffywR02vKSgCFoGnhwc3SmlTOqbuRfggddLOkTsap6pagFY6Em4JhMpHaeEyaB9x
x4aN9vQ7IUlmFq303UgRo2SSB/KYGGMOGIv1SR5iE+X+ocjFi/S5hEOOYeg4z+vF
cl8tOQp32IaOdswo1ZsXMFW2Wc/StEH8tOpvpds9q41AqUGuACtPTtyDbs+0wqCZ
z+cRx07SQCmGTszRZZ7zKgqSb6NbkXvzmL/s2abGALQvrwSw1dsWs49iLKMf8C4u
5MOj8rO31+AcZUPSEiWbgnusKoA3Is7iXptcWaVX/AOJr0CB6TIXJqH4yGAJyMAe
kvYtIguR1lu4enY58eErjRPDvKiVsgt7LCGNfZUEjOeacvUGjer2e+yI7Gt4GbNa
GVF/uZTbkcA3j4LZiRWPPDRPvf0St30laaWp3ChTF8a7lVZLNY2Z5HtJcpCKMtCT
Ea9b65lY7xzplNw6pVD9xdD+QxFrW/C19bk1T+00USMeF45TzseyOHlS+zOvTBIv
RAx4EJ1KCLHaYQRKknA32wBmqFx6AuVTh8itwHU/AYC32j/rz/e/YdJFsfbSLf9B
+UqrbfhruPw0ptGYLFHTvkJPo297HxqBu06Txekut9EVmdetlLPr4CH7GWCigxkH
8J1sl97d4xoEu5VkTe37Q6oik+nM6pwSsAdPEmfsLi2hnB6+S2eVRvNssM6VKqds
lI/JQ3aIGB4xExVyT4EdEuJLMk9qCgE4sSEQMgy3QbT3ajUtUMBQBFRUTe6vu44h
1YeieDTBx0TP2+xggd4jx+YN8bOpKy2TR6lXAyS2ds4IJdc51fHX9UT112sUIPmk
ERdrEmyLa3Prd5Sv49XWRY7a0uYKAa1cO7H0kQiRV0f2grDJfcmRwmn5y/XsZTKs
nOs9EBkOTv72cJUaeJjtQWlGc7PGRh2ehcer24OUu6dwn7Ak5RL2FnrAmP039zaK
yyY5OJIcYpYcSJPRk/CDezo+/vroumrkdVDVUBagwjrj9OKyHHux7OW5F/bXHgLU
NrM9kzfenQ9P6liok6OEVZDQTzTpDy1LqUhul628LXTpoVopYEEHNM2vfZOE0dW2
8NQCHR1A99X54JMK9lxjQHXpKykvpgWV5d5LSwe4cddsCqN/dfuLw3qKE/3l8ctF
uHyBRw06anYhLlrUjHk1ksCH/mlzvWiztPXJ5d1hzl5147Bzgzs/JHDxOwG2Yw4l
/0QQcxGi1ybzjC82txPz9UXaodJXNwCMo8aXle2irTGNg3XkXuN5nsW6YUDgJe0i
zq7Hjtcvd39po62eSDRNK42FjZldWyiaELE5vMWa5f72VTUZFwSSvgG6FrxvpLJO
NL9mIPgEyj3cIxyeHNqeT8UDxIuO55PSfkK1IgwpLm5TZy8NbinBBPeGb9FvT82y
rB4tAApoEnyp/fB2MQ2kyDmnpMFimikIQoL1WX1zPOgKDVXWDmlEakErmUQTgote
SzZjR2LmdROCnMp2eyKQb9cuQ5ajfGT88i5b3MYMYd0M6KP/iT4WRRvBRqc+lYsn
Kqq6NQSBmRy9zj9QIIuhf4PTbZLgaTbCu0EAhGTitxkRE06SqYVwBue7wtKQijtI
exMaeSQnW7zKEG03Xsky6eVJCKcbZamlqwtBdx3JUUgavRwnfJf6BNGriZZN1CAE
RQ8OC3l25rLHQ6+DPCF9wnlk0nMHRvzcASMwCNuyrm/dAYxwVKu1bXFz4BatoFZ1
dLmGkMFrNk30Jzljy9U/EIe3wENpVTVqg0uN2sGYDjKA+BrhGOy/tl8QMR1U4xSu
q3FdOOkn+M3jy9Xv8jw11CAmSzuxF1t+M3Ldu8EfPIak34wxZ8mbBbob9BuUiAtm
qLCyOg9a9gSYWfYbWLShP2SEPu7oKCp2NdSojKgMvD57fh7W6wNcBQTRjJ2kKd+M
8Sda4KgEgJGtqHNOtJbF51Gb//rZM7i0oYIuvQfxbKhTFb/3J8lRnUL/DL9otiZe
mFlr9FD0v98Rowa23eDtzZl3Y7G+v7rTUdAoL5PqRFO1SewTSdvBkTZjJx/Mwzdd
N9kGxhFKO3Btlvi/1mng/kJ6PuFXZBa8QiW8JBPcfKafnmonErwG9fzAnlGGFWsq
E8s1Ey7DBog/jc8+/VKE7LU69GxU2/Mgt3Xmo/MWs6JpctrtWBQ2xa2J8sazgSQj
p68Xz0JKzpfG6TI7yhTVm0SSxud+rzLYsl4a10sPAgGwkEhQBWpgODOwF72Rabco
MRmcDHeujRwtgiYGwVQ8FZjH72pPqhiLwVtvu89GUlIAyRltSKP/vLTp0xZuNzkG
XIFz+euua2nvnmwLCYcVrZp9KY++PMg3tVzUgq0mMSvf7ipJEbMBezdgYR6RtgWZ
zK2wteXGRRbuETFU1lXG8Pewaq9tMsDxaRe5UA+dpLUgnWX+CV9PDEI6wx4Cpiej
SKZ20OdztNG6/d7Way3ZX/kgaYCwPXykieetkOmb0uHqBLsop7UVcineVF/aNdRv
6xPuUW49CGI/TvmtU0jH6A8flVGQ2293sOsXvESLrYkiDwr6nL8YeM4tBvAYTklV
S+oOIZ1JBVXy2c56cITcJwkIgmzrid1zJ+LyUiBm19S14o4UoLUzMN9kEk2WmrJN
5HZ562gjhVk5+aNJWoF9yPI1oJfknPw/mDVRk5L4lc+Zv/ijjq6Ex7R6n7JMWMH+
WQB5p0sOE4nEVdrVsoTaJHL1VGSoxP4C8T8zbGmi4vEQde2y4h5nAv0WkzKyfN2k
j0AHRMt39HbebGzLjXlO466vjfeko//xytUmRX9SRZj0hKJxtySrD3hySfg6L6J1
WE62eU8y/+8c6y4YGTj0JfA6eqgEg+rF4e3zZQNj9LXU6VAd1Iiv17DS9rDsCj10
QM6W2m0PNvv8YNdGjbHdl0gq+gqVGBepiBwO2DRarg1a/qAXhILEdRbSf2jcDYg5
Q03JJJGr50V0Iq41DKycFclXu6zhNkh4Xdgm/wLFABgfFNnFR6R1AtbCB/LeEwZd
gBAXpKC6AazUftve+a75RzsOeA37RB+huv7tOMoQjqQORNvl64ibErUjepBtQrub
tPGVsF8hU8q1gMWggajwt82VD7/pMn/zzzeRM9CipbS5UuISTRO3XW0yNyvIBr6N
Jx4932msZzndNObypXFUZUbU6H7YS5NWRoXXTHSN+/mciRJxC6Dz1YzVVIwzMsfQ
nvIJh2Q6b46oKpSFXo4MdyguNfA+xNkJ+wCtB2U28okQ8B/MRmiftpam25cv+LRh
xXXNPjDuZqoOpB3o+AnXYj/VYadXQeNT8qNgVE02VMd2hsPHRrzVb7QFh70COOJH
W4FzXLr0BqaW288NYW39XrhfXSKUsS7Zvho0KFGjcMBjXkMkgDt/Y/FQEzY9tWSY
LGKHYf5P8MA3JqtFgzWbZ3AvQV5vZmYDB86JNI9WbiVI7lnsjSI8OvuIK+QTklzN
iaClzrNzyeXwEGLowGHpxUMWMqR9pWASRCNzVdyq/usNxZeGOloRIKm657gh0CPm
kL6fWuwid1P4PnjEWOCYbyfmaMltVJhvjrXhcYN1/9ce39Ub4BfNNLwOOuKWETEz
QVuX7KL+6/KNik6CrOSlbHmFn2LeFE7EkcSJCVQc84jttwYNhQXGAtmBXKSSY3r4
5QRhFhahcD+8S5d0VryHgt9Cuy6NE7rXpPRrxpfSuAuYznGanv/J4tMBG4tF61Wh
CD3ZeVZLYsZUzhepcGACCV68MhgDZi4Eze6s8Iz+C1YcnRlW9DHTrG6IzRfz8509
fSfBFkYtFjXzBI1TAaGdMo/CoWm0D7ryQfGhy9Xqkc2xK0og1lkkiZoZeKF7FRbK
eU91X0NiPKgLpdSJuKgRyWaq59BQ32ZuZcuV8iDXkOHSAteag9tt1hLXxSCwtLyW
jXQPA/MEYXkq+uw8XRBYBnSuKRl9FwpVzs1Xfiez2SfShfyqlyewDs4GSDwrM5ub
f/ZlzD7gMIZXL23kMJRQ4gWcLbkMXQJs+NWi0ixpojpT/0LShVz2hQ5R6HjzdJPy
Efo1ZhJWEMqyNOlzZrY0gSMt77TjGxBKwKvusDo+r+VxmJhlwXFM8+Jeygx8NpCW
iSMfHHo1yUxg+0s8X0Z0gpEB9zw/GAsaXU2FuHBtAV5dTTAfIp/ilAwMqR0twtk3
U706RftgH02n5Q411EpAaC8B0BuNkmtMKUK84fftoXXCPG6unOnOYUQtfwtrZQuA
IIX+2NYL+0KSD7Egn4NzgurSCWkK3mHvVx4ztbdMlh35MmzxdEcL2DEAJ0Y2pCQF
i1i3oIx0oSNgX6HoBOnoR2RxfKIxoAGeEkwjnJhbW03gJyImc+7WjI+uRR1QPdc4
r6oC1HQR33VxCnGbveP7SWSV1BQUYe9PC2NvATyw188YY0epgy5I3UT0yQOCzc89
WPYO+1zU7dSyuRiR+6k9egoH8zoG3bK7zpjZa1s+ax9XvTjGT4yMVn+y4vmWQZY2
M7NY+eMsnTbRU9kifgneC4zY0oPLJJCbZ5tPpmSgeTlNnVP1jfxoPJCZi9bF0gtQ
hnOPy5xTZKlN0P5mqpSrmLQNkCqwOKDfFlv4UYRipIUUpqlcy2oqrqZzejdxML1c
v+ZuhETpa1EBdpQBZiBFSPnXRetTJieGZ5CwzTHRIEvAnM53N7Kgs8r+Tmvhv4Y5
V+BAA8Tvaeaw9UaScS7EJgZTUYmSAy5jlZAILNXC5hJdw6/9vdVEq59fjv6AMo9h
9r2rulsaGr2PGJ3bSfcmIc1c0hhg7vYXxMlHzVMhgF6w2/ChLvOuEGPWj5lGnV4o
Ii49r7owfZwOnk87pZQvFQmQIT4isIbcQVvNk04Uw3VldNWKcXu3lMAe9AbR+ZY1
7cOISe1qvQZZevJ6KtOoPP24FVOMYUdnSogfy4RExd5JxE4l1VmNH9U5Aqr7HIW3
gJV/brAf6fk4boN9VUCVAp9c4PevIjwf9C9RrfbfNcV9bCIn/N3mTe4YAyiqDXVU
VaQ0+LLbmKd5X1/UqfTThAEFy8YrIkTYBvzqvYLqJMrc8BA8Tirv26AhezDTldnA
W1eoDBNjOC6G3aIqD1OOm0xiL5RcS2Y/mM8ZdqoI2AMXALBlVWK0hjSHlH2tDK9N
ZQO42lixa47lPNz12445/G4oqE9CNk0Gv8pbstWYoDWd1F0Bdusw8q/xI8Aa0tAb
ptLuS20Gkphcvwr4eZPKNA7+DHdYjWj3TSSthPh9TrhqNjqq12nR9QzM3Azzg4dw
LxjtQHoG6rsLLj44g+MU1zqfyjODyeZO/tbf/XlP4acDkq9gN6tvn/w3pO31sD0o
dnxa89AeH11xnmRYfCm78GDKmKSyTON7HpQDTx51eVCYGLHU17ioCfr9IACpHbMP
pjxnJo1MCS0/o4L2aEdFgv8op0xg4Z3XdLnnnvVPrT2ReNE7tH3418faIQCyEfQz
YC3orXVNOHcxkQgJz3a+JcVI7YY2QGGZsyoazCeUBlpvaZR7nPnknU38ca0CO+Ow
WmIjnFz38gHZq6OwglTJElj3mwITx/CMFVWRI+lbRrw1YAX6FVsQKpZWGvWmVjZ3
Xp8xL3jdKRhqxdGPcn1gi1HS8KsI7B5u7UfaH/bZaqiugS6OW4TMVvd6GgpkqZVo
T9d2ZEi8j30as8Pt0KoMWRy6VndLQTwKzDi7/ClaGndw2R8EQlyexqQ9UK+HMWGo
jhZUvhJatp+1w4SCyK77u7ZsQGen6Mh5JuExfO3bS6K9anEV1nJuUiJw9EAQv1+s
xQEY4oqzZUJfOw+zKLJRC6uD67lXrTE8mMMpUC+BcEccuxxI+jTMrjaYMiqt3Bc1
W0P25O93yTlV/SZ9XvrsRKmMAE9o37UXdbeChWhKDi/ceFqpkW+SKUc4r7AdpGf0
NJSizx/dEfR4DiOJKsHs64aOqKuY5Kd3lTocWUpKwTY/tIUDLsHlq3EAMxGHa4dL
AbUPRR31P9E0T1cHm7RU1pLiZZQEvAzY6fWoAYV0ZfOBeM7nCjpHw1BF2KfrxdbF
lf3gbLD/azCjQvu3iPTOkiP4+Ludnti28Ki7kQkLCvwjSR+K5VdCDLJ+dQa6RJc6
0XCDJvIm0UaONSVuN4Ok5kF0GVGhW0dHzJ+MJZXsWx+CjrPtfiNzsglasFWl9SZs
ba6hOHp4h475rG/pDL9XxrZes1jwGcMJKd/zm0LfRtT8w0Cp42744FeYwCWmr/0g
Ev4lYXZKD4a6Z2sIZLvPszH6U/EYeB0wNOXU2yN16OcDIe3Ei4FKSq71tJ9QFbfC
1f8hVfWmenWcwWu7imwVuua0xOdPcY6s2WaxRDENjyyeEkSWYP3sbL8ItvuWjC2j
wZ3E6vkPdy6JKC1Uh2AXjMf2pFdNCkTKkHKnAKqgTBMHgdxvWPUBGVi9FVl9O8CR
Ofn8KfUslfXs9zaO8RbtrzfgIlOFA3YuKC85NgP1wXvJHtwTNdg8fW+a70pSNDG7
kftt+vU1O0bYaJkuu/aTlTBXnGF5XJjv+SrSg+GK+fGGy81Xg16+PRBAUwJpNy+L
pDBkKJXPGF+RQUc/t2Lqfv350FpzuqRx/90LlafAgygJFiE9Iu5ftJMhyWIGodKl
bvmi4aMIqxmQXjf5xo80wCOtYgmXAd0sjqTkK1lWkvDERfp97VM8PU7sSVs8uSt7
7bnsVPTumcr1jNU7H4H58IM0ZT6Y/dTSCWGdqicxUHtsaoRx8bLrz4kS7P7momHb
Skcubn8Rz3NRor/cH0VHL7hBPW2dw9FV9aIh3CciPCZwPHMbJ8DYWNN9XvM00Ihy
X8+HfdeBKPDJfE0kYXAq3XZsQZVtlAtVGBY5tS8cEAPD4oKJucPG1Lu1cyk+NhXy
wSViLU1AmtOVi9j+1q0vktgTvDqVuv5MnkWt1IHD3VFd5U1jec4B+GhECQtKwP73
sFOrarwLhLu1u6budFrCKY4Zo5pm9HY58WRYXtD1h+xfBnou3pM3s042cVrEku0h
7LiJz6LiMgiuSyrQFOScfFEymTzehRJaCFf/of1aMfcpYn9uSrIZO389vVQNiKIT
xOdOjD6PdQ+3CCzJA3QKCaSQOXhHkxQ9zFajMPP10tQCwqPLoHcac81Qnl5fukb4
0pglQMUKlrZmoibIPue3XFCFRdK5wB1sTqulLtlNIrLW1UcNHf6Y7zHyVhAakjIg
dk46pO1i5hhnLrBb18EUb2FjzVDD/07MGmKGdU87EuADMY4GQNEZUjrYS3jk0G6t
0PoQU6mJow3Lg3GnvDxG78q0eOo+NGZCitoE4qP+/a5tU6M1vqNOgM7KxiyLJ3mv
LKl8fwNnlUzdKVgwvNDgF4pUxQl13BtWggzDvRSXVbtpIPBuuSdxxRXOrdqT4uad
uNpVSC4UTAtiTwM4RWPBvC/FTdJyEoTFHHEQed0Xiwemceo8JTjn+vkl/qAxXPTQ
Gy+z4kTuRUSCzqX4et3BC9Slyl2ctF/lJpmEhd+j/MNs7Rr7iAp1cpaHdVqEXmkd
gifwRXRa3N1oAwpII/YENRJudT4sAkms2mVPYvwbn30bYOTZc2LuAU6lb1wjIPFH
s5aTDq7SxjKAkBpvwbbdhSDl2K3ihrCIWv5OVGt3wx/TU9Pafs+clLck+1tqvn3+
D85N8cdVExDYfpMc2c+W19fLaZ9uSI1W2nl1cEYovzK7Q7zBwrfr+O+ps+f4uJ9m
VgEHON5nlzb9jJqmj3v6VpnLvG+rojiciM51UiHvQXKm56mR7WoRrxeebeQ6U075
wOVsa+BeCm4VwHi3Yb/7QBxxe4c0CENE+h4Fdxr9S9Oev5aTK2SniAoMzvNiPOot
Ao6w+2QRfnX2CW7jVL7mepeh0M7djnbK3JU0DOducvugfnBWjwBOzBc0IV5+fX6K
Lstj2ELLDXsqZ32pdavj1a1Gkd2jkgdinobh2tWj5PYEuPK/7dK2Y+MbfmKN3muG
iV6UM3gKDmq581LMEslqRYnU83yVMAaK4nrc9qjbhzyl1dRm7fivRQZAc1jQcGPn
IiNgJYKTtwE+oUlqDfN9Tuaz0PO39UJ8dnbobIphTudhMO2tdrmHGM25Q84O8Cgd
2DI1Bpg3JvnkcoU3WDdqGATp0F4TWoNQPmA6P1xmqHSk7YZj2kn6cNV4AvhQF+yb
bDcMVwjrksmSQO2lapxQSRjEz3f4DfAFdmItgt20hxPV00y94B9mf9/uXJCwFiv1
GSlO4VPDj9SwtUrserx4LqN8AjR00P1FLnRSKdbdhfwtS/pR1GW/8qPtNK9Ee3KO
qskywn8EZOpE5yjjdU+ou//pNTKx6J/A7v46jiSdPyGoK3FW6oqvx4ySgkKrZopg
SsaNpW+QXNVrntyEVxxpPCl9GM5Jtu1b88fKvWVR7WgKdU+xxky1pmwOf60QLO7F
E6H3LeGd8D4yDvUi9KDMoDkt8wLAsh1enjTVTg0CBLApq+sttu2SJFrOHxKTKx9B
zsO+jG1NPBl1UKafiAIHLxm+NyrcdaprmQ/urf/gegyiTTjaERVIKsk2naCyXooe
JcdzBXjIfK48fsNM2Bm++79gPy8foI/Jwfzb6WT9cOUs6bZTntbYAUAoEiWSGnVB
w+oVKyAohbLIX5wE7fHN+TfQ0b5yJx24uGE/Tqjv0lj+TEzxXhu8EItMZTtuxGaB
47F+VMuHkiKu94yKIWPWkCkYB1s6ydYVFBL8Mfndlii3AEs9OhJ199mhZ6QL75to
XfnM+q6CqB/iwxvHyVOmE7IoR8R9/39PCXokf0/Ix7SRTH7M5M7vUK4IeCHh5DZE
aqolD2hi7I9lmIWgARaeNw9nf+v+hcWXBSnAVoXtYO19AYkVaMQy7ZWPZ0f8lke4
eq1mUupUyw3eudhyDdNjiw3hfgRwJzUtqYCgz9gVjl/lJaMtul1MrgW7pHSt68Nk
9GpZdiPG5XXVghhFohc4C5ODuZrn/quOkv6XmaJowObbQfOrtQ5IDEECNukBq0sH
tEUMHM9rKOpPjLtCMzaAkMaP8RQ2m6J7DLm51D+KZQXlwZlovWeysKIDHR5QtNtQ
edKdJMZ/KUWUrfKyNi99lsRkVa0GyVucFS4NdvgFs03YEZKTVldNOR5UsHmLdsev
yLwr5rqKkqCQbjtvRUinhLzO8Sn0cljJVBuE44GsrqaMs1SYKEq/fM3iuBi9E3Co
p0Womrbh24e6DvqamyMZQZ3hR6xojkf8w0vFzaEv8DjpjL6lTcoY5g3voexvF29J
mivEfaz3XGAmT/Pjgxe93yPOPqwwQqzNK1Io8Q6bYPn88WN3F7S+IS2mOzXVh/eM
mkfPT0/4/ujzLIc1Mx8HMxR8fOrG02OykXaARls0yCNynOK5NvK08SEeHKCkWKoG
nO5v6iQtM3ZQd3dRKp58l2uBUwfFYbx2f6+J5bTtEh3PA5xSaD9zHgYQqstykkhT
XgVeUA0kk1WXDj0VGP5o+9R/lmJOTCbrW2bDSYf5jNxbairMOInOMykJcqHeX6DH
pLAs1NqoSQOqG5LbVQApbcPXDCYinaqeGCt6SVjrDLbG3/oAg27ied4HUtqDZ2Yh
7avur/YlZA6+DQ2yoVxvipSYGGqodXsUH+H0J11+qRW9Z4c3gnuLEc8+NrF21BQw
efgzwFZe15+7+MgD/806sqmlMPIL4/d3VH0Dxt9bKaJFUWZPa3ZDqjycU3U7+ewc
ecqHYI2LSnfa94Xd03/FwDNBAiPAGPXCTzE4dicNsBRymrUYLzcLMPqxSoM4z8eG
DarEKSAL1x8AFGyz4SS6UKP2yW1RB4OZ8xaCfwOCC45TFxWoTZDvPVfBX1ELuNgy
ZQ87HQGA7r4pJFBVPw5Y86y0Dljp+SPYNxKQqPjHN/4x67rF1tLm+nQLGY7fcCzo
3kl+03Y7Q6pwxoyAAAg4qRKt+1Of+b8gWNETkS52gq1SA+DbriTOPzLMSgArK8Tm
wZ+4gL5plQ2o9VvRUAxcwFTe7GvqiHGh0db1v4v5Fo0rXINhHRiRLe4ZxMpATdvC
aZu8JV36xkRnTAtd/w04gMk0X5FT+gxPjJJ6V1rGDuxkLhKzuakVnQBR/DJGoU2Y
wV4C1tTX3D6QjCs2nInYXSskhpMZKi/MW7fIv5CBPtqMHMA90CZOoNxceGaRJaLP
qI3oh4qfSus8PytWEgqdckbYtm/QPLf29RfR/jrVeev3v3R8Pa1BdpUE76xaK2Vf
zujH0jyYBioCzl1nq79PGJFvd6eeXiSZHIH51crQN+RmnNudWmdBIq26RM8An7Gv
S5vQaxLShxuq32BORz6BAey2Schz1L96oIRmjdBO6EsEeMdc0kkj6oyvjx2W2Cgr
qFPZQfQDrDfvRnHMo2UJ5TEt1WeM25FHWlkFtUgfXRaa4mm/Cnkpr8s2tw981dWQ
DRbuxtWo1iv3CNdGf6BDuhw0yjPGIv14dmjusbLVupKgGNkA5KV9w8k3RQgFx0qM
dJCF3JRyOS+sVSzji9MMtFTFgu54dOJ91KcjHBovUbkBV+z+NKRu3LzwGAVfHVZL
kkBNr9mAML09+Um+rS9PeuHHpTjrI0r+f+eVt++0Yge6kd/r3QN047NjHaNJibg1
hf6cN13Zao4RE4BsjvOyBqqhTZLP5RYzHCiW9ZQdS5lAJFMsXbWMufz/njifIHXZ
Fz+lxd/wBPpFxMl55sAQRA47xTxWkHYqbU6EjzS4OAnd8SI+ExUjD7EeJW62uPEM
AG+U3K0MQYUISMmBk97l1Iuff9/m1S5Ogz5EHCyzDqsyguYUPyNZRHQ/aVBvc3ZQ
cYdZuFlntTOC7vdRD3F9qbzi85g92q1mvT8CmoKBVrxX5oteTETQ3tY+voW6IpbF
D2MixxK/AIuQiSDRAz+yif0rRjFPUS9h/VQkR5mrdqwcWkC3j0b/gLqoGpl+1oAy
2ypEeKBrYHzlWdnFZOWcMdeab7edRfYv+jGxnXGyAT76XD5XLbad7/xR70O9vzRI
iOhCvrp+4/KFiTWjVLQkhXhsWBOOhtTRXcpogi7V5oMGVJ4toprypt9RZdEfuKHJ
4eHDR4QYbngR1xELI02eVGLa8+g7SZzjEGHEeMdacrsHSkJEPPT6GkL6b8IBBTWV
zScvu2kDbCXRyBYRtTx9+pNbiAOhvRRO1QxpoSCjEuy/ajJula/kcqnKznYPZ2RU
KBB4Kfdw10ja7v/GU+uAZyzbPM3p28X7ZCNzPu5cVB2SgSTkcBux/frAXQPdTMJi
U9eCi+yUPBit6QjGr8n78UFIH0tghoUwCSDHV90a3pkTd+Vjuna6b1QAe8UDjrTL
6tOiqCHKQDTb4ArQAlSHKz/zT+yzJpavNACizBec8qpLYvdTYeSL0O60ZKfLm08N
2MY030CPAX4eRMhk3ry4Ic2KSM3eNbSBRglK30RRdfGllXe/NkH7yNrEwMln186x
OB2dCXN/zL4M0WZoT1InQA1SSeoKZjKN3HRevCYNTh8Xx0X4zybV1zHzGqJcKe7e
P75+QvIqQ1QMXlphXfe7n09PAEPwPJFN/eKecNj2s7UOLawN9tz0nTJNcE6On+q9
GFr7QexHBHHb3HzcW8sVO1xeVsx3cYkJAIAXjYiIPdHdnAv4m82YX61xGeuDQMcP
5IMsbUwvMIhwiKo24VZx5j2LQFnilmVOD26Lr2VUWw6MLDmLi+ZAYJ6Hw1uxHY9o
+EXEMzlplaABYV/Pnhis0Sck3/wBx5WXfE9YS+JsyWhUELmbQN40ZIs+bwxCH0rU
JsGiWIVcerwC/PwBgMyk6la0jx6V6SRZ+9dfAgZ92qtm+Oid2S7hZtvA+O16A+mQ
wvDaEdfx3ZM7cMBdm48aSVaULQYuUJ4lSNaUIOFyZQvY5LlbHKriUKfaWriRRhdc
Z4VVXWFg31kYU1Fyg82hEpi3VnlZQtXwvbpFcUlZeqjm7RF1+Py7BSp1oUwHu5GN
7FrhvAKPMa0OuSSkCihfE2lW+xXdjpQ+AlQVaOoO9YO/+HRNGGJ4i6buRF31+Eky
45DngjsqqFLI04rH29pBX2CsLIpMoG8uuDi9mNvNVsAqBCfZQ98cUNyM+6xw7yIn
Bbd65Y/vHrMuH0bMz+fLMoWay+zDrkpFcGpqPCmNagrTrak/ad+NKKjTk5rjm//Y
t9GTmRlowr8iWFut/buF+dToyDtzl+MCiyk7wv0akLO9yjMyWOH31l2zioGbI0QX
C4m/hTra4rnX3gMAFwZJX6Rpc+xiDIyxaJcAh2bK/NfZudImd773eXdVBA1p0JV1
8XCumPap6EoEVHGkGAAC95olj+CB1cmzKi60eoELL6fx2Fhb31RVRINYU4M07G76
3QP9qclW/EmXyhl3OuZ9mLYW97NLNkfsX1VJoHjvVnTl7ZEf1RrwEja6oSQHUnq2
gu99k7kC1UoehMrAxzzE6fsrYjL00uBu4Xxe59WaF8mnk4X7EG+Jcswh2o431Bwv
yjuSFi14WP9JG8fXg/yAXTCF2jA/d+6Fuvp/78r7xtev/Fx1mma5vC6lTLOuIg3Z
swsaQrhDP3X8cwJEtqGOp80LtzhATHNUADLM678e9phNJ4zLwqY6c8gnL8BIc/Ew
QPr6pqV9dgP3e9E15pI7EzIqi4E5xteLajo9Tg1Ha9D2Pg4pMCf4In1c7ExwbMm/
yIMYMrtYTdB12eTn2bWPqaLSOxjbWkbi1S+F+E6NrETr6Ue3gVJBjWs4J1iekcpC
F8Oe8vKZNw9fTT8QXMr1DCIME6mnuux16G3UUfSokzgbNvToWK4ArIVuR15xR48c
prpB7SSEDNM7Tw0xkwhzEDhE8fVL165NtvuzVsaGyhxqoasqCM0uKlRXayhrIHIm
0DsOpe1BFZ9ILTRCh0V6bmfahg8LLNPke5jEBHq85YdDnXdHSzDCHwJh9fY8xOsc
0FxLpjg/Be6BbD7Fxss1HpGsh7jv6w7COIbky30rKPAu1yFAaYPMA6rFwdhTdRtP
B6RLC2cTMajKfYnyCujTcoexO3CDcmamW6Q55rQT6oFSQhbczD2h4aiYTnX3VtiJ
Jx9HhNbQ8TNTFwbneLNDaKh172lUDlqxmL1XtZvzCad6qeJmyd5P7fldpGWnSt10
FeB2rcGjSz0ed8gTM5b7d3BMnRZJ1rZV3Pkbj4XwVgQK7bADvoWQnKyIt1XJtsJz
QM1JwSrsK0wZq8qv9Ec1quHZWcR7ZsFOtobMdvRvVF9iOmyaHLd30/KcWQuG0x7G
BtQ8NeVe6e6ejkvqGRqA/mW8VoyM6bfl6VEq8aE7M/wjW6uOKfvoB3P9RTHAR5rH
ibtJ1V/KMVWG3y7NqWdjfo8RRTP/8Fd2QsX0BSdMxVdKwxJ5WBu3AYtTZBXcp1HL
ajo2fuVOGaL6ZlmwstsNfYOlHCiPW9OjtGTAckQ/mAoa0yq6UAaYLlqUVBSgPvKD
NMHZmyjQJWLM4efcA637aYkORzNPOIaGV8EkDDYLBMO3FqeAlxtdD1U/mxEoDTns
uRVxrY76S0iGeYY47f9mzvlVBdNSm3ocaffOedlG+pTxEDI5g1QL211cATB14H0O
fDnXEO92dJ9LeJAduS4Nx3+POS2ryA2QAIJ6rF+QwjzL5Q8bi3LE8yAO9zehBny6
hldR3heMlWNvuXJfxyhExuMNuCz5pxUSoRE2V8+BTEsnYxBDQHYbR5UvzXjf7SOV
mgXGbntX8ZESQa4C74018F1RDOGbOzWdMnTJ3VFN39zh+9AfdeXUTSukyRXl6GZ9
LAf2rehFBQJzWtcbFJ1S3W43qA2fRyTiTLvWNbJSin2rAoG5YzrYHcyph1P07Lja
A3uf3y9KqraLl56W55hBvOQONnBdh5vfHXO5hwrR9341XaKE0QuAMNZBvE96HSIP
0WPASTeNNQhs5vNNKpnpDE4yxdsol2W+KHbWdvFsNBOu7GI61EPxCICI8pmblovo
ft/Oj40F6dkYcL09VfX8bbWLkK6ScxrygAy06yqpZdLGpT5iwks7Oq9THcvqdx4V
DIdHLVe1MPOHmlnDyaqwsLAksIkcF5YC8dZNLFbeA5fSM7PW7zj3jiFkH6aS/7PR
28QPi5ZoIQVNJAnABOvqFBow4tn+hUZzKq/AtdV+440bSXesBCbRkeBaAbMX1ABu
Ytayck+PkdxvK7fdluXZyo2DODaWNH8Fo1ZTx/YXUvcdtPxUnIal3VJxp9TFImwj
1Lk4pvP89XV3LJEMoIN7vvXNwONA/LaRSvcT68IgJXcVBgmGW47aMkDJZmSfZ5Wa
qZoZjSyfaWBWSHu7hDc8Ucpcf14ja/n9qBR1fQWx065diccc0QjHql7KD2JbmI65
LAzytEjihnOhENFbhp/7a3mafZNYMZ2PpqMOBfSfLu6LNheCVEEBkKQt2cSS8Hmt
6oHhw+0CsXlwfOit5kXSdiNVzgEx3RMiPuyFfliD30y5Yvj1oNjQWUY/jF/tjtsB
cHow0Yq5SZqy487SUj6c0HWH7cSb50aoMF1JiwtoCK3QOJ/4lOetkevxeLR3Inxh
65VbV6qk+zRQCNAxUpUFQtN4XEyzLI09bKHbHvmA1auAm4BkFr19G5x51wUdRLC/
yh7csO3W9AKCwleX5gq0/X5bc/vQ+myrQkmkkZm1y70e6fu2eo4EFOpHwCs1L2qR
tUt2deSC95WFMWW09m+9XNoivmFCuhc2ifJfRSe1lrVui8f4twK1yNus50of0+B9
K887bb7rmRd+hl3mwZ6ZVscAaYy+uPNHr9AXFkMSyEf1fiYlmV3XjNFVw6pD/pok
9mXOIrV7I/eNRsa2XJkGP+OTunTsTMGCah9Y9cl3jUVUyXF7ZFKJuT6QHs/6wsPJ
Ia6PQ96/OzbN2Ie+kiJlrl+dKXUuWjjGZkEQrGU1YfgEqH0HZzPQPiv9cAYVGfPO
tRZ8KD5c2RoLG8jADHbMbydab0PBbsieD39K6g4rwZ7gybXZRXWiw5ejg/oC7vAD
USU8XGUsMiJHLnJ6psd0nbQ4firHTc6azdjeePboVUHowXdQHRYx0qt4TPYEVBHt
go3roTm7OWSkeDn8h829cIVlM3V62jgvsvEnjKLG81wMw+Asw8H/nqlwkbf2D27U
94FkC/268kcKLsX+q0i1Dy49AIyrMRRMzTruZFQIEewVQ8Vg+iLhZuQ7unDkRR4c
TFVH39PSU87Y1/2WH8yj1fOYqxya+E/agAV/soZKHmBGYKk84kZuHnn/jEs1EUs/
by/Bx7Tf5QDYSkAB/WYiSFlY3ZSGturq0gxtZcEtx7Wi5kTMRz0Zd9ZKLkoqwgom
0cMQXL8cq9xErLdIC/ApD7BgyD3vJF6ImFg58R3CRyugE+K9Vd96jAYYvdp/F8aM
WVLhdAkqApryqrrSBYZ6fTFzkrFbIEMVOUw8WG20jh7SdWaaYNJxq24ow4WB8bmn
Ck0q4mh7EB7TZlWMT2KfJ2S1PFdd+55mh8s2pvDmNCG/s8ySgDvpSK+QD0v2N/sy
xLSfAIbvLYA7hyZ4Ksr1OyADAuEHnrsCq+NstFkhVlGEUXYvUZaQHSXDBLsh1hwH
4B09NaNWHVZsDxrx6IVlh0KBCyH7z1yIFB+ZB7rLaXHNXSTZTFEZhstck3gqJbZH
XObzIYqXsKoyxXFHxIu7jGHzjzGGKwsK3OX4h9SyotmWv4aPgYHaNskhLVJMB1Q1
0sISVJwF0CHoJi3zbh+IXAIHewOfwh38pz/muXpHdnZwZ0sgjvWJ++8ofhg6DOZc
ArqumIrlCstACW0UIBkpSYgZVSGGf8PX6BBCNhvKgln+vhYomaVhikLWrjx/TQg9
Kpe5SQVmevIg08emRPLFUw3EzQ3tnT0NwtHisIex0MvBnzCPNubk98dg9tKf60n4
Ff95/RYf3vW//WqG2dYZ4g8kA3QKPJOpeKaM35s97F/Sq60NjuP1+kRfkHpiROdM
vqv/tFX8UuwOMVJcXWP96Rhd9ZgtLCxN6P5/34xOF9MxH6zGK1djrBwKMlHbuStf
iF48A6wyREBZXXI81sMou/DHyy2FWQF71WHwGidyY5NCNxdsp5I/Fed3djpxMLBy
iIC27e+IxjbzBcDwu/gqW6LJOnhBsSoi4rGkT5wt4tqPCpk2BG+1a69wPNqBj0Yw
v5u+CUZ92ncCQA3OJdgT6tW/C/rwVLBY9hT8AebGPITUROfs7XqVjhg79N2oR65U
ToC3gJTRPCqO0r+vDVSW3Ph/rm9y4RIwThfbZAtgfmLA8k4SLB3emiIr6narc9tE
3UB/5GdQoMDXgzS9yMH4QIrPq6CdZLAZhLiM7v0M9+sDF+Q+BTVrcfpBUBRaOx2f
o826RaqMkPBlaEkdWIyU3dCbAh4L2dDog8oyJdhpAzemZTdlZuSYY/ZWW+fF1o9F
Exd9tiVhd1oRvIXUlgwJJbGkggDs1Ex+zSVgjE4yC1TJnNhepnlR0lQx6mcfK5fT
7qwPW0fFOnIKBWiWwsosnsVWZXMKWNs+tGg89MstGcShKeW5vjkKp854tWuj5rn9
rzFn5vIKtKJgrKDDAbXFdn64DdndlDHyaXzlpnYPl4v+Cjn6FvIQeEH5e7ZSUHyz
CpgIJ+VgsqTxTBhW8o0wLHNVBrPoUiKddyn2eRtM1MTaQcW6lEke0Ue+vbodY4kC
Ehg4rBZCnNCnK5L6Btpe9CUKFcp7FFUYIaWuK9ESA4HxJxp4USf60T/6EzQb1L/m
Cw7yR62hxI5iobIMTIO7Ewvz6L1O/1EiWIFrSxfYMsExPDcLHensEuljESZn6JyP
tF5DLnqQzPTKl+DLlmifxbZyCuwgIIi7c1iotiW7LPtz8v9ZnJ7jCgSEjEZ8zdBu
3xEWSI9Or0A6Vto64xz/EET+jGatNf8KOqLsKoLBV5zuORGe9WnUrCQiI4hp+h0K
8A3V1XvbhvEuG1n73qKKkMO4Yamr0wtGFjQF8+ME81cxjYZdDw0m0+UeJf0E93sS
TOyZoJfaLLfneERkADa/TjV1SU6ylAdIVx1xNhPqnXoECfqttq/cNKzLk+Twj2rG
pzdljh5zyI1XONareiUzV3znLVfbZ//HcMJng7nqtih/EgGaSChlWKI1jEFB6wAg
dHnbj9/eGJeb3DHE/JBj7WuZV/LxnbL8Wq8HlwkMYGKtzBr5ly/z8dy8xNYp0MwM
nAjgn9BSuCNWKJRyGXdDgdIqEJWIGlvzTT/2cQh0kw2skJ9wr+U1tgq2ncW1Pa0i
wYY9jywfTReb8GkNdQUg3LinzmqcH0m3c6NP+ATOrrVNpr+JkbfHFG5CR/qALm0Y
Y2nukk/Y5LuE+kGIBF7BMCrRlQ/Ayf+N0nRpu6u+W7ND1BOAfenzL6AwMXf7KBiJ
1y2L+CKXJJZQ3uQSoyh+bPBbvDg3AWWSmunxREe6jVdfunMzLf5n2eONBOb9/ybA
9f+mCntFNnXd2HTv7jKmvbYM8W+71N1AJKoq6WjDmx8gg23wNk9AtPz2v3lwq4Pw
FS+sf2fjwtRok2wpfErApCrgqGP+QO5S2pk6pVnSXiFrWg8XquccbSTbslZfVDNr
OinJDiQ2Ezz9VcvnUWqlResjRNuAP6ZjHZoKZJ/RRKMBsZX8dv7X5TgacCGlEQaJ
evlhlkARr1hCqB7timfBMAv484ia2Bgig41iqVe7nrV315bjPpDQLoNEXT5JqQv0
yQEV65iZYeIShCLS800oCDm8/jfXcYBtFYkk/1l7Q/YEWWevawkKBtpKFNofI7KC
j43lev4AyDVI/GWG12jN8bzSws1J3kceuFCmRW+zWLXwqry3GIFqjO/pu4ATtUCa
cQSPtkEfzFlvYW2X5I6hZALcb44KLhIE6iKzRb40gKCovvEtCUWYgKgAaEAS9P5J
aUile1Mf1Pew4oww7ssxdd6ASDe9L6e4Pm/OR7dVzuErs9qTWn8t6ngEXhJrKYkM
KNscoyX1tWs9iYy6kdW33d9vnjaRv+lK9BeMXUoAPtKWJzRWpYVdB1nuQ2B3ps8z
SUF8zV2CkcE068PJFBvncWGCpIjay8G1wNjgA7M+yuU70gLf75MXZMwQ9KrTUKEx
WJXGSixrmZlhwiWm7Zro2KvSzDWyXUU1xHl2oshXZM42lSQs0u2lBSnbht4KgyTq
yZNOXHR4eqv4kJZmmUHVpwcdpD9wjU0GfsZ2Jb+1SziauKJtaulz/RvRh9Pcx4cu
x/K+d7CYjytqu0rB/kQ8dCNZIHx19xsQp7xRb+E1cGDfJeSz4+JNYfDhKFTrYHqM
yTors+sZuly8kzp9TNhHUg47Xi/7y9beYZhrfXut2Ps8CjoiPvzwPanqnEiM11Dg
vhWYhu7dbmSkkJM7n8qJKfzAWjdnUiIXWe2TkARbVzioMpKBkdGUrlJkYR1u7CXP
9gvUlba39pcVo6ap88cNfG+z6TKnddP3ZXnQ2xjGwuyMI1rtc0+SGRKmt/c3o1Th
z8nORBwl3cIFiZj4c3tWZ2QJY2xc9qIUZBJhHNCXVhzQvHM2SpiRGPQw1LAklH3V
l+0/eirj4S1aRWLQHydVrIFfBc1sMo7jSZOky6NY9VGf2HKRki7/lz3qufitNYQ6
pQADiVLqyyRJLZKOmWsmkPwwNCcCQnUEVpizKg75CoK4YcB2S1Lyr37Yzx5xxI99
TJj/waybNBGz6tmWenvK2ah824zxIBHCrBd22H9ytgbtLJ2Jsx3BqCZV8CW3KcjF
qDgOX1sE3KVYgX52BPcN7UUW9kw3yeudIENfKJzQRFUIWWnth16vsjBlNHY0of7X
CRIy5tuNBZoeDV5/lorhtX3lSNfeRLyDu88katSPy/FNiyU+j10TNptu/v87Q6ly
pBwyBi4ATiK10RILrNh0l1GajfPfUcgWdHh48qtzjf8ZWtKTMX3Cp8iBrl/MBSLH
ulbDIXHy9cB5n7SojXR9OYARQxC5X6r/2dmHWYrSPzYIS4n0GW3Xa3xwbQqEg2Vx
xQhtOyDqciAG6+Lmo2lnDn4hRz4ymGrqzLImXkHLp0QFof6P1j38APl90mxQqxm9
ZB/VEbiJ1o19FQwdkXWGMa/LcJakdFhhKZFhXopXiGZY+LfUqhrDmNOgz0jLI0s+
+Bbd4bNVMqHkp3rTFP6zajPSYubsw0oVealYvKjGZsuPNfHmNKpPmltNDJOUeTCY
ogandjTE75UdkDJchvGxPV8Lx9/9rRyzXhyD1fBXEPiHaTDL8fgVQcxDl2jSQAU+
o75ctJ14tNdVphLbI5cisaxRKYAR3ArfR+FM3MVlRRqjchDdTgJHU2Xzhbn8jBBH
N/PzMDNZuBxCKkBragbUuz5+i0241tbxtS8dJ8uBEBoSdzyQJwAjdhRIQYGfbLev
QP52SoISdKOLpT1ui269URVlSnuIbUQaN7wKyN8LWziVgFvviWrN4buCIb0J8A/9
iYb7Dg5UBjIp2ChnCSNWkQpw2+KGGyxeOwX7Pzej1CChu4NWep2gfLsOA244nxph
PGSZBOHLDAM8j3PUMfqqR4II9YTBPh+QuiArDGlX8ap4yPtXWsfSjw5F+hXpKPpi
Ao2MnPiQL3lwV4d4F8U7lAGHAdFvocyeLJnBKqsqplPkZtv0WtRoMs3GUAyG+8X1
6vYdPGAUUtkdfUFnV101DtZasyGHC/i6LmA5okbhUnk8zRlQlQLJmzy9kUwE7zcy
rvKHDu2505Y4r6jWSCtwXxvKtuEOXajqK1+HeGPJ9kHUZ5+zhHQtiZSY19Y2ySY5
BPpZTX4n4QIAfMRI3rNKJOw6D27ncR7eTvUOMcYAoLFIX3Vy2yVyD8rN0eHDDF44
f63mGPiwEGKRKwyRFHaMo88YMQf3a8Dcjv0uQpYVzzM35YJ41SfRYV9qa2tPV7Kg
yq7E2Zr+WpxWg3SuZ8BDkwskT/cLqATWkopt/VsjbdMwwJI+XmThcvbcBosgqdFa
CfK6wDOTTlyT/02+0DjQLEKmmixdiNtkmIKRs6+mj093+uw8zYlSL+8MBr26bYi3
hOEuTd2gU66ffZLaDERoGHdsPUhKELr1uuiPR8GeS0jlTwc8n2CNe105wcYRstwJ
1fl8bID9auzAQa12wUiwv5SbtOb7lp5HxMJqiZqu2pwr6ijtS2QxKTU5IbiKp3Hi
ZEwCLnW3sm6wsVdMq4TlcuAaNbXtKROf8n4zEE0KDKs8/rmM53J1tJetvJ4yH7PN
fJaQcOZGFo+QtVHZQ+FRXwMVWmI3CEIovGOyqTkiYPOenzavtP339IfdTjWtFYdw
mKS7mpCFzOVrmodmKhyDwazlOUq3NqKf/lwxnjsLCNviq0izD7v4Luxsq8Pkicn3
5USslu4KUEgaWkmMblMfu/MNtLL3c1CJdXUhnw9tJgpdC3lbo0uVisnytYfXk/H5
drYVBh6WXEDbVJg65ZUpgS9vaPU2MS7HvRL0b2Sx7onO3vgI/ECaOR71dLDKaujT
y8beFlFDzoxffDa2QBgK1Q+z8gZFlJRY6PlVnMQnZZ9QjI2Su74+lU+GtDDqZJp5
pu3/yCwattyx3w8/hte7WYW5ajtrDrdRz+xhwSs184BZgVLUzUmiHl4uyW9flEIY
tslE5qjT952F0OCTZzEvqvbq2eyGGeEEv5x1Q9XO2Id5EhwY6yH1rZjV08iTSOg+
0gKWc3cMiHZXtC2ToF+RByAlGJmFF3pJl99In5qs8wyFYZ8/onoGssO/lxRNZ9kf
Pik6dd9LdqIkGopJX5jjdoSLZwZxD6PHj9PzrYIe81Zkes2i6GZvOU9zWfw9BX2x
rzy+/+zCmDGmxQKZPKjl5y6f28Ns8hrbLz3/sKsHpCLGF2tZ3r+y5LZ265QThcaa
IqqVnccx8f3KkPMzPKmh2TpvsDl95wqxzg/+zgR2xvXnorTOF1MZbwH8rdiIOrT/
ibyTcam9D6qgKQRWVpVSOAEmOWsQZz5xp+ML1lT5o+iZQ1Rjk5XJXnU4numYQKAj
L0NN2VuhB+p+NnsZeDs3S44iR5e93eoNRhcSOmkOmqUCRGa5fBtAsDqS5tN4Rq4Z
3Y5JLK0cs5HzhNxmo2TgnTeEEGiZSRyvTjpyNNt06QlAvkQYZkSC19fPRzcfYwKA
WLXFwkPhiI1hsIXdklRFGnbmv2ntTC++zQItQ49Gnkp9gTCEzLA26AP6UJ8WyPSH
j93Tt/szHaWSbLiw73PPUDhCHx/2BjX3OYm7EwmEmXnC5V/AbaxyXL1b+LPsJCgF
fiRUcTg8S9ATA4hF2sAvE6ghSMkEzbuOxVr/c35oD77cFsEVZOkUl+Urtcx6XFvb
j4fTtAb59PR6osTmCJYUPM6Jgt0ZBTr/xJVEo9cMmA/jDvfsNmtQOCp/HGXR/bys
u8wQ1S3MONx5SwMWBa5vombw2/ZUc7s0y5Uy7pm8ID8t1v20gQb1IwLLVEs5OPPF
SDI33tRr58Y7XdVt/sfscP92HAKAUMETPHqz60Lpfnfr+AKe8t2EPacQUa2O08sR
2V2RsnBOM3u/x72G77LsAy3A+kce9Hf1adaYqhWuxiitfQ6ho/9vF6/m9Iin4KOw
zLw1PQvdbhjrzSYVjFDsHlo3NUAgN8v+POjNQxzKqFtJZ7yNdV9tfhWMMqNtGa8S
quoYUOuDGR9o4fRxdpnx4r15gxCznBEQbcn8A+Vh87PV7y6QgAvq2oOUIHQ59TsM
qKC5xPctF2rL7UiFVTSbdbn/rFw+KtNnt/eNeoUeXJ6TFbtthCX/D9anrFDq9Udb
Xh3/4c0LGvUkT+FOv/mJYVqe7mpPjoKD71DnVSlV29iyuxhHwO0DT+WIdYj/MBwY
IEpJHNHr7UZLPAjDRwaNd3rZO3GXIbuy74UK91YtTAgpy3nWxMcDSi6WAasWe/58
iK8FLXdoBJiil2V38bgEYAcI67lPfwoPJL/llwiJqvTwLwND3zWF9Gu3iTjIiXq0
/rMyaH9uQLHBtS/N5JS9XYzI+kltjO5El/kCmPtmrFGJPd9L0i4jsz8vvuLydBlC
0tfhpPyCkl/gzOvjOAu55jzg/dQL42wDZCdfWzlRIisl71rYQKkKlftjNHVpQsiV
T1cH84KRvgTI31OpCsCvdcuGmyQaKoOQUvwhWh2cXc087pCkJUutTjNOr+tPZN5m
NuoHbASrfD1ksYdYbxxdU+Roah6H1eZWRI0dW4SPMcTnoHdXSwgCnnwOoyBN1Iiz
OTsrxbLWa59rwkGUwIvxGVhKahyW9LLB+C6YIwD1Pb8OoIHOT80HsFAbJfrwLrTr
d9er3ZqO+zTnujXc9hlpBKVXWS5c72PRIpNqXXCY01LnI/2oJo/k/vZL4BbWI/zT
PGk5wgQoeKjWbtvkaDrmKk23wZDaYbyfBFvvVHdYCQN433d0IjQN9u7CF++0O3xa
VGRSM57t8Flrw/sql6T5bmqDvNc8UbOgB5whmaxslVnhI9i6EjEJ9hrpqyai+ju6
YBKszpLZ7NGTDwwIEIsykAh4CFYHIeGsOgpNdsIT4CYekAUvPUrGlVrBI2Q9sBWK
k4U+VF0xZteGkslGPpkIbsRA+Gk4SLuwH9wdHAhgauVr3x16ZDakBQ7/cxGUl5xr
bAiRxmtzZNhQJPbhjS3oY0OfU/1W36Z2HRfOWVN/xHNGdsmMXJ+qvYcTjUemvsas
HrnuFGMDq8i97DV6ChZuUH17C9sAF7I6Acwng+uUI+Czr/eLhMPhrmyMPPluhDno
jU2h3lyDZ+5jF7S5u/h2lBXWDoQJWre9gKG5kJ9jPii98LFDr0yOr4CDhDJYpZYg
1YfWPZGdPY1mL/53nk7SWzaGZEXeomPfXO8nResV14Xq7bNwTxQneuuntvY2G3ZH
yQYzU7pVS4/bSG37GS88mknZG5s9W0n7V0M4JO7xn4nEduKF5zZX/vDXg3ql+6Uq
oOG+A9GpAOl/bBWTdgZ49CCD2F8nqAjpQy9ctHNYdgNAWiqVzaFyroMSvyxNep7M
u2w/xzVkbTcJyEjvWvakndUeV00/En8sw4NDoC4HtgtyAvmxSg7kvtSpMuBrVU0n
fNIUAJkglX4MlJ3dgwoJtkxiiOVg82jfQjGZ1QmWA82MAr3PtbAl7tlz7OEIyZ5W
9xa1trtmsIIJkbVeLqkpmNBTuGQgP1VzJO5tiDPnMLu3eQcFYz3qXxrKF8N/66zv
Rte59XhK1GN5TMnVwv33O2GWcc5fPzQKpygDN6VF6s0vnxj0NK5+qhkb87eCxaAL
Dk/zmGlCJwhg50zlDkwoDvp4T0qIYkRQ88w9SAkodhJn53h1r42tUdQfYKAmCSUM
+v2RxmgvP4OsqIJVT3b5IydFiq0cIN7JPFrI8xscyAfCMxn5lMdvIA+gND8q+Q8N
LKxuN0zNg+uHqdlImRHs7X6O70AolOKwRzzjqLuklgtZwY6ujyiHzJe8Z6c+3uOD
v2ucZ1A/JnvzRPVjyPJ6k7SZQ5Z8D8LhBrjLHZZjB73qJIoiaBfdmVPs0ZjS213+
uC0kaiztGF336mjCld/UmHmgv1bTq7qjNKzcuPk4CZTThm33JIgcB8A+D0h4Wi2s
8FXh1GuDBpnwHEQmeVAVyNW8gIPjf4aInV2iuB5wzvOxtOk3TKarz2bhalQ6PGSN
ZRnPLMOfJcBOCLbkjZGCe4YWzQN9azhDO1xSHxNmnymu7BybwYSM0wNwWuGNCpO5
8rHb5nqDqNt7/bc10Lm6VOWbObt7CC+IpZWYfVJkHtGS9vd59cXBTMY1RFT3o/8K
VY59fhnPukRShXIeEUasvPaxt8LhumrLYPOiTCIu64DMRqkkI5o1G5IEryGxRZfG
J2qEFrf+2yUP3j4b+r/SCHZy6tDaNtQ0sfDErzK098Td8DpLxYuCJ/jbMOXv0Ijz
jEuqxLddDW0JI9ZMe4dY+4Ku6YQQisLNFM3Xvsm0stPw64aC6j331+mq2oJmNoQN
yewwGYzidH5/h7SF8NL/ZvgohoyF2H/5TTyRyJ4xDnCGqNi33E9Wks9tZKIWOknV
q25G1tFerUm67iRrFe+Pz0hV/wxpQAnSKVITmyQQI9Yw0Kdk2S25A4U5s2Oup9a8
XwkslHzVSGriRlzsG0KKmBiRrw0R4EG7zynGxm1tM3iUtGNQdi3pY0YtS7eqnatm
eD9Sox2TIcCLrYTKoMemXVRChmr6XWHKG3AUlfMoEQNYe/Qr4LkLlACxXAkVkf3X
ty5vK3tjx4DErHj17cE/rnhK1S7eYNx0a5ThoG+zZhXgvVhVDTCDgrfjFhxHJxeJ
eZZ8NT9gQU73iAj0Cqjph2nM0iBUKMoneg3ZBYa+YORTumqhLSAkih1PJQvyTCv4
PwiIHGDNXDjcKvrKyIUBZRFwrmjGVskhBahv6mAXbZrjMr+Xn8LhWw8iqtEMTGJZ
7JKWz+U9NAazlgCaX1ZA9L2yxo5coKh1iHuTmaPdDMxNSlLib78CZ0Nr4s9nuwq2
+WTOzol4R4TlwG65o0diMWyVoeO/rCkscet3pGQAjdECesw4VO636UGbXfPsPz06
YdSxKi6IX8+IGKm4znGIY8QM3ZsmHmAm7nnzOdsGMKZJlYlHEaVek4rGh0tlXzWx
bAxSEQRrfQuAqAfs66/DgwXC+2E0Yx3mdAZZ/Z3ETnbm1SkNLnJHeet+MGDlr2AT
LibJAVuPxRWk20lz8QE2PR05i+6BRwYzbgSK6nW1Cxm9k7WdfQDFzIbwg+jm1cWN
rnLe+ar1ILF0sgr5WPAwVmDYiu31v8kn8UDsfOsG7WIKMzNjsbBObZu6w5FQ3poe
3Bf1KIclCcC0JCvn37HmCobLhiR5CVa8JPQjzQohg4+Znku3eNzJVcddYxb2p1pF
plNmYBOnLXVBdNF4imQgwOqPOHzBl7jbRhk6avblm23QhhZwwCtKKxVhLTQM4HKw
iDr6FPlbFCcEAaRO+jESxvQHC7Y1fovv0NeXFsh+vFdb9fnA/DLzCOwiTkMu44qN
8oj1tpxe22Yz55J6BitExjLjJCk1AY8a7NT8dS5WUPQMxkyHhWwyD8jrl0Ucpydf
v8OhmemKhIJqbb2OaxhtPAvX2oPYKhI4YYA+28Y9HKi5jx3XTSvEAetMEvwsIcss
6ojKcDOOL5NYRuQyC75sn/iZGk/S51MTbytoH2bfMUHyWnAcJrhRxCjds+E3/pU4
qBKQrlB6Rrg+KGxegFw0irNLsT0K5JJuKZrjz6DYFmvqOjl8tbntZq5A9osmaN6+
/Vn4bac40YNIUCaJ1RDEqtprXgukNOzU/DBWpr1UdNLqu1Colg1m5L2bVlQyFEg/
VlUfralaTZwnpQINSSyXQsdjJJijLRd0A2jZ4RC1JzsnSzuaEQyyXTy+1zGeNknT
ky9o2V16wz2a0CVufxH4gPPwBW2UlTA8//6WHNjUFEF71LgJP99N/2tMGK6VwoEj
021FS39cQZOk1xUNdbZSr1YakaOtPkEX0hJv0BT957iv3idDun1IAkC4ZyTC9Ulx
eZglDvYJyUuqpJPTD8imGmloqc7YvcOwyZH2n1mfextW7zCKEgF9DtDBvDRfF9L/
fXYgzuq9e752sITaSacPykzOocftPbLLK8TyK9NbrUy/OWU6eT+jVRLkFBEAw7UY
y0LhK+QnDUMPRA5KKIA574RSi8I+gQZ5jpQYVbdrVFmbZScwxEHat84OGOOjCmcW
Nwd4ZZrMzSU9IUmcu+O0A4C1hIjQaiHypjvQN5tAiUvKPLw0VjvQCOcymoc5Dg1j
M1R0xXwmF7cLn3WtpvKiJiLcX1dJaquMJf9vSJtfjUZZ/H4OXy0lWo1GXeu/Xoqz
lrBQNn38TU0Pqkq+V9htC/CRkejniX5g7s5Ld9M5FNLEMgveBT6CpC9hN891ATR7
vQRH5KQlqkkeJAJOzGTDeWxgl8vb2Di739IZCK2lyvzcWCLrYncziP8to+tblGHG
cvBh/MvolzZknQjOmQ3BZoFKqVrJrjaYDz7Tdbw9BWe9xDm1t55JbdWw+WIQBx6N
LUb7uqtt40+4HyyY6wiAEwylsQXz+ftJVKrb03UV7aFqI8ehUzjx/G16RL8R29pd
45SawMF3af9aqIBt6uMlWTairajkbqEMSRDYKiwCBYt6Koa0V0JuPqKmbfmbteCa
DADxQK1as8yoFzip621+axTB0HEGjUPwgQ9eaoacb4SPIOqXr0zXib54f5amYx85
/JJ2KfLU6KQUkGt6SXD2CNnH2XHnVmd0MYvpJypFW0I1to2rz1MbQSOYJzVmrfZc
8Z0v1Sg9Hn7hTiECEwQsCey3EKgE3EECDf1rStXOkNf1hy3u+m/yGpbd0kDG+9gH
dhFxUDT4BGq0XVwRyJLY6a6HjyOZ74oAzGjwrQvsCV1QIVjFTuaD7bTysRjtEtUO
pv5sE8kMXIGd5fEttxdNzI7qQe1ULq5zVvFToK4hUmhNkbKM0iTAZF2vzesZ5/Ap
uyG/U4qtXIpOrHq3aAK0MeGqZ8gRDmRX/PyyRILhk3klKdmMtxIQwRCYQ00/5aJk
TPiWSBswX80cnRY69Lc6GmvnCzdktFTCREQTitFaCKxofnJTkx68hkZxM6wlywRK
aGt/Y0tQf54FFCfDhaH7UaoroargQj1ygkegFNM1ISY7VU6MKZc4XNimY4wcVjaM
gg+BJPdXN3S8CfgZPtggmI1V0w2/scgF1HtzctfAn0TjIO50eA5XHwtmeo8re+Yb
Fzwwnt7Q2LNEYlw4/IyUHsf+Mq7hDhWtkMfBrZvwcyvUr+o0eP90otG9z09oz7gq
2novoh/P/GQmNpAZESFEFM3AAasmGwxmwaqzg4116g7jDG8IWmJRow3e+LTK/2Hd
9vLILai+4HLYSReUO/iL48hvtlH2KppII2tOhV1t/PSzaif7oPVzF0sWtQuoA/ix
31lksOUxCxFPCVBvWoFJgs01lX3t1eY/3qrDx/u8aX8Ig7k5CCR750mUlVeuqCYs
eavZyaOWLCa/59pbcRUNGEQKAhXYPpl15xOLLdO0UFh2ko369Nt2TCgfc5XFg9D9
ORE7scGNnOyC0q2jDn/eNOT9iLyYbAnOQ96j+5RqHQXJT/5b3b2O3DZxTCuHSyng
Nx95ztD/jCb6U9+s5gNNazmwBqCV1y166n/UM6/jrexzOXs99ZNZuooqTxGdNj1p
7dQJ4xwUYfBdY1AWUxzjgPj951iuOm8LNDmJnTZsd5vVbxIyGgEac1SMIV9mDZq7
WX+1OT1yuhz/qOJy9UFs5BJinzneDa+7eUexpBKMUmR1mFgT/BilSBVAgLcxiRLM
T1fMnQTy+tlz7JlR7CLD3d8gOdkzpzGt4fMe+1mMT7Gz3y02lIQCK87AmVF/IBb6
3KOFVoxugdMLGpOzIiDLvHwVphr84KKHG5v+eqvWNWuLhYYu5RrGYGwclAM8ICkN
Xg7/cp0wkRQQg1YibEgBa0RUMsqtHt+y1Bzf3u88gbrNPeIbNOmSv15045DTP2q+
Nl/oBL1YQAuzFkLs1G3tr2JRoE2+D2SMIujCGsLFaRKW3suqChIyx0UTwm3/Xacd
zt/D/E+5PLhemj4uDRrcI8SFv511N5lxO904yimANG3hbsE0Od0Ad+EeDKeQcTwt
LgExeU5ulqb7cZgthPgVI2KeCWk4gkhDHGFUOsNi4kVQp7J8R28MhNxinwVQ1ntH
ErVfSf9UBoqsq8Hbsg+A4tc+2S9CBuOtzOsrohE7KxKzuhBfFUzk/bp/Df6SSdVa
HC5XxOaXfQa+KrPcAFpyWSMJm86b3t3oeZOAiQH8/xzrJNz/HpfLaslw3nG6CBky
S1zomtdLZFFKUQiUJ8jDPwjEqUm2yPEpqARHgcVpD+BBmetUyuFovXUbLF8uMHyU
1H8fixKd3iUtggklAjxSYyzMyvWlTs/fw1BOviemhS+r7TntRp+zyjK35jqay/PL
T1+VFuNdNxwyZ8warl3/oQmYYg0hmS52JnZasMx6eVedrorJMvpsrYcn/OSq/ibZ
QCzCYg50DREIPsVazZ0QhbjlKReNMQBSxB8biWg/Vgfs9BcwREuyv2wg6IQRE0Ry
9VWmNeD3krczAbSqBmaWs2BzzFFbDO3tsYKB0Rw7FoEwBVpX+XLeodjtqvlkhsge
aWN8iSzrf+60ZZsgy77rW/apYqyG4M9udkweznyF7NVHqaVwow3Et6mg9LYPiWtW
+rQrVa+eUWMYANR7az4WscHViXTayzOhBfqNz8dIMM5mtN6VBlR5t3FZ8u76MLsE
rb2hR8qz4VTilxJ1ZBmRzh3xN9VPmqstwwbbL/MgANgcK6ITvYA8WnShVDWQKQMg
A9pCP9dkt5rmTqFHtLXJaCejwwNkfWf5/+1ojYcS/Z+mjuerwNCEUzfNEWFe1H2p
K+KrMTu5es86udcyAlOVfzMuWb57BzTssVQuQo0o8ncjEXlyRg2o96yplydQhbmB
kfLYbcXwHxOjg0dgTDzdYUzhzKuLH0wAXW11uNjp0lB4LTXmtl8ZdpLMbnzoSy/d
2lRp4z1G4kI3DI5rShMIri5nzGz03wDItpoJDdH03UbaOSGdB2oT0Q6bSIqOoL2j
f5G6bNRJkS+helhna3+S9XuR9KXNzsktPtNX+/VokOnLABgW6pSjNkXy4eZkBZVe
4dnjuTpEbXm5NQgmMoltwQUHU/CXvc6fly0rTGsp9WxNVXNBMOaMh5PExF9Kn5cx
dj1Yus+nbqJaAb3zb4YcGGTrDggghtLx8aI7HSPiQ/yxxCCHvmbZzKGpa4BKw44D
MiGdAuLReyZqfI8EsOndQtY9mtN5dreWacsrJsdGcfFZ6hYd3A4ZCm+WBkm4lIeF
+ccUf6P97vpeQfVJ7znHEw/nDPrveV1HCuRN6jAQsaRdPopVJ7gr573dvToKsGwx
paVBCxINSVL4PiUPjeAz5Rtaqka1zqkBEBpB3/ZDdoaieuwhfTdnqVGQeNKRhlvu
y7siz77qKIJS7DcV/BDr3/vIgHM0u6c7HYNWJ0t6D+LRbIkcsn541kcdjiV3s6Hq
5adgvVSQjv8ppkHzxN2FpsbytpVXwb7pTwRBPfWbyP92AmsXR8kc6tlFHjpojkr+
JmBR0WU+Cz/mq20FnZCjG6QfwLSJucSdMyaG77IEAdwdoovQyvzAHVN0HGvGiCJo
T0AhSIIXp4GF6D5tH/1p8v6GcQxPbOCu+GGCg7wlIneDZLclAeMTdwlTqQ/4I9kW
3EIBSINDc9r0MCimtTliYhDFGgbn3P4XnjJGHHpqzfvEO+BI8VLEAE4TJRdlGe/a
MDl7H/++T0WGiTnuUb5gddWTGnaTj3YlBHWoFU7R/+xlm+fq2y31AdDddrvKYlNq
AHb7Kd6TDSXVmfV8udS/9eDTQ1fz7yDieSugtrNivGvBcM6+igRr+7L781BXoe4l
r01es3kYT+ZmJRmCu1YeDB+5zGxUMDc3deDJRiFt8EjSmDi9TAyed0FGLB4osR+m
gWDhGKvom5oRHijXkDVQjJq8uID93hQk493DBtgUYni3kNtgpz0O/lSAw6aigZK5
OnGU9MoyrfjTa4al1uYlo5nXGE/XGBspfupvlZ7bJqD1IaabXknqN3dfTL2p6Zsa
u7j94IlYZ0e9ptEX1fcw0yEaMWheH4N+YoNKdihgc0JxBL4KO3ADy/4Ay0hF3QrY
OqfTROTI0WVpZmWGdQuWagiqXUypOLxCwU6OvbW6YkLvK41Dcxm2AZulNSmiagGI
+34xBKPfKLyJI1zoNCmUD0ixFXk23xiVLW8/+TFsTCaUxBOFnvSheTw+HA2/9J0e
B7QFBRDlqIqhNfAT15CnlAeJ39guNFtOxO0MAU9VZzMqAagfW+1S3btVspHC+XG+
tkoynCzwBUL9Ij/hxW7aeTGCogo9JJdw1HDcy7d2nrXLSP14azox9vA33uu5p06F
65Pkz6nQEo22YuccR/YmOXyMGeMsMf1ZEKRu6zNSuYW907BpMUNguX5m3hL/KtZC
PsXe6OrRRlvLomON75MJeP/jI6JPBiX9+imaX9povL6JEcMVWBoTAJjw+sUvXz6z
74m8IN+PMawLk+ZB+Y+2FlZaEvbv/eNi4Fm8RjhnccDwvC1cUJB+8bLmuWyqUCLk
eG2BSlrxR7Jr1aKtciPFMb+8pTA6WoKzQ6YiSy4lan8VzwHpUCEuOND3nvmacfA1
ZxcdyGrXWfr8X/RjKs7isCBbfnyxvmdjbzqnFwhCNWATM+ePaHbM/R9+UEBZV2jE
t9o9uEkEBPBdv7x2gYHjQiWmYz/EMitFCWXVaazyr051h3At5bJWVOOGp4Ea4Jd/
RYnD6cT8yIqdozyN8jocVHoQ5xLLB5ohYuTIDtC62mnxDUCzas8OINHeGb4vZYTq
/ywnrddCFewx01NxcSYIRpDrJLNPprf5Q2+7wZA0rWZOtHv4znZrDMdsbGwnFnyj
eHRYmC90SEbUSLUhwbZ0b3xTh6cEc7T6fivjMVidzYDfXaoDtrOe0srJNbgyZB/d
UDVc0zi4c9vJkXpfkZgZnP5/VZkoxYdGAM+oN2It/oR4n0Gu5GAuiLY+OTtwHXcm
2VPb9THYIZ7oMTvOwH2BQj6990fBQUN2YPcvwz3HUaVI724scTEsvwQhnkUjPJUl
PihjocdtEKrORF5Q2I/gAV61OQdkgTPA507cBecbTqzbGUnK0BzwrbjU87GvgPoN
ukqJUht4jaKH2Dq8J3OjdTzpoP5+gOVDlnEKooH1CqtPcek3USqX2GoFR/luA7gz
HA/MHnOrQfPNR6XBL6L9LTLrtuBttqLSzsYwe0G8mfjczdDzZTXw/aoHtrYvrVAH
tBoBCACV5KGZLtZU7e8ik0xC2paLrAa7ZRU3wInO6MBt9v9PF8QPv98atzPpFviQ
EH4cwfTLJobwzncawzbSzy9S4AIaFCXfaiTyGg9IoiUpqQW1n3NSFmLX8jayDHta
Vs7vgtoq+KDvtqkjEsUJaBaaXhXqFAUYC+jcsS5PlSl7U/yR7t/cNwp3WEhgYR1j
fHk0MQgq7IUr/VnE+uQdKzhePOibyOzb5QoUVhuYRtXh90LTHM5r2ODPMU63S2g5
uRAX/pmjW1RgnYuDLf5W6DMGPV+BvRgxNRnfiQMK8zBx8LL36Cj+/dkqrl+x4L15
zPL/2iJq8K0CUBYBAmOLhV3Ic5PClh/Nt6ZH08LczLu/o3wUUeygVLgfKxhfGLa+
/tRfzkH88i7d+wFPW+gF8LufRxDXaNuuuCHxDOH7Fje7dgVLU+/vtBpb1w3YXX8g
1JvVSHYpvlmTpQA0KU0rMC1DmQyrMKjlEI3rTy9t/2ZWV/a4n40Wz7qar8UhhmQT
zEqy8oXGtfEkzrshrIU/Bzs9KifcLgTb4DwB65TSKxlbBbAcTDxeaxNK6w0ETbIu
ga6zYCQMElhrISyfq+MxQXtOP2OP8TN49zvOZNIfRJVvr05GEt78CuX6Epa7NPIr
b24eN7Vqek3/qyxVk418/gnXElLRlbjRWdAhln1daJEQYEYLfGhcEygLNu20Do2d
1tUqie21RT/YhDguIuVfTLF8+r6Ec/Rm20hLxVmIULl5ju1t/YULbwxEtxRqQvU9
tr9MqgYErnZt212rRK0qq37tR3yEtnrJVkn9XO8zTE+kq15vBeAWA3WfGOIpu2Jv
rIYB0Bj5OQheLoMiffcTVMjNx3IATXqoiJwa3wCLJiarGttTIaHolDeWzCxAeIfd
xIFq6iB0lU888QSLAzJLP/BjIZUEO2fR7AuVXNkBXNB+uEiGUSOK1jWHfUgiAPZV
2Ej3BC8zwmFWJb/1deBlFnZcYIZ1EkblR3Z+KEvz26jHTWMjzmRIiUZHoy4Hxull
sUxAqAL/MC4yDn/IeZcR7Y3D9ISM+17ksyhZBDm74BKBdZUDo+XycflAqyjijAAU
y3r//iiIKos2LmhsTaTQqY5qNJ0rKNocO2wUws7bBARKxhsz3xCXv7hy+ICkJG4g
+si9OwN2NHEK6Eqv0Xm5giiBkBEvW/p4Xf38IYoiaAXy9eOdCjRGGyraRcFIR1Ja
vLUEtieHyJVPhj0374iEMWjd0wxuamDdNaZQlcnuPSavgzdQHNIlAABxKArJNYOu
IFXGjc0gr6nJl6NPZ79XJFPqVREGJ//3VSTV8LmDuha19RnIcO9lVIeAEuRYAcwE
1KBkjQuKxXmG9DBU7hkR/CPzB/WTLX+/bSBwtDYzpuDd17dVmRZ/vwPBT1nsljOi
0vlb54OW4mVGYOeZ+utEJg5hk0/OKVjQZzFbdiYycBX1ZnV+0zAylunLjat42AJm
gAll0h2qCwW9JbWVga3oqkxwgUlpujA1XjQqsCrujYk+I8jKdf8A+oeEiSWAIEAG
TPhutK1QMh216INHkMV/TjWSnNLJchsNbvzXq5eu4EvO4Mn0h1Gz9eMNDnpUNliW
5QZ4j2vyLwr/67+6QXHN+txbW8XMyhDKWiDu8muDrTWTCnmJmJVldxswHuQtrx57
FyIQ2LpyHSvWvZaA1SfWbXuYaGM+lYfRdxgJd7tWJkHVERDAbAm0bshy5zejm1mp
KaSpzYNjejDX/QvLlUuD+JeuF2RG3qtqz08e635SDaB5TuwoYhnLcnklN+Ea0Rnf
TjgMhmN4Fuc23cloIdwtpIkwpq3YOO0xUgv640/ASDxAqTOgqbXMlM/cyqMol3Jx
8VK9gi3FEpETTK9J1LBoEUiGUyvh793ZIK4u0o1tLDU9YHymREeSsDTOFpw7HwXa
p7VDjNE/EtT25q9yjhrCoI1bzGCytKKFWas90IHWNOCBqP6USDzEYh4y5kzZ89mL
mtIqG2pUKOEietaVZCo2fA+dtdjf85BclyPp6H0qnJWvfM3t5VLbjr7/hx+A10lV
vXjM0asSsEJoVWkYrOjqp38YFXihtJLF4pH/i/M+EhHSqDZ7y4+9Zt5daMjxfQeU
/pl4MnaavNmXI1ez8lGxnSOKuoH1PQL5Cy8g7NfPv9kBSTR1GyX2iTPofDk5flWO
r4ix+jnH2T7hBodCxvCYSLHPL1/FTEgKyi7vx3MUGFfMRJpfSObtHGshjveJgPAc
c7apmnC095T4p/ij7lS1IMXl2DeSd3MrZTFGiyLMdnliLV+7Pafu8eeuRrXFDTIk
ghB8tpZMvTT/sjfeBs3QjxxB06G1cYTuUSy/d1IlcPFLdScgH6IKgD8XxtSpNLBC
AepYQItVDFFrywbNCfS4ugbpsJ4v7cLMCtOqD8l5i1ChbSda1GlY9OFYoq8O3uQs
lpoigz/1vG2zbjuYwEW4KtQcm1OYHNnClH+3j4+so5ZSJGVaAAxedh3wTX7d7WaA
+jBahIiJ6DlihYcF0WL9u1RWjR2L2vCn8cN7CXAb4l8hwFc93PiN9RS8+PrPHuzZ
+np7nGMiaIf/FJdsPpP9OyQYOegA7soQSB36tfwKREgJgNSCMBmq6GYw5mfKo53p
DU0pO22/rZqt1kqHFQcWrbtQgq+gxaEzG4D+roHVMfQBc9BRr+G1RTyZFbLOtp4s
zj16u2SkzZWpGt++euuYhKDCT030RwopRfjdxgMw8eF0FCYaWO7bLiWxryKByO8W
rFGGV3ku0AsrGmBy3Ej68YNu2xmdwhVMg5CAuBUEBkNWzqvdaX2SszK5XfyCZ4Pd
oXGzoSBYOBaBhMpar/zMN38Ba/3Aa70kFaFp8cR7aV+IeO57HpThXZ91K7yJVT3q
wdKbGJXwyXSBMKteH/WLKIU2ys15gwbAwoOnh3QdzLLINlSuGvNvnnJjM34uVslu
1/JwpK9EDGq8mJoS2iECTuB6wjgN4FgFVZPGYi2A5ubco/5Xs3x3mn2SvReUB/Hq
LTBPLpqnGXe13DdiarR3kSGw6r+UgDbaDBddECZMB3TWaYkg8b8Cs5tDqzHTH8AD
yIR/ByIQ0V29CW6d13SyHNT8+59S89bGMDk8oEsAb3zRyGfqRw8EIZQHMPIN4+Kp
I7JnBOmsUJktE7Ro51lK6nPQw0PKVLKYN0ibBtxXqD2pT1mQCpFIdG/TIvGT91GV
NgwNLVndrkgLy/DRjnf4lgnZiWj9e5UHESMX68OqC9zjYWlwq+tIjIcyNWQ0Gtbz
E2F0R3klQvsnd9rE+g7inRC6cHS5W4joAqioEQmWnktzbuy2Vit4eNAuUY/xvQb3
jzSPQTkUcirMpldKkZwDWySabFRI2yyu4+zbV/l7K+e/Y8Sxp3WqnV94rs2XEb3N
M+3n3mD5FnFp8QnS9KMQsmOSaAMxmUB51PED7hQreNf8Oy3rAAeoffR+wr+nw+as
v0B0cxYTF82qR797zYGFtItwiTQPBivSvxcn1lqbmkzv1iK7moRLDLXT4EgdMuNE
84182MvdqqI+JQq4rJ3q2CZNOe6vqJ5lfEeDEVO3EtGR+VmDs5nS5bSIbPtQvGQs
PfSgPIekcHrxhGVh9gyUjl/0Xb9LM+zop04RKxNoAra7Ad5VSYL159MuIaL2wy26
Y3W5MenHvw/NfjvZSmalWaHIzEj8Q2AhUOW7Oxn7BkqvsFzkPgEbikMmcF16vtaf
1IDwHf/59nNkhJL5G8l6Oi8vrJXY4/sN4kwEIgLQcsHNcW6Q0EnD9FPo5BwOqe3q
mPmaGfbU+W2o4/1sW/n8NTYouW8ANlO5dLRNp3MC8Vjl4CwLfPhN9ogiklQhSzo4
KQwkk8grJV4hHoNaMIdrXbLBu2gYcWldK0XzcPXLtJvvWxR+kolj1XIqWq9Y+7fm
LcyeNMvNQqnwNaODfBU5/gkOedQN6aXV9vSJ5imNECR/nyxCjRTem3wFYsI1dZBU
Us9Sy8oLr2rIYwR4yrvqreQKPHBGCEBkw1I4EsQWGLQM3J5kK2M2pC+pu0FyHTpT
gySyQwTSNVe1KCm6gnX4hXJJ1ZDABQ5RGWrPZhpoKvu0AtDER3houC+3QW8F2UGD
SLmIr32oJ5lbBv/0dltSiCDS7hE20f8QtemB6Ifzn8JNj5hnCncig+1ITmIWnq6x
lnZIljAVXJCAYwg0wLfjdKQGCqdBcCcGnJk/2kgHyls0siv+sBw1hOJYOG36EvcY
gOThgFork4yTa87ZwwFV/I9fYvrUfZ3ZXwmfnm+DrB+vURGg6u1G/P0tZ8/5oEX1
R/CodFHEDwxLW3YO+Jtlp2X1U6QAviylnt9YcoSMk3ismVUWkUM0Mnr8q9ml4FO/
M53utTl8Ii6dTvV6zOmiNjGQFS6+norWDUnggQ1xhFiWmMiF4H+Sg1wR+ZvESyl3
Y74Xb0IbHwrj1ZI79mCVnY5tbVHsBELKWwEmrxDtqK2bLA/F/lx35AEQh8tT/Mf3
75NOPVE/EdxaMA+86EY1+eeEdOurkaqHzM4A0PwVRcTIDErOILzYlwVJExn0C+up
BT2eu0LdNscuoyqFPNMGhCykSM4IXTsfeKHbwKNpp+X+8V1kJDDRtuh950OhFDZv
LOk5tjEyPeszbPkhWsu4LiMMnGNmsLBNqgeyQU5HkdANwYlVmlmvo4LoYU+IgFUV
/CSOBbOlpq7xXiEIOnmTuPyYuv8GnNCKyv+VgmKqGAGVUAiADrYsSa54MrOyyNRQ
c2wCff2XiWayidt8MAL7qeEzUw4JghOSD1HiqWZg/ygzhmJ+ykDaFJcotuTwELkj
kIPikuYGekUC5Z8M+bIfwEy69e8zZBrdHeGTCFMXQ86eGrp0BtpUOZfVU2aVIxbf
LVOGRpfVE2Uykz5ws+TGXUIByMhmcpT112UpCZfqzTVGwLVl2thCZ+yvguhqkAqV
cw8aPTWzqlxECvehN7xIpNeSa0fI2daFDd4cpYONT/QkY8MGqoxFGLNh4rVOvjUB
mRz20uuGuuQTZwKYXLRbce0G3ptK8awLznvadm9feFZdNHNcGtfnEtTBE8PovvsX
B+R5S+dBEjeEDOQk2zqsSmWSEqygczr3cu4DPLM4ibFpbO+zV850IrX4fUp3N8MK
zY2PfjD5Wy88gcg12AvQATezY7rMy7WC10l8TxIR7G3kCrqPE0M+VKlbhrh71wVx
BdKjj7pSmccDd7PZLR2Ux7dzsF/vgZj/9pScSJl+q1bvCAJGqnTXDdiKAgZoyZVJ
sjmVrZxoMy6nXv6hiq4XJGg/WW162jO9Q/cu8MKhhTFqrTZzzwl6Sq0FAsjyWbRG
8EdLcah3UyKAMlqGy7LyAV3NcQte4iPll8JnByfdT8QGx06xGcJbisXoMJoDBG2n
bd6nbTb1yE6tWXoGvl+DC8XCqMSwqUALNBBKtHCOCzyvUq+WwOygJYIR+D6cTxeh
Xm/I8iHt7hZFah30Qx//WACdJcn2VWiDJmW6dnkqtCxvtBNegNtwurPzvX4A/7O+
79tYEHF8Tn+78cnv7UhC45DaRPR6xItnAUSBb+vf2G8cC3CpoNFWtPCuc2tsReiM
qSvOSTRFFhS5lS8AH2Hoz24/RBLBnl3Bx+zRTec5Mm572ugt10OGRsaw2NV0pUuh
0J+fvSmdSolomvGrEr3cQsmjxzsB7Va1Xx7y56k8BU2hXTvYirqZz4REUuAI7gL6
nhQNFLbkpgNZC3J+MMmrmowOxdPZp9C7g5RL3n3U0aHmJoCAsX9fSMeymXUhf2cq
e/kOwUyAHQXeQIF9WxgcpQyK8EAuF8S3FOfOPm965HM/TCLuD9ibzwC/Hfid4vWI
fyP027DEGHrrRIFF/qJ8iQBoRIldr/UFc5fTYyZOrGufwgdAGcUUGqMTJujx5D3/
0xW/yE1gX2kpclWgZ151K81o6gyAa0EGjHkxPiGvHM9EEC7XMIXWbyxtFpDZqIoa
6gKhoaXlyes7Lrf8KopTYGsb49KwUrP/x25ZPzNpV5YDJqZ6V/zq81xY34ZWROT4
tnuJNyn+74ZrMR87TyBjPhhNy3q0mwUOIAaLdjQTELcv8cYAqypdDLvoT2qdqh9b
7hiTOVV+QaYGOJAQfxNdmJH+lnznXGdcNNHFZBq/lg9HyMWs3WRt1n1P9sqvd6U9
wd1kmqkkBu/1CwML7I2O3xRloAybIG6HEf/DhRgLO5C1p1UVzskh2UULQ5xZsm+A
S/k6bXCbtroULzaFye4R++mxJqav6CYyGAJ1V5BKtcVkrLJmNt2Lm80UEUYmpBfc
AOMGAawr8n4D7OxmQ/nOuEWH9XqY/5vxAYeGBvVPc77M2VkaIJx5dROX17En6YlE
/cUIQ25a6xXP4DCs1FT09ExpSDwgatSCoRAk4eL359f+LJsm89mV+25TLWdQq/cn
CYDxc9YpEDhIVbk6OkEBLqepwrE7LS2DGbroG4EijW2r97rYrbOj/I/RPKpIU2p8
nZgMxcFJFlspJ2+zVN13gxD7StESi1U1Oxknm7/JiOwROdj3CuNPKEEN+Psmla+e
2ucL8YVTljFvqk+G3QAcz7DGmQhyWQxUlf2Y5pjuHDYekVJ+u8ZFWYuvn46KAV8j
B3Y9B5ohkohMQfZbkSqcyTsAfxWOqtvjXaDNApSra4U+HP1Y+nS2Z8qkSWzezsJG
xj/FQVf92OyDd3UpfF6/Fctsf0ADVewz/AdlEkURrnOkdmosw6jjWzxKyuN5/aJu
glxQlSziOiIP46k/D5fJJx3l7euv9HZTd/EpuCPG0H7XwB2u++Xg4d7pZeUAyPrw
B2i7QmfAz37G9/hKsU1S7tj+M0Anf5X3wkWcBNMZsR7enMPI6pIjIazCMJ7dAd4I
pb+h/44jE25Bpo36UeIgr95BMQYxvaPH8Rp9WErq5zsxc82Yba0KU4R1SeJqHXne
73jwRKeiOJtsLMzla+kEPf2OBo0vhJVKGrWPFPVbU75KDCNdb90UcGPv/Nb5b3Ez
wW8K/K0PeT7KvIQVs4knnZTSNdfWGN2AmiO5A8eodKXju0KGWbq3ZqXazMOLDFmU
oXCWkM0Y5D9VrqjEYhjRiJTkZJuJ/j/LlLmohAKZ8fk45cuAvFyiBXChmJz0PtmX
nXZZQiLBAU50vJnb8DO3DjfM3DsikYgq18SGsgLOEZBzf1M3uifxS2hJrv5U6nKH
KqZFE3jJeUzuSKXKDaC3gGzrkE3hzBgShZ6bRWjhEyhtteE4mTvpCI8vOwJWZdAH
RrKnLyGoAoqSn+TW+jsXMZOE40NOEVADU63/2M4xGjZN3apVeJfL51Z3idlyhruc
PFrigWhHYX3SgcOjfOQ6H3bCF/wGl52y9Ceb/zlP/zHvHohoPRYvFkWvMCtiGm1G
KFlxUE2B3Y1goe6YQ/jnp9WMT/qrh9K3Idsz1YGagXbwmLjQd4J96AaCwfBH4R3I
FuJclt+CRKCC0pM8q/vlk7uuI7BHhXjgkorRrfKUZs+xeilWHaG+BGFxooy6lRv0
Z3td9KYbvjReuBnxTsXywWgdRuMEz2ro6xtyOI1GjGyqF8ymqRqkT3sTb+OibEe9
w1XUIPYniEnDIzx/LcYebQNImiplcQzmfS5sS0Zd9jdMYTOpyeyUU6HHc7bZ7Hmg
FGIN0VhGby4PoOeU79tnpk0v6HjGIR0CaUzG0tOC38AlOBF9kAKunCHWC6SXwXTP
q9dRCIqqhrQMTwBVjpOLuSpiaaDLL6ybYjEOSRDD/lsnnuM4Crv3atyE/TocihiV
hvKt5JyiPzqOc9GxjbELZvED+zYmU1ssRCFZO/jEGRA6pOf6qmvnStBIFwndAAC2
CjdvwjBXWF91dNBuswHb0piCwAWhfmBFfk5ZPfDD3wpmLXbeafrgCm6DuedvdTkY
O/2pYOWIvkrqEBP+8NNkvHPYeyTPMX/8oJBRm0882ZDmxX9uhAtXfYdU2nI1FDBN
/B/JuScTR1V1c1YUD9jHIbSas8K8MQmgtJgxscbTvptQLdWQB085loJ8Plmh9iOq
3z7neVXfCHQznxNeuVVzUKHnXCz86WvvrH9RpNar4MaFHjnEb5eSd3Ut6QOlaJWR
g62+s5RMutCG54x6yORamH0hf3GGaqObN4NCFKoHQy+bugDrGIlDXOwneQCdsRsb
zF1bKNFR1K1UDUmcfqMHVz/yZcBk9SaM0ntERJMrnWsgQMpkzm2J+QSYxoX1laS3
a7mV+GfPcJZe9LrmOgD0unfooOrRjY7SIJo0ZknNO4s0ckRggPS3GW5QmaIjTRWO
gL5WiHWUITKdX8h1U+E2oBlVm6/AaeZwKg9RttMyxhsYtGhGjbWMOi+HqN2zr1vK
I6nBAeyEXQVf1sFNBXuP76p82DsVeZFoYDDC6dqt3gV75dyzH7TJzzIZCH/pAV36
ZvFTTY0AlXAcpG5v244BTflHLA8xeYDyGmeksq2vFoQhsOlzBJUUL3cdyAwRKKYR
hQyTwi31QbX8WrXdK1wEwplV6P1NwvDl40ENaSwwtPWqDnNZSZUISgn6bXQF7raM
JjlKRn8bFbpADUoPyJF66wd1xzfhvyPo+ma8xpQ0nV7HX/7nnTcQo0ffRDA7Oma6
thtU/lcD5/oYFu1YKkvnLHZ1BxagsMi05ZAmuKAPl3I/JUjGDESTT7/8gJRYueE3
MB68Qh81V2DyMCI1Ipbogu5YdmF5rfLovKJtnuUSx1SToxUyaPP3w93wgvm5B9HD
x/O87jFfs6JkoJPpH1oCn58Q/X8ZCi6fWn2hfJ1YumExoSWfjQParskKIx1NOwLz
lnMef8+O7HpRpCENZuLELKuJZCcW2lOU/wDInxznzQI82nfZEufGsRKWh1HrBx/r
s8RRbvda/QTJ9kIEcB3pUChhcrOdfsNwaXGjntPIUmMHouYqmPM+cO8Q0YqyKo/S
zX5Aq/3mpw/nAJXnu5Rx6OGO7lvKM3jU4LBycETM6TDzKz2GhxMtjFqfZEfNt5wp
eG8vNZVCqMn3yOFv110c7ChAoPfpeqzyxWsTxWsE6v2x0Kj773I8/5XSxAy1FOFE
OvuPbtTAz9bvmJ6gwyevteWd8gu4cmiITtk1/Qs5jjWMCUpWDoleraJBiTMUP05t
/S+S6u1NY3StvREc4UCkWuYlUzzrDYLFLHaCtQYd5sx1BAJ9vrgtVK+8E8l1RGFH
GoMDQ57jgY9J+HVtLtUOj60jLMmOKCbp6YTntpd4G/fkUdvGipJ+PNh+hAytYOSS
biDpZgAYtZoeRcO9eGSpSeWyYkqbXt/+fB5bZEXrDVlOPKk+yn80oWQ4Un0bB8FI
uwvslc1qyVHqGyO8VQAae4Ikr2scJafUeShqs2RKoRlFMLYz3MZezI9P5nvX9sKU
oTh/B6zCwG9mbHq9H0VRR87PThF04jfrBXC1yxWo/tK57WtcTSScq6/W/TxuwZhY
hgoUuFQj33R33Z25AP8mIxEkXkoQbqCoEk7mvu7h1sIZN/Bp+95934pa4BETEGce
yWi6l9/kYmuKQl6U9pvINM12RyWi+e8nEm4djtFySUlDrDD40Jvn9hlXJXgRvir0
ejyHzTaLHtJYlxGDS01ZRysjtvjo9WZO5+LdwxsPIrqKOP6uWHOpXRjrPRS59DDh
m0ff6UMuR0wN0XY0kQlhgchmnBSjEidedx6RpoKAng/v0Gqwuzrxhm349woqQzAk
Qm8x6ey1dG9gGT7t6GGq+A7vRZ42KsiaS4gyuLdNvyjI3/mqZLfnfbA8kwYMOnng
KAQssEMm2RpiRbnsYE/h1belJQ61pOieKpwGnMFeIdukgWIfwdGxHLVygCoM/b+e
OSgCM6xeRB0KP2A53XMz1yk7X/qsn7xThHFCQgb1Iyt218KpAyeZ4XGBbgkPTcj8
8caoq9VQnMsI5lxVBMZMidcKPgL/0k6/d/KQ8xvOEIwYIc/wi0tiTwyM5flTYMib
aPpOOadsYUEB0+ZidDL62P86+NLInyVqvakmqTDQZBc26eTrYxTploQ0h4n4NWjM
C6PNpnG3jolTYmQpbHxQzk+g3MeR0JjOlYJ6r+Pu8IG6EPz51miwBnuzLZH3le6M
zM+OzXrKCoT47vJ0UZGBDtqqtXl1y2AgRkPqAuoH++ePmHl3K0LZK9y2T8QXq+iU
hU8k4UcE+SI5NxT2CQNMqjX6UQVLTWGDUAvJf4RwtF24eTol+GWX6Zwy8PsUQbBh
6xBRNaaCgOiOBaeiBDQmSwJxOTtBaZYPbfguNgKDO0YQYtz+XnfUVUaICeZk4oOb
1Mf49D9UFTrU3PIT8uXrWtu2//8bTwXun6bzBd8xaHsPWVWf6XhbJ6/RyhMJXSg6
Y9p6wUGhJzlQ3gjyAUX5K98ySgUqY7Ae6UWb3+GAPuob3I8d/uXWzYrHcUUrTHay
ZLdEI3voNJEpgUMMhSO0dwGUP53d1MDmsThCIe+rlR0AETc4xxYWWkgTEx94p8Zb
lXIERufVNiA+NzIPRPqWcs7m7IeaK0sjxW/t7OXhuihwysXYKtrXEq4BS0SPSlYh
RT/gOMnbX0BO1rGUjizjmbVGCg/Wu62jr1X7S3T9SE2Kit/k29R9zL8ben+smxQ2
3IuX9xwdQvgiPns/UdjvvUv+r9ybfqkMxXM1xlOq46iydvGY0smKkb0tLOxDloVs
fSHJ2GDwsys+NtOdf0UOx+zN5y3FWL6+hbfkkZtZkxDkhJYCrTaFsK94pFTKjGgp
eYLo13gCthIm0G23mQJQez3QcgErbAvSAM2GGkDRh6aEtTw7RwMfTxKKLmkAkU+B
FswJ74x4ds8BE2jxZ/bgkfLFy//IXaSW4sd/BvV9Mww2+YAct7Vff7qaJVi6SKC6
r3DtI5oIB6fiEe04S2diF8VTevAuSMB+FORv+/rTht3G8H70mWWAQeC1b75sghNX
AUU9BLmA5nLb3ipRGQvjzoGpbECWHwEYwkueTdH3LHI7rAHxOTvrAO2PlOsTBboA
1aP6ea8oRkqGRVTvGlDd9uU3ephGbkMQf7ShUQi7+Twde2coD0/TDqUcKyZ8Dpr8
uK0hS0qwz+QpqjN9qPxf1mMdX1TpHBME5Cym1lvSkwO45vE3cCRELnlARW+JtVAj
HX0+UG98TyAFcNf7FWTUetO2VhAX+AgeIdQZ1saMXguUj8cT5Ygkb8gFt/zvAVl1
1pD5yvNyDnuABenJ/X9xtV59Ef13E6SdVWIyIkaTPAR57YJMr/z7g4euvj2Ino1i
3YKmSC91Hd6HGD/C9SfEH41BVCSIrXjHJ7pZ6C2kPDssw/2O6hhsN5LcB0FlA/fc
MsxBmVOJGOudv4WNd79UM+Y85VVPkOlFdEw/5nLQvTPlrukdBU60qEU6qDC4D0vH
G8a1hqBJKmHBNmPsTCA6hkjv8c6F3WDJjgbMldQtAKwm+tIpBLb26txN5lqwipUW
OVxie1S5nXUfnMy4g/aSrh0y69Te0b/eOxMKLFdET9XkgJRut6oB3S1oz4YxTkrO
E8iPlt0SvgpI0X/giRm24K9XmAtrvVlja6bBwf8toxjfnoAh+ZIxyoLm3HT3CPlZ
jzCk2H0ZeV5xJUMLcakn4TG+85DvjUZ5bB3N6DMbAS0RO77PmTh65Q+OlnS3xg+o
6POucF0/kdDUns+L4PqntskvHMnC/dsqcxvUbVCUdpKoypogmqgnFv2Ae+TDbrA/
jo68i8f28ZhKyLY7E7Zijo85OehQNU0fGAZUfw5NQvgOJpS9wPsSeBdHFFAPzmhJ
B4hh+n4HoF3KBaO/l16v9auxzdhTcefybVPhPdAubhmktTebsfZoIrAyG6PH2Sxa
QRTv0BG46Gcuva8Lz4QRSH2XugFJmksQ/Fs36NDbmGwZ6rRkUxabDZ+EPy20IUto
+tpVGoqngBvVmnaKC/oCYuZHSLCJ8QjpvcLHa1naDSAbJsqnUM99fhA+htKQUL6E
pYqHthIApYvTsRgxlYDTwKDRDmZ1H8Rt5c8Bgatvlaires2OO/BIjEFEsvAf2VHD
j7EuW5V44XNKmx9bD9GmvJHd1eq/K64UmU7ZpHTPZQ63SbGoVoQ/ZKKCkvYxn6Uq
pQCzqSUAQj9uwJbC8OkpgkeC4nc7Gmeztgnh8S2oguDgyR1MnoFfDbD4n6AHMMnw
6VCZewUjWVFqfSdJDAcJpMXr7xS8sZPmseM1Dfu7rGOfXsZDXMaT32I/VRy2aDXk
E/Z3napJUJcsa3ZLW2WxNl1owdBdr/WvFKY7CNrEnsfHeGiuf0Qnm4Gd+jysMNrW
69fL1lp2ADvI1ZtC5Ah8AGgjPz9JA5ysRoYtq3Xeb2zIvcKnrVSzN1GwDUBr2efe
M0EAdrCqvqdaDiSGl4ZixtPn3xBCo1i8HYynpCEgdTpNL9qkk2owLwmUbrdZBVUB
hY2OBLE2r0JdneKq9lc5lD3G51xrTz3HWY+AGUtTtPeyz0/1KRY2BQAMcFozbJB8
EckXSMubRTPgFniw0Xn1wvwPU+zp5aRU1T6LyXmezpX2M51BzVyh6bwYJkC5TCAk
ivF96odmFwx5+dAIYoNOkLCycpGGM9pif5Bfel5IO6CqDA9+ah3lzNXVYd+yDC8J
NGizW0yRCgV3AOmQpoAyayS85snTcEtVrE59RTXRNrqcIR5/hvzs126aqXi50TTv
um3T3hYxqN/gTp5pWy2YXU1JkHo/j73mA/AoB8RA6ilI+2pL4M6fgNLrBMlDl4fs
vYMaHZQYJIthx/GoMXf97S4jyMPW8iHtJ0M5Kab2nsLnXhzsO2zWGjriFe6XA1i0
Gq7KPTelf8J9p3/ooBjTdyrPeXdHgIrvBHhInXYbWklprIT3c0eYWszJkf4OjvcX
Q7WsvxLs0hoaYsorfRf+zIDMv03EfkB8KOmCaQiGFH7Z7TVmEwpT1vxJq1tmnhM/
oxtkDSb4Z6zg+InAKnVF3qoMVBnlsUqrWXjAlowZT20OA+9rrNg6/xefVOcajr5c
rcn2NFcfPojWAYNN6IFnKCC7Dji/MebqYZXFDoili6WGzBG47M5mhPDNQQOeR3YX
6wtVfBsMTac6r9NrqV72qtC+MYP69PHbZF730kxPqu07zTzzkU3LTaHwuYiKoYoL
OdzFZ0jVHUxMc9L+PvYVzi46c8yY7V02Zv/BbwyBRRuQiZaT0X+V9wgSIlpoP4dU
OxImQDvRQW+bJpKWu/Db4lrdpBtQpa9dKU78tzf9wnFYF/MDL2683MNax+TWxJsW
gWKQS4z22PCn35LGlf0o80fGLcz1zu+qJMTNO6jKZTVPrT1TTQmBTxkFCz1WWAS0
Sl6YY2YTDZgJBk8NRupk5Mfz2laCjaFFZ1Ysltg5Er/PicY+NU5ew1mL8sqhbjde
SC6rqJB3zoJoSwbYuXkEM9fzmmpXJFuvyVCg7pgooIh58XPHbxYGbizLYb40RdFI
ocnkl84f7V23+l8ycXleZx9h5zkYExpzQ0ppovO69GrYGfbMf0zqwH3jIZp/cgP+
a9j7PAkO8ifQVfaGGomU5wUDwiIuFDmWu0psqxkSFex3sE9+HxVwvrc8BpHsLQmT
0n8YgUxFqcbQ8ftGcbIh6C0PSqNE9szYf0ubsKWb/CkfYXsop+gJI0tTnRpnm1kq
td7KFoBZ6kbvbj8j2W/M6LI1Tta5xQwDFF7XPm4WpGzWAGk/27dovvERFjQpsdlG
MfZbRkbIi67vYR1dNLKxfxjHXFcw2ez1X4WlXrfmhOyqmLsDDabfzT5RRM1/Pq86
Yj0H7pMgUR00LAsR2XpRAyiL6D7zpPL+oeM4uBk4vbX0rGJ4fFSG+6ChDTHgoUTo
5hcJtXy0MdcPp2k/RjqkvMxPPo0UnRAGNcRCAt/Fo5av6wypi2mJDLHzXtVHf2NF
Fd1HEyqsA/LmXWzjRCWmiOYQ6qAKr7O2tM26jZuGhM3sgh+Vs1JFj4en4pxPKmjM
SbjThXIrsjxKGYO3R3M64WsU3r+3VY8nM4sZyk7vnRrG3U4M/0ujjSYIQeAXdx3O
veCOvsZ/aLtVsKDs69goFGTqtIwPVuappQaE+81RnapNB5q7L2miAvGFFAs/KnPu
qCkX2xqciiBj9ZuJnpUYy1RUZb0pBRyjRRV/WqGdDimQoZB5/kZrNRtxG61kBlPX
KQ/3Udz1h/5iz5toUbbdimtyHnARU0Mir8O3cluvy/pV6hKagQzgyjBNeYtvKh8l
A90qG3JdJy0psPqYPWQRbNAXdtuFjj89+R8zB5XLkgUBhV3MgniZx2AnQDXLh+YC
XR3WYvmWdAJEkxlKzCCJW80xuLX4/VAwcTZqhGABpQ4ja4q6b5NMJ2Yf7ydZVDsf
OVP/VcHYReLKTvRSBb/dtrmltsRU47ncANHZl93UCHuKcYy3xp59uStzc8HqVsV0
Vc6MDDDpCDPD8sCg9eaVBjdBWe/QVukkqJyrLoyP6AwxZM8S0TNO1TqrXbBFq2qE
yavw9B0cx69muu0piAGi09WAhfB5yDyYwdoTBk+Kz+U6yilRZHM80WPJm//kaTu2
L77wu4ng77WuFJbO4/vLwgFKo1lNTSU/SuRJaOzHt/2ZMc5TKke+PvcJ1DrhBgQv
KG29bp3jNPD6pt4/NAKtLw9XOr6hh70zDfO7iJeHFsft8iiOjUUHW7xBBRtjnkAJ
F5gVyGOKwTgnZQPSaL7i7iHpUiiLj+2QhqHFJZzol1k0b9eP9XjmMJbybBY7Tctm
jMLSIap+bfkPe3Y2KyYbvz/fbZ7kDRKYbYCJIeA2vyHg2bR52IqBOiIF8RA1O6cg
NTJng0cY/Rqk254VfIXTDBOPASy2uU/VuPJrmAqN6o3y1kr1Tao9OpJzAa5sJPIX
HjZirEu3NwAwVmUkXnDIrVrNLf02yWy9z5mUKdF2q1iIpa3NCHwlIxuc8WZlynVS
2LmW0L2ux3X5jDziUoSxW2z2WG0WIaT1tMIfAND+6Ee0DsOaSxCB3TUmT+bFPxmV
eIRmmZiT9XYO+LJfW2edZEBemI8vaDB1KK+DnR/Anx9VHCmn2yp9s2RjEd/k9wek
JGp7Vke0yxq9qPxHyeuDfzr614N19dOzhGKwpGhKW7rLvBP3zFacjLuuX3oNV8Ip
KlvOFBTtMtP3DyNvy+T+biKHZg/q5YVol2qjlzv6tZkjjDdvS2ggXusDScXbtV2U
lcEB4lkGF+VM1AJRp93BWw1w38QdBBk/7z93NjYS/Nf1VcLVINcg/6+mGnEA+y+S
wRQFFjZQXSxJi3Du8jqiRaxuhRc2v4NjuoALnZ/VjxQyIlUz3W8xbvX6RKhL8KYH
SzPBIMZaSdYq9dNC3Yz7tfmO5jrpOPheKWaPXQNdW2giFyPLr9Q5a0YnplxG7q6p
sx6ajQpjZleFlzYGK0aLOVZ2zddyZt4mAMNVWKqi5oF6TVNUoFYBixrXXl2UaLGh
Xibj0EKekwF8Ez80m66a4hUbTosQe6Hf3sy3gqaPebPoaFMl3VD2/9WBPB/MTeJb
ejjKIxqXJOIyHfe1xLzoEC8W+ifmiJ0BZO+h0Yv2wU/8JC0dqEwJVH4mivW6Sn/z
/3pRT63pbwgJklMgW99OojWJ+FU0nWgsHIVURZkJ2opkHjBoGGSucWMGmpgrNrMH
tGZ0EFg069+brwNoCR+lZMaTxjmVZJD0GIcE6JhQJW8kBZn2HMHqW2CLDAdbmF1T
4hdribinvcPA4C8IvMeFcSS06siF/QfyWVfXlHtpqhtoHbX569Fnbt4lu+F1xe4U
PssvDdYjdgKPBGtwvHKfDxD0vJrRaAFFcX5hDZWb5zGOVw7PWftXymiwAweGJGxH
vvI1WWuSflmmOhADWU1ciRSOQwsemB5oejKeujsJ26wzHjOQVZ8kIrFc7YGFZ2fN
/CkGYh07A03MBOryNeyKD3mJf8k+yqEPv1XtG+6GjIdxeuXO52MqZrBTbmtMawEf
Kk2TO6gdLp7WEEryazz+OJTtdGSBQCHQBihiJod/No+cCaf4MAgWp7aouKZIn09U
ST+NRLduJU/+/aiPnqxAVRQ3Ozl/kOno3cDGtQbNI+gRNt1Y57W3VBkFPLzR3mN9
Nc6l1x7vkJ5HwBoJPTT/8U7BGuY4vl+Hn5xK9dQUiN+Wj5ld3wAu2OMXUFixWvE2
c05l+5gmtqhkVuBudQ6ZjEXNEFGn3wN8ct1djxxRYtfHGPUiiOx1f9jWBtxpSruD
jDWeoZubc0QX0E9DCnLrnZct7ub1zOTAk5u2f/uryjHVycAUaFRqD3Ht8VYin4tE
WEzaR3lZSx8F/zU3uDCTZLd1fqw3nEEQo41LQV3RIzOJ2YL/66JY7w5Yy+/77yub
/sAyErf2zTQQqX54UI9ZtV3EJGk4aZTOTUHGcgQMIDnI4LORTTkJFO3k1GIyH+tT
qJfd3SvjfGo8h22TjM0PcQEHuaIJsHH3yiImFmpKV9pXngZ910aoMXz1o5yGI9fs
brNcjVBaIc2yO/hNk2obM/NNe8QoEZ4LjUj0QwQQTZy6iFVtN4KVcMZMNF4LdJSn
No09R6x+DM0bnq+MjNplxq9hwSvkHF9NY9B0s7UguTb95nwPE0GIk3OAkvSegk6j
wut5NbQLSeXmP1yQREBGPDoLJA75Q9YlFCCjRM11b+1NEoo15MTxPsJ+yDWL1aoM
Pwc/WOQ9miByjROwoFiyQJN/PLE6mNx+KNI7BEOz0nWh8SRKgM1gnj3t/br4gRi/
8fY/9ehhjeLiQijUZn6LAvNhEnY7ZzdBixnXmM/wEXtkipYUoGTNLz2fkXNouBFI
+PGmSiSIHfArPSVF5xoMaJlZhWab57wou42ita+UKoJZK35di+rFJGD9iswltz4a
wNGBVvBil4hQAIXn/bixbSY1lW1F6o0oATr9+AHjrmoCvr8/OyC1PulYnwr3c7Kz
AvPPsq8lpTCYXE1ihubNmczx7YJnmv8kRR0TB1NoEk0Hvrs07L+zVORa74GDQdpg
pseTveaqLz3MDtCVHfXw6c7PGISyeGkFQj0mrTuTRMG5Ki/5/ZLNirZuvaQsB2rd
Vv+i3okUHUIu2grrSUZT+A28KFOx8Q3WZ/pWwCvFGp49nkLOwDjh0X3trKi0jcZ2
UQsFBQxn5x8f7PGug8/KRt4BMX+9p9ThW5jH+bRYG75l2hTBB0YR89aDy8FP1guw
rviIxao4JEob29oPLu91zeZaJGUhn7a4GeGUUCP1wztvBl4jI9SZUBQA8IkNewEP
aTyrIIqKyf0oz0m0G89y97SXiA8u2ZNgWXAbAHyTjy6UoScGYqMAfpwxszLUMa6G
GkIMsBtraP8F9myaxx2cBkKvx6/F7UxU3bfUwnI8/5AuX4ZLGJG2U4g6ZbjavKol
CslGDUtpd8HHqlyxi6kVoIV0boIgav9MXPq+qv8AAo94RDO6RP37OCJVjU3FXJDu
4uV/3I16HJFwHXtLWFENALja9gA9BVYF6ArJmvM7aogdBgPU+zWL0erwTkuF+gRr
iM4pCcC/l/bV+CRxmpySWnDjwpyhL3RhJm/bkqIoWT08myfkcvrra4qATy+NmBWd
9IB+l/3s00QXVLvhZgNmDJ722XswvEu1YEVuUi1xLDi4DJQEvjS+1+dTTmACTRZS
ci9y+m5yt6CAE9vDs62R3iYdQFCR69SaeOuYqgWYjQHToZ+UUZMeWecwDgALqgAN
YOOAh6vYxFu0P/qbJSJF6mt2zbcJFj2fKTXVhyF3DZEEG15vVc3KWxJ/qQJQNERo
ffyzRXh+mAdezAMhznDHfQwA/1wmHvusS7xKklib6lfoh9bncOz7aH6Ih7AB+1Ja
zRu0or0H4YuDiEzJwwqmW0SFOTiBDXm+1VutVnh4bivFNauWi8hP1Nl8zYwhdCdE
LL/czhMuHFBdy7FWZ1VyyeujOLgL6B2ZFdU9tdISeC0SZz0ryKQi2+xiqyo8yBe9
iJVaXeVe0QIWWJFHEBJQ9cCKXTN6O2N5jTYuVNEg0/G1aPb1oVE1xIIc+BAb8LRK
y/XcNhxoVC34LZDNa4eu1kC7opR4l7fwFmcjho7IBKDBdb2aDWhYd38fhl+w1DV4
IHvToVuA/+4IVfY/8mYoNWMBGr40HEqxXtWqF42U8Xo/w5dK173W9ULBJweGFxd+
5MSozF0r3v5mwnI7YvdrtoqHGrowHsRVr+a5kyACvdkKXSpTdy4AsJ1kOeLIth64
rTOqvdpq56ngK6qBWpF8ydRkDbNrPFS5Kfu7wq3MWXT06dEi4YkmAn/oY2m9j1MM
5B5uu6tE8ciF1t86gG9Ipvc1m5ayylmZVBcIOrQtvhwZsEL2Qz/557NqwC9ooJOE
eFY+P1kKwW7VpmtdSRqhOS1wDKNnwy60msCFta6iR9vq35boyB7WcWfQEP94v8LW
nvsDflzKlXKxVOmJE2iVzZa2zF1LhZXOKmZ1CNUgh4+fBdgUXO+kwE1CblJn9zr/
Jl1yt0z0eNLNsr41KC+/H7rAJFtk9wZ3kHhq4CCK79CzoSOE0bVcRuncFiC2i8sq
KgDqyKY4FelKsGdUldBGdmF3m1RpNJ3uOHTG+wbQRLJZLV1Xipd33DByqzqbWkmu
ZAyyZ49XqR9Xa7eHBo3NvDG71tmDb1oanyH0d4OyToOVpCpCCzs4UwEPJ/e7xHvn
P4VblTKDRSBRhc9RyIKC+lmDOPrdvYuVzvsUrwEYF+mx20Zz7wCvn0vPVaUfAGHv
PxIQ+ZSzOYOawQFJN2xVhQNcWXSZzdvZg4vmWhdhHCVHJvsdrRiT4/TwDwluHhFn
boeG9HCM3bvnAbfULjQMr3ZR31OTKrlnoQLFD5rHd0UPPkPuGosY8ZSoZRuSTNAx
XY6PFnhcx+Mlh+C1VgH3+kR1Zx/5tYHTdXbZ8mnvBmjxpRiQJn/pKf6GVXVrY9PG
gnGpApyMKufsJg1adG2OdRhpf3L4v7eHnQlNFEe7upvSaZWFgUl/vQO+JKHKrCr2
XofcHqiJxpoSJjkmxFYcL1NDmuWI1zKgd8+3ysZoIcLNwKZDwaTRVR/uW9rISWn+
Z25h06wVNJM/Cwa5wn6WT7JkFS0ZiNzH/3RkA+QXbHS+ZGg1uKoz3pxP6fgQjzay
dOz0yKR1y2pX33R8bbrZE4esQIStC9Bv9SiwR7Q+McGkIGbRYvniXWmwgQGri7iF
BdtTipTPh9q+c8IqP0f7f/9wqNodqzUVRdzRULNix3JFhf51HXc61qfStUYcd2GT
wcAYvNGjgniClaUO7k3YAGN/yC3hTfcpz7cCf/2wjY4BPi4+1HJSKdtFR26yPshy
IDknlAHZLInhVjixpyOGe4EFcklR7EZ+nLyVBLKTjaT1G12MAEtEP1cJ7hf2X+0j
HK3F7CZMTQGCMcHFXGfbuVcuohBTpRjUSQ63e6Bx0B3xn5tiiJnQMd1b8MrnvlTl
cBYBEUl+BDImKTFwq2FtHlt2aXyPW32TCSVZoi6zGxH0HVqpznTRqQu6RjHIkTQB
LJrv5LmgCdbwv17Jvqw2b0MLLzJDDVZy6SK30cGGA5Modt0S3PbTseAPkNTO7mOa
dSsDW1ZukZ86eA07BQuFmMnzLlMsplCNfGnCA8hI/+KxQuRz3ELsIHYySQ1IlyZk
w0iv/KKLUxHfWXjcg7oNkzQeNz79E4eyknYiZesFw7gafXSFU//vtslELvO97Zyj
mqEsPSLwuq338u0oslxU4IM3CQyMBqWI4nFKPrMFJx42ishCtvd8EHxJ4k+T+Hx2
XJvXqHEWeajTe+7UL6Y5bfob+tBJhjphn/KziCWxwWtf2o32n9RhrSaFZCnhoWmg
MfXyNi3ZbwKRqScU2NBMLpLK/abup08kM0v0/ondFKhzplkXIcwO9ZymiE8xCb/l
pmenYpv7bna+PYU5Kh1oeAIsTn4vYuZwoAxlFG1CGp9mejam2P1s5/Xs7EcJxzcE
73HDQ2ApV/13a5FSClsKgpDUcG69vQ4QXu/UCybW+VEY00yX6nEoE5Yi9BY9/vWN
wW0VdqkeiVjrP3RszEDjz81ieGxBO6M0kxlz7v7FliiX7/IDes9TOgYcQHwFPzKr
g9PChV7E4+3PM9NjARPL3YE0FKEkOl9rjL3QYUj1lw4wXS+Vprjtv4tfpPSgii78
qHoRXxdLRiFrdDXRysvXi3u3qiIvGHpc4yYt1tsGEYv8IWCT+fUHxpxMJMpqMSD0
kfngCGNpCsiia6lkA1XxQxkPYLTO9bYxiz9o3LK76kKfGsMHuyOnELxMlFdrDo8b
UtJ++TVXsknh0D0RtoP73WlADoIC6RHba1ik2pR5vkwqzGuY87igR0x2nGWiDB6A
foQYFtzUP4P0VSrbk5beXehDWE5Dm+T2zS7K8jODpyOTkQVuxyqHeloPcbXAxVS5
ETzlgKYbpGmaoCHvXqEnsHzJ3g+0goWS7l1ZMYwAfE5c5GG1koy12NnpvAKb7OzW
uYEtMfMSe1UYPXsZodbUd/kMJxtDGw5GoCs35XAEaX6K63OTr9V3rYjD72vvQhzv
ft30ROvCxfwSRVWCNZpEqiZcMFz8BtGOwcauwGokb8w8vzGfjS5Y4PEVy2VakW7A
Ia/cobdGdsmb6rN8NpWKnUBy7uGID4fFJt8SFqzcWkEz051cFM1P6vBmNnsbc9Rn
R3nJS3OeACDGE/XGIGaIiA3mbnj3nD/buwF5GeG4FPZgBTRkK7QLbR5r6GxIPko4
mLMs+as5mcmXPSRDRwlOgYoUTMxn6tppFqyHQ6u0OIBRWTP9xbSJBKEJTGRrl5Q0
jNrtwHsgi+FI/SwvcrFvYGHVSOfVIoinmt3yws4kKOHLq3EosFHXrof+b5bYiMEb
ZkSk9D2XqxlzWUC9IsBehayRd0ZxHAiTw4VciLUFxX2yYPvxR00aNgkDN1/B/9+c
BAcHzgYTLLr2wJHP0PgBsqYVcgZLfg4v4OQusVo7YJZYoZlfbkCzCRiqPr0k+BRb
uXVxsp8OXLquSidAnvFIWmUuNwREBwSxb+IGuOYn1XHnMQSYJOPGcHCvOWvFWj1S
4b1cX6wQckGn0+9tfPJcKy296TTOPeLMeni6+vqF2y2qouKnGesFGhlnwIsH1+xE
fNGNz6mKiwceFtd67ykbmABJOvWkn58dJktKXmcsczSHb8PQq2oNLAFQAY5TiSJm
UkN6BgpVc3zg6/zEj062z5+uWqMb4qxdYhHzm9kKHiReZ5x3O/tO3zYcuQcFyZcb
IT7H6x38r5mOhEPQNoJEuz7Kyi5T3MOG3yQBRBsFuC92OVXzlc25+FjtzaU9OMNn
Hm6Ij/HFttz9kW5YwGrpKGXIo6jQcskVuj3w/fBAKxPmDqVAERtRitZncjz1DoIb
RT+79StOIuCrZs7TtiPvfyPXSZIMrRApfjHB+GBDo9tTHgw8fTJu807y3oizgWo/
MFMQfaR5/w0G8LZ752PXzT9BgRWEuex1Yd707qUhhzsRe/+bx3Fb97eVd9KGKlMF
AO/OhEHsUbtLqDnmBdGbMkvs5Io02PRgSiNL3sD9B5lHfmH+vcMm9gV2NGKwunVX
u7uRRIW0Z9T3HplwSSoyBNZAJtF1ZN5Bg+AEsFz4U9knwBY4opcCQaq8K6o2qx7S
rWHIqy7bqFekyFQ226AgXLOAjF24xz6iWBoMX8wZyWGTlE2hTDsLdW/DQlKV7rcd
vtwbN0xZAP2XAgeNvztrCxxZ8K9BgHiLppxTrLf8ZGamgLkbIAhKM7Gxb5Mf8a9v
X78VUMPqLFOkPO28ELs5srYfZ5Bjgjv47RE7oqjUVpH+FpyAbJcqhPKuA17Y+TSG
f3v1Wntf0ovSFtnI4jDx9qmgwESenm973yH3aEb+jDsRBHszL9IYPL8kPISb3wkF
gVaK+rOBgEL4KA55NQ9+uEMfobGJ6IvOXxt7YH6Tdg1qjFxwYLBEgODSiqXEJ+KI
vOvBOBcl4cITkuRkjCwlx5YtCs9aZqjNu39munxsQXd6gf2N3+2hwwDnzgEfp/q8
6JxYiuHF3n3jNd1dYLHJ2C2ioumxBrnU+nwN2Se1WD/dqnff+B5eaECYBy/ToMHg
xA3/ORD6zgkgLxEuhUILoMWw1657S4Cp4q2Ozne6Yc85CgHRgIxByS2dqLULJmA+
51TZ6pmvClJQSiVTDaaSU+lwgK3aqbFcDBaautFam3J62Asd3texBb4aMswTS7OH
FbtNGQ8H7ccX7vTHuQaRZ1gnnEF0Dry8lGbZinsdupkvm/q4EQs0Bz/kOoKA1k2h
+foK69/OM1f1slkP7bl/Oo7M/tIItPGbcPH6tAz3fZQVCKIsGYHHvBBwasbCzsE3
qqKH4jA4tiz+Kr20Fl/7LG0QRFDBmxgWHzmpWmCs34H59zMs4QJdrC+R3ubX8M3V
kGAanKhDWZmGdvAB4oyw+yfSN9CHO9+0D86plhWjdLHNmaVeiERufDqFZQzL2hht
vNdeJ+9vhUX/lek/qhMOnCzV9J7Z3zkO49wHLq2Ti7ZI9/mATRbyGmNr7NCXKdVq
KYKnplRiJhGBtr/g6p7BvAESE4e9pF6ZpnO9v7zo78GIsiIEUMm02uOKUtXzH57E
0EfbdNEC8WaqyZyA/r+qNXdtsViYuGQt2SiavTGmxaX2VPexD36WfPvphEgJGGrM
x2JZEJgHu1BQBT9BXDSeax5Mxnpg3yV2E4WmuqifDVDQ3i7UTaMUNadCJFmckZkw
hf2mSGW+iqlKgST04IJx63KAmJ+HCTWGp0bAa0heYW1IsXirKJi6inF15aHwl+97
/OkdV2Lm7KpUnpUeO1Uv4VOf47Oa3dhmQjpXNkfygzjE3VgFItredU7B1/9ZTDcl
vSB+HUQAJlhRx9YcSQDK35k6VavJPiI0G6b1B85vkvoX63cvUQbQy9e9T+K5cvgk
YWHkNVnzuEygMhGi08m6aX2D0rd8YyZmoIrZ3grJ7tiEMZBoXKesdTlDesX8hdIG
q7M66olWS1dkGJ437RIkz3DprdFEGVFve/D/52Cwtot8t6qCiXgk0JYiGGCJcKn6
fMGts3jKHGx4onGPPw+2W8m30xxvFERPelAOAUtdUxpu3dChPqNX/xeHUL10ncSM
Un0QWSJg6AlJ+kwhfX5UiPziGsaPT02oHLBjl/VvvUl7ORAH8FQ/rYC0FANBbxbT
7CuEwInSi5du8Vdoxq17yiEt+g8Llc9UbbCwgS69BLkzpQwxdpX4Aixh8PKtLihZ
/wQCsyrwNSinTGUavx/qLD4pIIjPhRmGcOiask3CjKESFW8RlFNuNHhzNVijJCBf
w8WIfCOjGNwZE+U1L2chzu4wIHWArhQkpo1oudQNxUzoTHpipMOPWkJihV3C/xp6
do7bHV1DxXXg9uvxLQh2LoEICavuuLqpBsfX2CAVWFxiWfUTqMSKU/dcLT3hJCD1
ZNyQTeoLC/VM3nFgeIi7Fe2MfM+5PgRtFyzi6n83YU6If2njPscudGWmig3Sgh27
9yen3F01s58vVa6ckKVffkiQ5jmAqWLMVKJX8suvTFuKbXjU3fDP41q2dqfHLgYF
lH0XhmXCGoLTKL1mQBllajwLYtk5DT4GzNf9biS27enh++fdCwdMzOnNyxhkKh7S
Bo9ewDMjA6BYNGtWx8RJ0WuYcDL3+QhtoT4TXXcMxBwpStqvTOZCH6LDBAzCVnfN
fGL8ybyG/F5rfzP4isXqSol41p9h1fcpjQ7U5oyoFQ2GgZCN3KCxIo4oHvqLhVC8
1ojJ9DG4FclLe5uSIDUee24NXn1lqwNuWO3Oy1YU7WKGTvsVFxRze5FlIrspCPSM
PfWmeZy6t1jEZxCXCCYwzs6c7W/ZW9PkrrYiSBUlclQKsSvu+lTRLdjPrSFUP3oX
FAGTS9K9zP7dA392aD98QpjBvhtZ/aBrwishw3kx9o9w2O+h7IuWDWiHAuhwpolk
pWcA4c5hf3si1Fwiv0LXSY56BfkjP9aSZZKCF9JZfoal7dqd1nEPKABrBuQf5Ias
SqxDjTq9FqOT2CSAAQ/QY2ocdPDxE7S8Tztiknl5d3g5K7TyUTQ6SFg5O8oyYKqf
wS2CFLzM0/moaB44mFPrr5Yk046+hSZMXBqZwQFEuTu6dhch9a0Djqmv9KKXSYps
TUPd1ITdGRVv/ERjHG/G0y98d35g6zT1cDbDl7RO9NzRTEkQJ/ZIUOq7Lwoz4Npg
pJqTcZTS9ozN/t+olVtEDUimonMjOlOnSApLrArU8ZMAzfmsR/uV78JkyF0t1Kd+
uuWinO2ETzPnY++6AmfKmBriODr02fDtyiQboJkr/DmaEaJKwI8HKKV5vKipKvL5
rDibFkPecSlMPhrk07D21mY8V6cNPIeQlb6y3SZsYuEcwIMrfrP2N5kyZzqy72Yb
mVARLghjs3Xk2BQG22f7JTrKAhLTZykmCjSFoBuMYPE9ec2S6bccuUO3Zmj27q45
aWOQ3xUJHPN8iD+nSfzwTByuSjXdL2euhG2WfvmqcR7HshaBvszd4H9rqs7WQqwA
KM8oAnBnk2pApZqMFkmtIR8GG2c4TcJ9CXNIkMs75JiRNooZktGpvTrrq8glPmRn
36IcslghhGyPKoY0rTmXHdHsoZfbSwtM2XTFDJb9iNeah4yWpX3qU4hpsIvm0oWG
GrcO8m5MRGowEqQB2JCqAdcmhCf1N3wGidDTMK5IJrz2f1L3JYzlNnfJ3QuZd97E
u7LhjG9aP6Ewzjb8f1q+mjgRzUqVaBdzymdd9C6l2ovjbDLobhUgAmoyt4cvVkJc
pPctAFawqYhhODONT4UJvB2AtjlI5JjlRUHpA1nMuHT38FvVqVqnI2uzzpzTZn6R
12h8pBPaB1i9syHHRNr3BH7ZYu6VUw2JKuxfG4lys+mtwJy4JjSQyDCN5O5stY57
XFlAASS9OSO3AFMfZ+v3fG09yQp247IR6sCvgH9LkBryRRI/KqOyTetPvO0PTlVB
+QtCMxMB6/ufP0mp3mn+fMrq55RrYGO14qUODnPQXc3kB2v7TAWSvB6WcAM361GU
7g9yNoZjLXqVPR+b2/gp5YCJozSGSHisq3NFnBDigHSPKZ5J/KOSPbyjH119JE95
oZhlrGghOdREUq4TdrSGWZtRrbXdnqLvM1GqXgQumOyDXq80Hpy3DKGBVEx9Ghjs
y8sasFEa7NNS9J37Y2RLYFo8TAFrBaAJBbSmfZhXv2Pux9j47BR7KXsEmw9yAPx4
iDAvg3BGEVjn9Ap8dJvBQ9LC26TCRdmJ2cukOCkwaEwCH3NAJuhWb/hjpzIO0thN
CZL7zQkMwSbhSF0GSQuqlyIgUBYQ+z65uTsCINtOOF/STaarY74UAhVuys1ugeYp
sWou30p8yZsS+2yuIgX6ZLurUz3toVuxxDPpxpTxKCqp5QESwrWc/kDmUi/2uppP
xkBxO24x4uR8H+HZ+h4r8aKZSI15Uwi8h7b6fuAkx+PvH4dk/eeq+nVEkv6F4D2e
xP50xx5Viduv1P29JgViWwSdhMrxst2jvOmdQfz9FqyNgFwRAvHYVE8kNj/3nxoN
HedV8WLRvV2uhPXygR9fdM6fXn1sg2R0DosNLQja5OREZ2V+6EXaEkuCh8dzYOFr
Kimq9hcAqnCuUvk23eJLfgz2NtFTGSV0UpQOUfeRpTKaQkzzfU5/B+s7MnsRRBox
EjaOckgt7xQVPPh7I/8VFkEP6++V3JzTutNIt6wRgTn0XYjvw4gL7ojdrobQVWQ4
HnFeN18MzduzgytJiY4VyOX+mPT9YGqmS8irpX+pAcSrIp4i0MXJhfmGS2tzQ4Fn
nQFeVkVsHgkwyQVYl6BW3DmSyV6lGWSklGPyWUFg2dftFqQu43RWXUaba3CiKMzJ
pC8uQ8Cra48Rapql4+x1XSe5OVM0PjwvPy6a0ISoLL+i9Z/2y2mh2P6lgaRubEbv
OLWpSwGppi3j+2ORB8dZomP2GBUd4CxDYTLnH3PZ987PvbkcbmegKIHUNEbc4Xp0
auITAT6HFRQzcwqYxJj7k9tSilMB3GHcqiKpE/wE5AyYmjBW8iU4pPBNBiMLYYnP
VrXi1D5h9Kn0dPsKA7KS1wuP+VRHQNm4ex9C8Ti7oKnBdqc1SOd0biYMbmKbBpVA
CEs+64zHouDS24lITKCqNws4JfiLOPx+QvNeU9BOfcv3H3lsO4kQpGvKCJi0Bk1F
UtspXQMwEuOl5AY7wZ1m22keNXKYBpYXRDqNV5AUCY8S+phYPOnZCZhGArj8yuWQ
9RM++yN2+VVn18/vITPcVRAAE5rMaZBF2L3cJgZhZ1VPd/+39CqErGUhjVJRZwtA
y1LlRGsRXM5XH6yf1bBra34uI/AxcnFoH8mXIi8fbapL39RV5Norc3v/KLECAOFH
NCJaomc5tPSOcxuF6M56LnqyOexr7Zp7ilCNyqFwYgziKaQUekv1xlMyKYJELAjx
8wnFbnwD2Nks8brn0UlpqoZLdi4+CF43c8/NrZ6Xp5eE8pmLQBuHZ1I9FjRMSV5T
u4nmAS9e5yhICokrng0M26v/h9dFZabcg3YTB8iYQ6nuSLKfcRB3PfljTT8TlEvd
Q6ievdmxHARphB9+2uD4H+zKsSSIDt7Go+OFmG7tU4M6UOyyTd/pLDM4v5dgoDCe
oO8ZGzJYMDlaRH8PdCUm5+rzCd5HiSSQvp81KjK+U4vFIS50xcRiVIAVmWH+5pVI
8r9ZOsRyy8ms/1nl330ffkGIzUW8tOHxgyuracthWSFE4FsAwH39t5K51dXLqtqY
83Zjf9my8zciIV88HkKZce2z7ppdY4y+1N9ybzyg9gqBMslNymoBhlK3ykcwrjvD
a3G2JRx6lXLUqqsbzVEKqeQ+1+T4Qp6IFEJ+KOiOvLG9vIqfP5heNDu0oK/ezNxt
uz/1Xz0jq4gvCHXwvii+/VGnk3qJ2ULQbzNc0F/bxscrAgX2khthGWbKPaUASOB4
t6/oKGvcBREkzf9Lddaeq4UYVy64B/yI82N6sD/hH7uEC+L5WxmzegnERKyEMqXN
Y4w+VNqorD50oxWuuCHJt4+VSgEdFBiwSFhjPeZInEIiPieU6CKxtp5AtvLtBe5n
n4vpl5CAOmWAPr08OboPHZ0/hLxmpWnf/MJOk5DldU+uz2XOuzNZs3pROmJFyXpO
k9vmA2M4xWzJrHSi0MkbJk7jNazIVnoultFaB+HyLRYayiI77uwLWCWgAfJRGl4r
xOf5rhX0IB63sk5/aEwdwp98oFJfANiIa8iTd9jR7qWoB1jikIWc7+cP148igqc9
gcOFG841LBYAP/b1jhUg/g5BFpHlgNtQlodByVa3lLjHKudjpKNWgQ2kqS6mwG/h
SuPfeGa4FpVYyRMAw1KBPmg0ME7ypEIiI8HCMH5hks5R5tk941d8RDhOfNllNyTL
gbpYYmBVu9zdNyHOggpGrrXsVCmlq0sKxl3E9W1kXi16Ad4QeO/wsm3Cg+DbHKgu
nCffuA+H/lbkZz/G8yaoHkC1UdR3RgHOm6LyE+fe9LuececcJiJngtyyRmqC+1Bt
xzYe0ba+5/PdULPs0OK1ZK0lVMfeQYuAfww0y0SH54J4KBbF4FnIylNSBYXXe1yl
0+NxBJuEn5NMsAJ2Cbl0h1a805IFUZz2uAxbmLsFCooF4yc9cBxKUp6cgAY+skAX
Ui7Tpv2vbswQ0ppkiy3fuI9sAcy/Pf9yrxqn4XbnqEQjMPY8o7z7OwD7hdrxktKV
BiA95V3tbXZeKGzdlMx71utAipbDz+YT8Thx6TBvDUJntQCCyWrd16u9hpbEcVAe
0pP+8BxDugFapk/JG4ttgP7k2hmHYfzCEdt0O3ZrLvbnnIqTe8iDFj0k1jg/Zo1s
2W7j3WOBuJeL27Ghcq07ipCU/rV5puHrkP2BHV1em4dwCvKIKaYbcRuYJNx6tbKl
7SFqSJf5qVcc9JRVhIettMd3XebSSfqDOlUtgZidcbjITHQZIWTQrl8Ju7sNG4Kd
/5kVPJbYqKj37DOXiJBxdgnR1Wveynv6jFckIIB/A2yEhzQRFooiTdpqpddDL+ym
ZjRupnBrP34WXJleBD8fc1Ki5sF8ceCNcV47Yj2COq5nBtqiSjKAJ6tWMIJAfEN9
zB/5Cs599OVHzXgdffPFgW3e+00x4S6fDe1dWRmJV8zXoP0wgYZW7+kRsyCjdcOC
nVG5pbGzH7DHV4fZmoZdvziTlLuuV/kQEpHuBAYVmtBG4uP+vZ4UC+OELePpNXIe
+aLgocUjOITFrPTyqcG4UErkujS08870nEukiHmpRHUitadNgyHnBkgSvAyrC41+
c+ydQeGoE9xPwN79u02gQMBSXdvZ1TjiknTATxVSXgoNYKicPNodZ7fkdvoGtQ8I
9U4yiDSFf8lxvKFG8Sfxug5+OCuBApLAUyOTufmXCgFkwgBQFZxWiB2nF1w2kZuy
HXYMBFNp831xE6ixoohcbvewbtoTVJiMcryLYwvf4CV/GS8AttDcQiCTLrr9utAn
1uP17saNx70BFwc5s+MyRVxjxWAcJ1KU2qs9mCPlkzeyBWPgtFQc+lDK7AvaJSX4
fPtU0p8mLRTrZkX+V5SY0lvzsHErPIqqRzsmHK64gjbJEAPZrrcxOdjBRlg9OUZB
pVcfDdfNVHZnnJUmf5BiKAlXpksChhHaBRRtmGlWcFToasSV4A22vuJSKh+l27O9
ueChCsIWy8w+paH/ocnrZKWxcXYFkysZh33BwKxLf1EjueXGZBaDf3V2ETWAcdIx
eNtpQiPOQOA+eOXpfCyhfrQNGW2Rub7R08rvXY3mUJZuzPwy9VOJMJSCHjA/ZvXW
EF0v09VU9t5QDFkYhmvDEnJoyqhlK89HX0zG9GyEaNTG1AzK69a8FsmHRQbVzxYi
FzU2gYaDpURZxU1rkPm1dCK46MPNUfuytb2vLBsjpzxwx3Kc+eQFXxetvVnQsJtl
qbT3SkA5Ad06o736ZG2zuAQj9M6wjnOg8tWxylG4jDs4ZuJVnbH61ETd0qRFkpKN
kr5r6Op2ZbVcvDL74KwY+MzWwvV1VnhlPypgXvdLrPSP9D4IkERvnsGzSfiofxm1
BlTQ+Rtpz2T+DuKh30sXiZQvs0sOpSOGtUg2YIaA41SN6Wg4P8+MFFgLw0PbHovq
K9qD31d59gg2cHDz08v54YCojAtZpLpGvPSoXma51c7VdKd+OajXp9FziVgCWtoy
p79vCjskivUVoSAscsK5LTuCRiM3aVLuKG02F0xHhAdJIGFawk/xDwMk21qOvvA3
yRz6dbOH3yhts63/oyphy9Gu886wiEkueKrFJezaEJqd60As8saYyoivGfeWyC/M
D7l+k+ArjwbT0tzAjZe2fqKGVq5Vr/KzuPpDDbF330szVfOpbbqoGmWfm4AkXWLg
xcCuQs6zamBpfgBwrg5+GhiZSivmYUQLtVNBeIkUayLakeLZgq3omYetfVFx+NaE
mnWKmdQckNbIy4qztqp/CVBhTSGMG2aDhn5SdNXyi9Ii4RtSBG7fkC8CPw6x6ALX
tcsCLHZm7kdOsunWLDRiwz/B9GaapgxruPXfT3CUEVCVzRQGy5JH1GlvrLnsQl51
69F9FfyXeuIhDmaoKqDI5KgArb9wabstNqN9cfxDfWi+6rSuCE4fUfrgeMfenxaG
Jk/Vs4RYTvyZZbSjc6J6SYQmxzqcTF5Rn8CEyHvK1zldvWiu1eajJnbioYtL+Q6s
S9lnERi4Bjhq1PyZqh+tK2wNwM3CCO9JXJnAQvLLmHSZf7sBhpBOsQlSjoovexnH
WAbGtJzcQlsZLh+CtFlSVIQjbchprB8VJZRZDq1g2uRSAPek2SAI26OV11hBVjE9
nYkS2jclFdVo8M6Yn1zD1CMxfiZNiQYU3cVUlFPK7QkcwzM6e6eHqo2XqKNfTTVz
NeSENXcm4HARBwbzkY9VUpFCntIe0RVLdtX12YChJ5vneViAOOoq6wvgh4EY6jZD
zsU5iRzdTKoGClDjentL7zTTPqSo73/otzz7LjZ7bUiwYeaH+0piH7A1NiGrChNU
N1hp+2Pw1OuFPN34DDX8F+6U3A+RQ4fxv4ZIZN6tsxI7r2olE6P9t0olW+KahAIw
Zxe92sqi9j7oyQci2LSbvfUydIKmCvMbPzrn7QPDtTgc/y0rwPzDZwGEyXZ1nakp
B+59kLGl56hb/oCQMWBnCrY01ofHqpT10aLq4HTwsMA4k8OT9naUixePL0kSeNYF
H9bktpB1bv+ucQSRqrqmERMFZH24qrHnUXJ3csGIOoShZwFiOBnPBcKGH//ymPoJ
cpLPMTfevXfsQVa6Nd8cL/bExhMeOZKqvK1rpbHkF5t0HpqDc6cOldDmi/jHiAAS
LoK8CmlmpO+m2scWaqooj6ZFuaFQXBmhwV5IRg70lttmEkY3OGEtbczDCMODUoeH
HlvTTyznT/DfK8xmAI35aO97/kfHxtSoFjiudS/fEzA2AeVXS/tqZV6iz5pUhBIg
diGGSFKw7CyNsbCyx/60m89J24+vpVibQ6h3p99gCr1fXmLpYbBbOtlW8MyzPPlV
Llseab8TpkTBlJUOPVE72XOdAJTdNf8zVPF60EWL4D1XUObD/4VP2My40xW7zi2z
ZC8hXz+FpPKJwck/nfK2FU3NoI/m8MbG5/QAvSttn6kkpaFuiX+rsKIWwGveR8wr
gP40Kz33+9Iz4s6orWfQ4mVfGo5MZb66f9BMjgVaGD8zQwo9mZXtJtk2nph/UPlj
T5Od/tbGMvFa6TDtBJcjly6XhR086hkYcGdFe3fQZFr8D+m58xz9GBQtYj7fFfTs
ZhPAM3iTybtPHNBCBT3mIUpd/Zlxn/2cTFQc035vWZV51bLo6Pg5q3i9Ma14YctO
QxF0S7X7uFzFjZg9A0BBD20qS++Z+IeeAw/5T1CgICAxwnzpEJEwM+OddsDVVI55
CKM6hnY0rw0Koh/dTvDqP5yNdO/Mw72kxo+hjmB1BNu64dxy4B8i+mvUyMxI8QCx
Gq88iejHRZlLrk1o0z1Ysm67p5XC3GElj7ZiUEEuLegSR4NL/aq9ovzEJRXemWoD
FJwO+Rbb1Y2Q9ifxAoZqti5FH7Rxm+ziI4XxjKFSlpm0cpWg4YqPxgn7p+mUA2dL
IqgWkDb92R54eP66TtueG9y625Rq/c9Wy2qagoa7fUq+cjZ9bq66vLF+DfRD7b4t
k/m4qkyGZUOzuVGZBP2N2VFbdedlPmbzpTjBSFlKYbCXd5SPhDQjYt06S3rJft/q
32kD/ONGyR0lYSlcNUE5jiSOp8hBqjvFnOZG9x97WJkGDRUW3LdqL2u26N5zayuT
sa8bzosq1jj+DSgdBidk30DLBdxPYOAVpI+OyObBooD705RPsG6Ztprm72zylqDU
xrGLrMzBEZE6irfvXibk+/ncrllSgBK0M3/+AnWRwbKAfuCc5XJaPRTfQK749kMX
F3PnMSVvBYu89eAIjzLTjctqkw7UeUcZMUn3l1UqDNZoxkbeFQvMgawQvJ7UW3Je
CAoko0LCstWaf2qWvL2ol5gu6/JK3IPhitiy8NjrkLIXHwcz/fJylfwDJZcHC/IC
QYlYR5XsmnY1Tj8a5BkkmtE/gnaRI4K6Xe0zRuV9hVkE/hIBK/NX5q8evwicf+np
TABjJWfHKsSDeaPDDe7D+hjVGk0zOj5pCPI9fE9NIQZzSbVYnb7HuA9ENjdY5RgH
IP/5pJIDDNltlUUn7A05UZmmcowUncVZCvxUNOKcwsclY+w98hdnTGf6W2o05pR0
dhTQDhGzQIaFx66IfSqTcnJ24u77WjsELoCYdOCLVn45If92p6eKKzQV5lOwtmPQ
ypRl/gOnRAszRf5nQ+RQRIFdvWiyyooPZhrC6O518ttxWbbhiEX3xAadOmJKeRwX
P9tvkkUZKG5qcxbD013lP5u8K6MnmDeugx1Um0xw7d0v49pVcg7930d6e9+AED+2
t3IekJFTFl6UhwrlVbc8WvvCuwuZ/70iJ7WlVPGGL8HI+P7Q9daFgxmhb2ST7ddz
lzXlsbD2t/lCj3+19MPH6j1P8XCMd4H7ebpxej7PkQk5FJy3awqG7g21bBB4LdC0
3wM1xu4lmciPBXx6k0nwr1+N45JJktBKNoUA4UbxYUJaTl78Vcg4BHgMk8JIgSTE
I7zasqBywUQ6C4UguG03Mib48SP+WQ31bLSWnIIwZreHkxBvAVfWv2dMgiIXcab3
bcwhWfaRgSUdH9yZL3XGjXt4tjc3qCGoJwrPRM73Mc83y0DyZwKnB0CtS/r3Cnfw
GqQTsy94uAq/pvnyE1sBJI152+qGw5LoFdAofrJbuPIrhifyELpZojL2c3p6Lo3y
O3jNvVmFCrSU8YJM/vt8Whb0VZM0XdfJDgCxMobtw5DRzF/6Jsq6odVwtaU2WjJf
Rue31LB7nY1psaASG+7ysQWUs81ZGxF/Rp7bmwm4C9Gj1vFfebeCX0mf64kIzZrn
noLaBnRPl2XapnE8BwzHwsZpU7apxFHMRxi3/YCc52kVipZOCXsSSEUSZNq7gPq0
KjHeeQIm1jAE1X3uCfMU362UEQmkhOAFHZtXNxHvSbHu9iiROYZMDyYTQ90s97ws
a93xe0spl8Qw4Pb+nWcsFr0atx31UYtld29qlZiNAosdM/YghpaFHyQfhsMjhM8T
eCc2WLGXpOKmLK5h6NCTuKKOA6M0w1pTFmNm6irNFLjCkMeBp9oeVJQwhSEMuP/X
1mXaN+1iZPjg6FPcFcttZsJ1E6ED4NtLPaRwmCbxOGE2uxLaFR3sXBG+G8DoRIQ1
8hpKdoBriu9WrUawRrtkBwwsFy4QJ49Osr85WaPPNTL92cON9naYJa+zkm+q+ExG
YmY/3bxCzmn1/MJ9/OP24q51x+hIX1GlQhWZt8GCqyiKi54WkeC92EX6UEnzwtZu
yxKT/zp2wImGIinE1TMrcx8+JghnGeyJJfMC7qFqxtyXxqIHS88WCyqjcbqHvIuj
59MrQpLMc98UHW431WlUEmbVyzzT+sd4WQEJZsWfkVQ84s771mYxjc2CDMIQRZ7y
bW4JbenB+wxifHh7Bkgvt+KOgZBVeUP1gU04Ah2U3sZliFlBFv1ox8ixTYVSWJet
eXHft3ogKRa2VqBKOV2ZLll6gmuxnyDvHAcWOlu1fTEQPUU8Q1pnrEBWTYCIkdsN
K5v4Rf3p3h/AuUMhZAnv7J4qhTOxUia++wwwvnEnimU9g4tIO+WSc/RcXpqNYhvO
I+m0jZksiw8wQVMz7gyIsX1igURP6EsTFMawklyzl31+igKKDXJaCmF0v/3Z6wK+
QSA1GHLt+VkRyatzULcCDMjCJ/tY2317Aj5dW4YYo6oPLOyBQJwLcyTlBQNApZ8R
63E/AauX04Oh7Ng7wFGyG+MQP6nnC6rQyNaSooQV+IXOt2mCzeuvRUQ8v3y6g3hE
INbZeAQ8nHTId2IFAWDrWR+ELnedGOShcYXVQHMrnfUOrzyUiHX38/G6q4uG6KUl
LvLn1Af9M1RPUz+12Z5qclyD5NZ45hORZgHLHpUr+YdqeipQDbDZxVFuyFJIrCiO
0UnR5tiOaUvA1b+vr7Go4ZeejSF5krYPXRm+vMhYdPb9+g8Ak4z7e1yO5iC8eOtd
aSXMnZ3c7gBC4/T3bZ9d2kQZymFh6AvosHIBC9MU2Yw8ymJGFGvbjbSsBuYqKdOK
h//+r4c4jWpuj7pv8hKLSbH9gfmbASLfbj9cLuCCmZ/7DYUMzzwvyYtaANiQ56p5
KbqK6uUhJVg9iKzPBqBcE06LGgAy63B1gLfN1CYaufVwDKSUZCMlpX6Sed5g9owQ
PKV87AAmr6Ii6zJJUYiuisELr+QKkNISJ014ryJie39QKQMtuFbbmoOFd1Py3UK0
Sfaa6/5ERKd55frwPqOhiRb52wF31Dgldfpm5zbvBxxxa28XaGJxXLFjjVFCEK01
q0Fes0v3opGlFbPltmB1sGgFDAepbM2DG1EGWQbUVcfC5fZD/TsLFkoVOrm+wKKp
KU07MvFxsw8Z3CPv9jIcK95VfJryEnMCe9wzf9nU6v0NNelQnAbeMASdloA0lldZ
rphh1Ie8KhTRJ+yPtwdPP5ar2Y1bJDH6JiOZWP5gXwsryGlw+4HB2r/Mn1jz4NEr
AUysGVtsgcSbxI19SVGkRXyohVEbUDspcGYVfe2iYpkF7tZPmqIwJZCZcQcykSro
qXzudwFHlbJ7iwT65meBxpw0xSbj4yJCTCiX8v6vjzfsE+wegSKsAT4oUrsLFEVR
iKd6U3CtF+E6yoUEIeRQ9b4qaqWOU7VE22Qp3/SnXfG+9kx0DyAtZcQTvb04V7MM
k0O2R8m1u1wg/JRKpHFJZNEAG5ju3JsDR6UqWcZBIZyrOKdn5eWlEn2M+I5ezFal
DbflobQ7v/OlrZj5AhExHiL/NGFNGt/zStNMbfHeT60VD9aAlqzuvBR1ikytoeB1
NV/k6XDpwOZh/rEBP6Tfl3a6EdOvUZkFK2/tSW9uaf+14kgs/OQwQH/JSbVzixuO
lQdn4j6jN/AXFsTckA0vfDaQ7wX5cG3NbrZv68sLnZVbzqOXqbmGjJtiV+60SPVG
ayUkrHDRR1rzKIH8lse5a/XkMRajdRRw9kp8qrYNEV0crdyADDOG3Jjh5xWRiDoH
YzhYJkonKu0z+GrRWemxZfaq2tS0+ZZBTTdC1i4NTV9a5cKfL8nHFqvyUEwpsy/5
SMGm09iMGfNWvdv8pMtN8/aG49bh67TVodLjzYE79hR4eb6/z6SMf2QxVWi5emDM
eLxBx6+8O5lffIg5S72gfN6rCd6vYO2kN/DMLJCPXXM+O9jG4UN1pN1bHrr1Xd5l
bBdlS4Fyyu/yP4hgfcxLdcOSPeKddMcp2Q5h2bfOFyOgg0huajGLswmKXSU+v7lF
Rpq/UG/gIaatEZDIGHhjiK9qksDihKcWctEiZDv0egD6QefnCT6logvZmu8r4Wli
dopa3DeeT/TbY0VE5h67UqdPj3MWzH3EA7/yEGWza6l9HJZ0kjRW9xl93TCzl7bd
XRPk1s/FAZhpQVUUzL6eyRVhHjkfvB1AjVHhDguDrYvW7PHmPZSG1gsxNQf/ueCt
if3DPRWR6IFNn5SbXi/fD3wTrlz6vs1Ep0FmmtYUOjzwgwRQQ+Y/yr7SSyrtye/s
nD6Giwpfk2oimIZsCt132iYIF1cG4eES3mYLuNxKS9GrVpr+Cx3YlXv9Re98ZEDO
saMuleNP4r5xMrCeAJTWtPiphCNDvAi0PtfnoW6Q4fVYFhN5/THrtPTYgGnr7jYp
xEJdBV5+2PWzpM9FeUQwFCEgNi2ycj89WQ7K7d7py6puD2OgPmjLwyPq32jM7gEd
EhIQw72zLBiBvWEUwlXBhLg2MrcF/OCg9BqOQnqhy7bzP3LzeSBonOT+OA6zuaP3
PuWPspAJIwYh/24uZLXNOh8iFVdtq+3s1xfGzODNjSwHnOeWL41vYKyiKQuMUemV
eGhBVQh/RQ5AWvUfCmbEQdOYwgMv1KUudmLm49Q3vMkr3kR5/8yjiBizc3QIiVes
4NfOc4xU4vGs5Q67XtYpsEWvaBy5XlSco6TeGdOgukvN5hUzdQ1mFwc8SK62260Z
xo7AvjFHA950quBoMNdKtFq5+ycCR8hbSgnEwyMPpGGXj2QXo7G1CGQ5wNd2jjqX
eVQfIG7eNsw5fszXe7wKakX6ZAkB17S5wOpjhDC2zdULlXhP6PohH8LU7pHUISot
w3NGIuPCAkhWE6CxryAvkBScS/HFU36hdCeWIau6dfFGXoNaIPu4X339o/DFqfO/
3aNrL8FyozyMDwJkBLcFUeJnN0/BHrX8HscvyXwllzijyBflJ7dXzbhBv+nZYikS
rPygMsZSreAcMdaaBw+iaPajW/sfkfnPcQ9DyvWopcnym3WOlRXJ+WPbI8U28Exr
FN3oXZxvQ8ThLYCaZNT1o/sY1DvPH4LTbqHXfsQo1cJm5uWqcuSuiT+g84s1dxc3
Vbc80V2lX2smDrejucXJTTIcRaYyK862krMc5jjTk1SfSYmB3mTI+ytURD9Uz3Al
TMokBMgh//jVIudOmNn+cTIQrTWj1R+F+PmNFQOXfZjT9zVP1D6qx7SjPUyAEo9i
HiYxK7tqZgTNVsqND0fCaPPl22EntzF2Wp42n8rQ7ip/brk3Z1FRhACqNZvwGFiA
9pzSAJcEQjmT+L/XR40A2L+KcusrX77izEjN0B51kYgy+ypVDrJTt0aDMzl0TxH6
sYtQ4MOV/+DUWg3vzJPY885XnAVuGFON1L3/LmWBL+dY9IwuaHc33FL6JPRlkvG5
dpuAhssyQoamvn9Cy47JGRnftSJxZauV+8X0HFeZzmyQ+dN7k1JzUZnyFKv5mXc7
P1y85x/U+8ucU4eof/6h0cxgdN3M2eBZX4WYLoFqNaWvDmLNAuTseY23YkKNqFyr
+BmTNBWVi2sUSLahPBWJtRJi687aaD101HDaRwkIk6fV8CumcMuqnrTI1mHUw6W5
6eFGSy/aeL3mf//iEARzLdKCdBgjGKdvvHj/3KIxAH7fqo4Z2fTTHOiZ/7T51qUN
xjE6nv5ijnfNQP98zfZIlgQAkXVV+/YOTSDxNShaI17wyy5f8aYDP5PWE4+ymFwz
rLe8H9X4vamtBXDEWLwJYxFQP2w/Uw70kSxfxANxevJ72FP4OYTOAcIXZfx/83mz
k0UbzUHXTSAC0xQtpknMPT5uOeWFAT9VfTllgHE1+yk/5pGmQFSW4jaG60XE2Tud
+JpFTmQAIsXUb8AyeTDeUDnCcDmVz88FhklC2mMYUomcHoZj1Np9quLzMAmOEq10
joRaljX+quVidapo00UdaUud9jmXw67FXSUA45/H6l5UwOMpSWEZoGiZBiSNGHRi
ybx4NDxFUJ2W3J4meW11p2dwmelSOjsFvlVDSi4ufuTCDIEtsZSQR1mK58ypxBdC
pI/jRFIyYIZM8OTNgjbLi07/pD1W9rFXF2A4SWOxzD1DLS5AlmVvjSxC11ePm8DG
lnbHWBGqqQs7d6x46p9qA7PqnP8iYUzJTNAt4+9nfg0Fydf0WQDrxeuCmQCwGBwP
bTozASte7vp2trAli0JkusfHU2ShpGmbt3O3IDnbi12cQ+YQnOk1eiEsV9pp39/u
W7BR1ietmgV/ijb6TsGizkGLiBHvndt5wEY3WPETZD0rM1KMni04qN0QREz/QMsE
O5HydY9EPrZQrzV2waLoMxv6fySwmKo0LOiOYs1Eu03pj2yanu2pME67u/BMm3P4
TdxN+x6Doi/nszM2JIHO47Gi7h71OI03bQ9p6Kt4n40KhnuB5ez/H/PjbunN3A9I
BxPG/58oIB6FfckXYUE5sQ7cIGsXgwjOo2ohjMN02Ro/43JlremN7+BemZBz/XfP
LarA2nVIrI3gsnLK2mEAs2VNVwUcCTcd1a3t1fMPaT9FmCP6cudq8cPyzaNaoW+B
a5dNm94dZaHy+M4511al/07JjX25HjOarIC7eIHpQiwu1TAToLMfFocJeqAXLJBu
H+XQTHy57Li0r7UlH54Owlh0jArOSgHCK1bxbRelWvtTTupn8tqdTCb7u9kaEDJ/
XEf8NV4YiqbJNfVrD/6UM8BceNYsS2G4V8aJxWF+sLGLGDD2a8Mqf2+KyaMauvIQ
+Vg+0LouE1/lnDxBMgAw/AVM1dYB7jOkGADfI7TtaBUU/txFRN8qJtYsuQQNDUdG
C7nyQ7WNDMALb4mt6vSPsej+GXdgTAY2PNZwWYDNRY270nm8tYW241S6Bgk19ES1
5Djqjn50p2rwlHnyf3QXF/f5BCxOxnqCZ+C2psI4SriULfu8Dwk3Y3f+0K1mKf/Q
FUhCCAFxSPFUbcHxB+iCig9hqSFjy5g11+Mpy74ZD/nYrz9Xi93QIJGC5lnKHWvX
wOxB6uyJM/Ds3Ohy1mj5HbtVON7Ck173hFm49f/6wyVMLWO2CBEFSlcAGrk2Swpb
jwfoSkos8hu6mvtcAWSIXz977lMbqVLVpSOhk2aAmOGGowGYOxrCpwkH81ykGKY3
0tZWeYomAbiB6gfFjBVTltThzZOMJnArjguUEEWDlBRl7q1FIk3Wlv5sM9xI+PBJ
ImLKwmG49YyVQ6scNQziz50Yw/VDsuOd3wGiKT1p+opi1xQWgxjT17jBzPx40nSi
GjrOT+Mj5ktTtF1VGFAVLbloHEcTl4iC1EpFUz+VX5VThHvf40JpjxNk8ufXMoPh
EzodJzoYyyzyKc7jlm2v8+p+cA7T0z3ObJEHjlkHJV1aGpT88RAUgQadIuDxo9FI
eiSbWEfz+oerARjoB8eU/jUoYRC8Sp/au0qeuVRDyYdgySVVtY7kIoMby/WKoI8z
my6T8GKIdo+6+a44Qriop6xt49nGInMMa3oukJXykzahzZLOi0qyL9dXbjkzw0WD
DG5Izt7kwMbwPq9TL4xF2Wk66u8l+10LRqUIwmJ5BwXxMOCV6+jC0yhZHPxL6OJS
dt0r2r74GMe3ZmyImu4guxq1xOzTNUj3wqPv2bPkblaZOF2JfbPCWwvhrJGy+0yk
gS4ySB8y2q+zqpH3Xow6tTx16S3xHupzxAtlGtBupuItr2g8q/ZV4vUo3Czp6g32
QvzPO/lsvPwf26W76O2VXLDX8NcuNMEtPdNvp923oLzKYL1X998ccDNyaaRm2Usd
h1+IWjT17blNkDitq2GI5v2gDG3pspZk9mzkwMsLMYPSmGSI/tXU+jV0WYxn7MBq
GUPUr9t+/3dgj0i3RKffMneGZHBR1IjmVOpYXFCoolajaH/Xz3gPHJtkQEMZgEW1
pswZtbxb80ActKyRdUzqz0x/vVyXvgpngbMzwarCYl0lYKx4OqEvWxjqpFvRv9ra
9J0gP5tRBV7U+MhVNEbM0EGhw8P9qoNLLhkYXLBepK7MMMxLuG4HVqV8j7KqXxu3
dizov47oYD9VkSO0cwbWYFAabK6FG1dglAOKCx5eb3du5t7TRyZCYXsQ2+eer/z7
LF6+K89pwIzJb/rYZ5A6osTnBpZYyUebOn4W2YcbskP6btkOEUp3QVrgH+gy8iQj
2nNJWd5JyM8t/TEaOIVCeLYNbwwnVEb6Z6IQSUgxO9KQQONoar4mhp/ZWoDG73dn
4wuxmafmplyY5rC1f2X6w6nio0YSqn3+Wao1w77uKODc0g1ISpTrZF2bjga2hOEq
XPDwoKIZJOfdqxftgwDavN5ptOqCgGTlQ2pHadXIG/4AxtXgd6ybTgBgqlvLYDdW
pJBYNLLYvWvaOPcUL7at94aReIxQC9YtoO3bRhzii5r0ShvMrOJfWGz9loZCC76B
uz1ONCwprBUmMzphchDHB2gQY+NIjSWx0NIBElX9ZmlH8Awy22gysDS7bieINhLt
oiBKGvEwqiDcoXqMDeGMwSUzFM1NT9NmuKS1hpTCamjkNN18lMJ/6A/za/g9KRn1
gCR0UtJ8EyGiNdNJnG3hG1CH1b9lt1ybhxrorl1yzG0AhXDDp42DcBl6H7zfGNU+
XQcuRNAD6yqB4mgEEg1JA844W+ALDgJ9RCoJn+15rbYWOsm+HOThV5670lOGHj3M
nCu7RFeAkNm9bf3847ND6/65d/o63aj8yZ/X3YQ2n7OgkgW8iNWak6ScClCG7imU
4xbLLuB+/5Wh5g+t62nNVvqXRNBLWruhHrb6B5WpCkG9m6Kx8dcPT7VAghvWk7Vl
OUL7oCJEDwxuUo8pEf+66vo8JyjYOvdTlYfLMRO1QKhGknbV1F743kEFmm3njzys
loICSb4iKglnUY46JQjkKQXxSyyLi2jgHPs9fxlgsOaeqC/AfHCtRNttbsD+MGjU
E9776Dhe9kVWBHVhQcUWokib0B7OPrGmNMC81W+j0AnK/rdiR2M6cthHOvwCJMXS
kebgTvDTMSxVYFv8l2IWukC6QGpDvnUO1zyEW2IRIhi/l9pnL5RmAUKorMm/kr/E
5fIfGr+NaD1B4+gv1lz+6LjCt6Eb1n2P13FsIwbzvPFDwIdigmiaJcR81qPsY5Ex
yH0auU4s//dLsmiTuiKeHFs5S8ynDOpWYDAnQvtn1G/7J7ZrD6OP2CM7EzeTN0/3
Nh2SjBvMEG5Ybyn5LB89eWQZkL6YYOCLeL8u5ZKx3EJhbDAgkounZWDtnWBpFTQ/
IgJMaYLXXUSn6SVR0YHrEBiboU7D7bMwvrt8lehIRX0GWl0rRZ8mT5nOxuy+xPaU
qXH7hlxkyaRCARcvx/ox6BYpMCND+W2c+htFuyTTa7N5SzcUz4EG591+0ylMlsuH
jEImYKJtE+zeRe2qghCvjPSeQ6OaGr5zwyLcnkAG34hQ/Drg5baAGZVZzSer3Hl5
I1cRQ8yp6Gy3XjVw7r5A205+O7XEzv6zZShHqLmJPtE1yr0rfi65TZT+NWGYFLy8
LMk9qE5bw+Lset6bzLJjJoUkp6XilK2zFBN/UmFkQP+3nWY/zI6cufyDQ4UcV3NB
LS8nOF0USAyr2DBqCBHJS4ygi5Ri3mzNEabs0xlwNsaYTGI3jxdHoQ/kks4pZND9
6s9Kmt0IZsOLDuYZwd72j3qyIn7HL78PP4DkNNPi2sqTj5FFPvrjHDoeRjBYicz5
Pr/yUD+ttqOcnrZ5xE9SLeBxajGx0G9gT1LfdPNgnbq4gGot3xaf1WYHW+YQkLmD
PDgTZTBMIQBh8yHRAAW9fQHGiDy1TPHEmGm4qB4GDa7ItRbbR3NHrL9LelPlQieu
yqoN/y/KUgQVuXfJ5q9woFMs0CYoA6zEf/Aa/Ub/Jb2L1Z6xkNn5XPBcWSRLpXPI
xi5jMCtCiHdZvgHPFH4JolB5bd+sR+i3bQndsVIIoo7ij0zf763uQ9HhHF7usFhX
OrumbGf7mqyDG4t21L4sE+nMmpf1+YHFy62Ic1ZfU/RJenECTLCR2Zjmpm9gHQn9
Fp4FJinSHzX2pobf0y19kb6041fAFGokRHjCgNXPgrMJDX+DMFknzFjn6Tuq2Od5
PxON1wXv5tYTox6iSUreDOoHkvDNS2QaFCcU9h3EXT3qt00w7v8ippt1nwXpXFWH
NtU8dtiVSMnpAzi0L3RWkIez+Ek6SHOvlcVrs24HDhAa1F8/9FEJXqo0rGsJRDzD
9KeitEv2fjvOrxPgKFp4Uub6droJXzQP2yTept3qZ29ZFpzZkYQLH84TrK8URTNJ
TkNfvbgDcgU/aQGyeKZodjMF0JSMu46kGuMGdWxRD8we9qruxPZAxLiwz2zGgNMb
PQzpTcTuErseuqU4SmZiLq00kipWNUCLco9fYOA3VF8IBoIZByTYA+/4Urr716BP
mJPhC2suetihH2cZY6aVkT2gsJzQfWhXVaxpufzUEXEvuMsi/7gx4yOT3vI1dJDW
/p+kQvrmAvVspWJW65b4badBfZQJjA6nQ9eA7ydXd7rE7NgJpMXqO+SfHsPV5KrR
d3MvSBXXMxLH27ZdBaRA0YxfroBJ9Iq6ZR2ZmG/uYYsor1qPIqlkblkK8pIuPVYZ
yZyvFHMaFDTmamSZQr6/8pLODoplkMSEwoWrFMjx3XuIZ3Z1HoC301/JYFsRDkrY
drKCMe+EIJS+yy6qqKIOkcRr8vjRbHO5BZAsAE4/mNq+Y85D62Jk+aRtPDHd5pvQ
z3juRE3RJiqAjReQehlSeFE0sy6jCO6tvNSOJFqpxcCRnojYlFPw6Qh0T56NJ4wo
nuBFksX0beM16g12mCmy92X038woBFbZA/eYKqH1ABCNyomILwE4rk3R5+lZ1sCK
DL7QPhfzhm+CX4YIJRXUnRQiMqHzas5xG0Bvl8qFHpgIQgzfrkHHXt7F0hfqUezl
r3C9rs0eYAFu6AdF5j+dI2RBUgfSYSl7IliQW4lCn5lQN99oBKTLGHI+FbVygh1G
+s2YIJ9Gs9lX1qUghKTjmEtR1BGuT5HdWiFui1/wWtxJi6VawXFwKzcphmLFDu30
IZ2i6xBKXYk8viWjKSqdPHD4zBWE6KWBqnovttNmaMFyOv3rSFS4PoAxdI/Hk1NH
oe72o85bEgpJBrUiKDfeUBWTqQAu731Wal6/2GArOQD8IIka/fHr9Zhlp7Bxd2xB
Eh3+G8rtB5qrgzGNPX46VLdcphSoRXSY1Emt1Kjg4HF7ZyWVD2PNwYjvTj5FQIeT
N7/3PFxW8mpApCyGV9L3l9EUL1TYeckwnf7HsH77kHfxfpUmyWLW3KGo0+b+dhX1
6uJ3z8b+SreLsvW58jQz+0NFZGmafbfd42nhTXjFZXAxh3gusJP8NwHXN+AtsEIK
JnDW8htTbnFNnkO8h5e/Pigl0QumKXq3KxlI7pVt+XXX11hhnvYnJjrGz08Tvb5t
cdReYCY/A8P5mGgJPC80khGsnAYtntoYYCui6w8VmMS89ZbpQkJ42HzJirBzJb7C
9u3VlsehO5oldvfK9p707Y6zS+EdPeBqG2ePQ2o/b6NaEsdKb5S0qwIDSPnie0DA
zCaiQb0icIQVFeChixKyT4VNe4Y2qdZl3RdcqrXHOgbQiaBDh74KkkiiijoR4BQc
66pvttZonJcvRO1uhDtd43YwvC8YuCxuUSmOCT4B+di6JysNeCO54jujyw4Mxc+f
KsghTBTEethmHM7g0/fg+aqWY/eqDcrxDcfEM12Bi7iUzbEceBUJwqA86K6QbPNo
CgfuececVwof4N6GZFWp5B1+64QEKOHy9WLGTXvL4emTd/7LCm8I7ktUx89DmPDh
xplnhLhHk8+xHSTP27ITvwslpCZa5iXLnHIl3bUn34WdX3u1t38xu3k+ifKSyNor
c9UekaB9dZaQR//zo5TI1cfuy5g4LgGSDaeQHTj+vCzkRncd1b6owBOIsNEfVZCJ
RvzCov2HDM+lH7zAAml1aTvudMV05XWeD2ZWBUX/iJTYTh5Cgztp0s0mFE9AqecB
sEW3pCvi5CoRsJh4V424VDMNY6v3Sp3aHjoWyMzq94t/D/ytXm8iJ1//yYKD1JAv
kBd/Uwf9PID1+SSd041jRBKkCdl5JngLfzTupqKMSMxHixCtQI4AOSPE2gyslK7w
qfAWFUI95auRL5w9mBTjKd28A6Die8XazGn8n7p8BiEDS8DpEhLKQafQEf7k6tVQ
6ZV7lUPhKByKj1ibRPzc14hnO6gCH4unbpBqo+/oTFn7VDQPJleHmbet5Lszhd08
nvCju2eiuoJGux4lAOIZLGUQ6+55jzgJRMm97v56zmcV5jmnu8HXPicihrcrVYuo
sdhxPIxC633bWnIvZ4SXII0GsCf3znFGRKezMscMv0JkMlgjidqw/+E+JiCturA8
sAK5jxXtnW5jmbmBqcMz7N/o7IT31rmKw1hQs/9LslzrHdxA08OwfVY2Q72nVff2
VRY9HznynrSHZCqZ9UZ33MII/LGMyG2Z4ZoOEt++/So/pr5HaDmLTO/iIl8dnK5p
BUq2PwJspAZ9JSeuLl7uwTIydpqQXbV71cN4nzRARz/d4jYk6sRlqcqoSu7ti/0g
6eD2iCzi3oMvuYZEqsXtazxBVRc9l6BiEBSHHOjV5VoG1jPgyLSuH4WQf1yAd+bQ
G3bGIHz7sJCQtA8ImwIl8NkEJtSebrICC9/5Jl4vTFgqbPI+k3yamF0Ypp1Yo9Jw
X2vEzTwqQJ4moJXMziv21T24TBYeqBPijFdg39XiP4T7Qt/fTnZN1M+q8BLqkyAa
JS1N2z5hmDVLuoKjjmu9fhh0OiUDt4x7ofQBxrGgjTmqcVvu2CTMd3+YPhqLoRm+
cs3dy66apAzE80Oyf3I3gQlSZIpe3ZJGqBPeqNLvtmJH/fXar7WK9oADsxV9n2x9
dTXPSRulp9zsqlyQasmBK2Gt+yilRp1HitrjlKh5KftpC8P0u1XrELvnSiHQt3xT
p8xXk3G0hbEsU9lQoZif/a+F0KIxOq73vCHFNdWgsjEbrR+3wWNNqomwtIcQsx2N
VxSnypID6nHkZS4ufztv4udM3cExjEZHhr0UZBfJ2MegPNqYcqj9I6r+yrXO2Avu
QysYz649Ptr3W1OQhwbxv+dddKVMZUE2EWjE7ANRml9bNGHXcrgluwU6pejhCP7m
S5TCHe1vkxjZg92iNbJZ660GosQRZlgG9WASuovLH9lctwHriOMofioHoaOIoSm8
NI9L8gPsYypq0Mzrjt2YDboGtmuirGgDI0Hm4IfRefVRNPm8ildFXFL8DoYozgPh
D4GKfoGPnTYp3PiNF3mQd1yJ9BAm5YkWpdeTxrx1g+k/LPWU8/CP7sC4/cRrxvyX
WcT5Ax783MpZ9TrsaP0d+eas7bTXuSqUqY8Dbbia/FipiEXoGrtBdzj7neojlIMh
TF/Br4UpCdFi7hrgvV44jSEKahef0SLkEAsEII0Qc7PEusY+qn1xu9sglqXajH3j
FWs1KrWm+pllPXRKOQg6xYB0eCg9pZtH3QgWc4uC5GnWoi6kCTy3KIfloepXXg7g
CfXX7mt6w8ZsUDeT5jG4Ht2O5lw73z2PcF1wtScqeaHmdGPR3EddX0mh087RsT8/
vaD5Ehb0r8JkNv385ZNh1zQByKczga3hM512ZA//nn6Gb700Zoy58KlG4Z03uS7F
vEGgZ0OKXoMc6vJuoLJwDOWPWZQBxYNp1+0t/WTWbj+z8Spkb82S5HQnczPfBe46
NnBcRw10Xs+mJhd7XdGx8s12qsg8rPfu5V0dLJI1jno2pnoa9UZFRs8SvsGUGw9D
7c4Ni13kWsSFGVKJb9vBBo7hSVGbnEAsbGysHBxbMDfhgGRrIb85utrX++IPn2MM
8IrDz1AXBSnmkhob40RYo1Wn3G3DXtHttMPcotGpWvEpWTDfHDb/OHuL3S69fI4+
meRL0qtAfc6klYYcmQldKWtPSRAgCS+VrE0Vho9DBOVnO/nZP4+djP7pw7KCQk9B
ufu+jkonEz2m8Dj7mFTbHeivOpnK0R+A2ekufEMwoNqKuMvbDuNCp0tgA2q8HtAI
42VFRdaywMUcdX4tIf/Xe73YbytaDiDeiGapSovfoT4LaheG709MKCRW0vcX3vKX
HJf31Qdr/crnE4QT+9e0T0SEn4IFcZ16mt7X2VQz/Ryo6k9/9yahd08jpo7PO4I0
UILxYcreXJQIRMtNxLE8cIlFerbhkBPrzIhsMDVMY56HqRysan8v41QR4Tb3nDqM
GrsIBHirDVxatvoKx4Azn1O5FAPBgc6hUlSmt68DWSZVAyY9x2e1q1zSNonYQvam
zu7IgAWd+di2wrvA+77Uk59LxzDI5aGSUUW9adJxOFCUlHHX5lHZThRf9nWxjpsd
mUhFPlGm2RJ0BF7a0zdknaqna98VkxmwXd/oWCNvXcwRrmyyN+hpJ+aUJfooNi0E
oHgwvolCc3JNM3eBiPN8bYxo6T8hFQYN4JSs1FOc2ASMC9vQz+IxrWy7TLHRd7uA
KzkpwwYj1yZbIsIFvE+6RPuKRvMF0aU/+db5jLcEMT34beTtNWih8yzHDrSYPJBg
NyMQiyMIBsGA3G9e2Fd+mA35ed1MHvJaf3hjPYjrgsfqNOXagITuYdGg3E3UfTGP
zVh7gdkSA9amcygEYf4laYdUav9gfeTzG4j0S+mWIzPyhXoA6uF0pXBvwrdvvLYH
peOcSfV9pclIptCObS7eXEqTljh+NtLeudZTZsn+Ge8PykgjVXiH4jQibeBcdDlF
wvvihzhL/PeOUaJeahAIliQUI4658b9FhphB5IPnYbna1D9V/1ALYtPskTQz7QMa
VtAvSg8VIRGLpo56Bl4udcexvBTH4H1m+Wh2EyxecJ+iSoYKSRp4pXLF3dH8oszP
FD544EiC+v/ZemP8BF/rC/50ZBfbxdGQNCQEL9wBWVwtU38pm5xReKD0cdqMpK6j
10OrcUnQ82W4GRog3FqP/NXgJivJi0+3YLcx2WNdHVI5Cqm6gebLb09+POqN+W1r
7VJpAwTJ4fp63aEbbqruMps+nge4XQo8atysYi9+k1Tlrmbx2JkObu7FqmoH8fAq
/icCBWArDBJbwLcEYppBB5c0AKpJPUgdEGH5HDVHW33MGDtFfUngezZj5td1P4xx
7vGQlfY2rSvPAUd5FZPEoIJtUdKe9n4Q8Lg2YJxxdGyy4ngCHZfhBR7nsXeTjalp
TsYZrV732cb4mOf6WjFNFvmqNNgtM8cFy3KH6p8IqaUXoKDO2hE44fC5AiiJKrWM
kgeFFMn4JfzgNrg5hqvdE+19FNzooNfxEsUtK24GRZ4+Q8AYZoKIuWZz9pVVMZNo
LEjnnHH2fFpRCh98UJ06Rv2xM/siZuX7AXKO19vJqcIWJqDdolbkbrJ0sk4XmeEi
erTbxjUGPGY6KAXKROq7UOc7n2wz/Y2n3LDA7bBQbowfnLTSYnrhUlwRsV7lO9bq
tmQxeHF1PxHFnxd78eCT+ZoL2Ed1l5gBUwgSKEYAkhBDaFFu7HmfPcjW1tLKwYcA
74Nnm4Jkean5q/wRWW+uuwTnyhwTZPl4sBOGIqvMG/rmbanHi9+KcSlJgspY9okW
A1P/E3aBnWXEocJk4khMvCvzkjYEw+Ry/3psKb9bHIACV5zOvE0PhmM5e1qG4iO0
yYx8DpWzcb2U6RG3EZbTIWZ/PRpo4Qz+dWa4aKGzuab+w3kDA/aOvVokzOFElT9O
x5aBs/9JhhyB8jGFfxUynq3RchRQ3JGZjj5tV309MSTx/icrEgm2ZU/Uvol+sBfa
98/Z5sYywYgaP7r7kw40+JrKI57G5iKeW/Mi1nl/n0Kw5aheDEdCAFXuViCWO2+H
giDy3xlADIGo0c+SkKWjCIP+S/22T72KFsbqwvcQJ/cIpP10o/Huqt0eiIY/Lub1
XwovvGv2oSh8HprL2nAKzKUrO+egoM3Eq4E8oeIsRe3TQGpWtXcwF72TU7uqwWFm
wqdysr1kekywiPR4GgQL5GFWlPFdrQDVb8lUnw9UAC9JpyHLQeMJ15irOmOSke6x
vQIaOj1ZB1jQ7mu7ABXmz2BX1Yhb0xY3OizLPV6ZEbuWJQaVrdhxGWFkSCeVg8yL
G1nCUu8arvZFYWU0/0QHTY0iyxjLBQrpyvKT+9iVbsLLqhrcB9YqTnzWd/FQoVfY
Ch3hZlvpWixYoYPWhGg9FKIK87UixV3iJzEFXu4YEhuD3QpkDRVOkxbM8vM/9voP
QeeTARtpx78XXhJLDYcHpWn+9gmy+kDn/osfik2J1r8iTP0F81zN1xUVnh6nW8GP
7nU5UvMZ0qTxGY+Q9kD7I6clDuZiPpaE6gmlZQwDL1GItcQQ20AjgSPGLKCnahIn
CF/6XyEcDWC+tO+GM7+RDV55r2aPy0Jd7lke8ow/2EcoV6EtV+SHt6wvRdq6NU1K
ImjRPa4P6xEx+r06zWBozIhoZ019LBQ847pqih/ge+CimB76qCZpDWq8J0cmpeZo
TbK2T/DfcuhSxj/syo9FCe5R5ZNPtH0t2giQoXyyN9Xx7zNVrd4Dt9lsnF/yIZD9
Mpc5L4aOEKFVEzd26yZgCLZD50/oOL1PXHQObgmI3XuXZZdKH+6rJijF6iJM/Gbg
bw5jqnyOp2X5UR8STa9aPhfRm4qL47ra74yIcEn+I9ec9kNgbqdXvV5o06FTsk5o
27Dpm0ltxNAswEXtqpuFtNbzeI5SFW3mbhndcI54Mxo61bv046qfjngiMfhVy85N
Uebc/Y4JrfEMtRDtTFnLwmS51vLhxmKFS+ibdC7jyE+DT/imf/86/zUT+oj+2yTw
YAk88Qpcv34/oF9Pt4N3YsEeMZZd4+g25HRKxlbWHMhjTb+gTsdmlu6rwkFAP6v/
yJiofhsfRiXggKJOAxUcfxLTIyKGscVG0cu7GuPkrLOxqZvMWfyO5T8QTePMlfqG
1OZDMmyRSpyaOJEPjeOxJIopzKeylD6plJzJjUtL9MHQUN9Fgh8IQgg7tv33nGzs
WhBJCDKYoBXELPxhW+RDqwbSsqMJapQ7baBK3PJSqk+au3b1lbzuaSWjEKO/X4NS
PWGkidnN05KuWV+v0TaML305kTgYBoGIxByj2ok7z7gWW/PpI92GvP0MFGqT0G/B
3jYb5BI1KfiEB+1omgaUUXVEIym/ROiW7BZ1puICvyjigVJpgSWbAjNlrIoH+xDo
LMTJVfnVC1ktNymrTODNRetU5nrGVB/iYCh56QAe0XOqtR8E6SCSV3oY9sU5R9kn
jhlghxhKDaaj9Ftbl1at0M1PvELSqzaM5Gdm/tLkaH8gs65weR8l+/vzBuuycoXz
pa92dFACipY2CfPeTEa5cgauFHBx2lKobnnsRszJc2wB6aDRqslCSrnNcaSK+MPm
3pQbPcMnwBfrNMnQYJ9B8SFW0Wniq/uXpUQwpyuYT17Bh/1BzEZn33O3EPfwVwKi
9cgAufSI/a2yx+zIe9Ne+b3XX5tYtUMhiJ9vOi+GyvKSNVVGO1PhS//pKN9F8/OI
1P1RM2w9+P19ZODUm6TwfbT2AeIFOsgISAZ5kTGwslWhQjTY7CxxS20r8DSwomCp
A81exHwrEOlMHx/hniEDUc9UwVLA8ks/8Ef90gZDCsa0pxjt5d2NrnLYs7lwx6Y5
2h5GeKdrOceL8qvC+CrAd+gnnV0dhsNWd/JO8OrdH9bO/X7n2P8be/s40sxhIh4d
yhuzds1RjV5uFUK3CHvbgJAsrzFHzdE9OUplZjukfi4nfNb+F9hhLc6sqfPNAi/8
aIjukqBq8jjmAqeUsdYlTGhhZni/L/cBx8o7d2iuhJh1aKAHqAqif9/+zfTkYzzi
ZYgwkuB9PbcPJF4zmReuAz0sh+j6drXTqTZLs/4abHA6gXJbOEW+/8Hll4l3judy
24JioRh7QxW9jz8mACCRlGZtuArA5OovQGrRhrJU5lGZh6ykeciK7504dpjeDJiq
mMOojIdrUqXOHl+BXD/kCBZpTalaInGj/KTJv1CQMnDwyaPyfv0sQ0i02M2CYkbE
/zrZ70anmWELjUrAlwxBdX9GmC+bg3sZFH1/bD6ghKHT2sY8wI3aqHkYoK7qfyRV
vCncjlXdG/koLmJmWdwAxn3sxMCy6TVDbeQXuDyMiQ6M5wL0rfPK4jerLA3kwcSc
g3tViiB6f8DtEfj+hByXsumJC99SOc58+Tk8Ps85aZKoUG1KGY4RwrxeuSTs6LAw
a5YJ+Pldzq7XGivWkO+3gRn5etl2N5hmsySY+eIjWe1AQCmxXkX6fNCqmYdhZbSY
FcXst2+lRrr7e/L0Sb2LERswY9LHgNw3cfwrcbG96WWH8uo6YO4M2PleMrkU682e
7cy+wMSlsS/qe1qfUXIZkB7RPiBfANslc24XfGHHWg8mv/ektT6f4XOOF5f9Sv2J
fB+sALPzYpGBjaUMw/jW3InwUsX4V50GLgjlrYV09sdRCf3uanFlbtNV69NUO/p7
grbmWJTt6sAyqduqpuhpiOA39iKnow8NuQlz+sguoi5CXIkA+G+/La/wpOsxlnDp
gYcI5jZEvXSIyar5qnGXiOSzw7GQWehuoPguWy2HCK+8qa3nL5WcTrpI1SuSlRL4
VVTgSvsJQR0lDYvts9DXuAZgNjnLGApzQhuUkr92V1vrWBgTN+CnuJqu211jSfFK
1FKxzCxjmoWCQ1azOiX2Lk8G8cBf8aShfirf+Iq2V6ZyWW+gabb61isdSPn4cwXY
4mdTrO0Jh6w/hfd98hTJZZOYP7myP3qLcT/HdN6VjPvhq2O+HZGcQPFao0vi6B8F
aoAIjcITeGqLvHCx0tOFHzdbEOZkCKKvskeUd8Y/Uy2Cjz6Qvu1dcTCVP7UaBV5w
WW1ejB2WDvtNYrLVRaNDgUHl1sK62aSXrGbzt8nFdqjgiU5Wqw5ZbDTIio+907m5
nwCEyzijPSiRQHMbahV4Y0dcILXm6DrWmfHMcGd9wshoxFGNdU3hNsEoB5Q8zobe
o9OrKP8fIiXM9MXO0avu/1Gaw3Ja27bfDZTvd64LZJB6wggJakxRB7wG+8W6lgm4
gYZnamXqIp6UiBq3Nl743Skhn+eQBhr8pXvC7lj2ubyOxdWEGzyvpRmG9hosqMbI
YhaoIu9U5BsNSbdwkxgWR8wm9aw5mJCgGM2UjMIYhm96GqfwpOfEvyIyI/F1kh2Q
dAJy4FVIx+nEQUtA9uKDm+dHUqRm5u/ZFGh6zAQFe3+dJQtwtKZguNtpqiyzVMjz
mkv3nxG2jrSZNGXiYd2sl7iRx5O5PzqKgsUx/n3xSx4Ow7SMWC47gN1tZj3n+U9/
FmTaSJ46VeN1Lz2OwoxCEmKGuO9pgtxzo2cVZRkc2Zj7I/k4TJzbsTzg4PEMRMMM
MTCDGLp/PjPubbyUk1qoQ0CP9SCGy79Z6mkzbb+/dFSjWIsSVZ1Li056+Odmovc4
KSbuDeklJ2xPSMg6A9Oo4Vv/6mKB1ekaeXBIVxEj7B1bhWyslLPdjmNF9gXiPWqK
24C8uoehLbfYm1RjdUuXZHHD+hdw1Hp3jLMCBeu9yZyRNcUDhFtlToMQimGXnRvG
58h3kJcp7MBnKYi0tkOQrh+Ig7wRxhp29ytvEr4spqRFy8M8vdeBn9kxMaSdv3O1
koXp/PczioysRqeQCb0GdGlciy+ovTVmz4nFFhdcEIW1dtZdH+Dhc9wHjNcr6/Pi
qK4WA+Ejcau0b7CCQmGjgdb6+ZJQ8/V7d0JJSia3gcWqhTuIwvXCoNyTqMZkZhrZ
FBp+gGT650LWk15qz6XCEjDU4zgvRJD0eluRdmUFsH2IRVew33FJJhKSKjEhhcI8
r1EzJbL4qxEYnEz+tJtnhmQmvTUtzJeyC2A/+tNX0ZHkb2H5Q5DInU0JwE3P2Z5C
nrGf40vYpbb5n2cN/O58bbIiN1zkHsQRK4xoaEWeNP/vel+yGDB+GwnTGJGgIVE7
mjmxM1qDTFVjTCwoo0SAUiiUKgElulLconoKxtP2TiqHBxo9gBSprvv2le9ZDMs6
69aiY21LyxSNY1QlyX+iwW4333iRaXDbSn0M5VI46yaym5PJWVPAf2rEySe44x99
UYou3vnylWZu21/tF3kUoW0Qqtnm6T+oK9V0dfpkfLVy3iwUVyiwVWmP/RpMJvD2
hwmd0R8p/smx/hAKZT89x70uotnyqd3yY+SWrFvcD7nX90Dn7pGn+4RqGTVDvFWg
Y6N1r+WL6GYRJZw+pd7RSro2gcWuAMtJYaxwNJwTQJwpI4Nsp+dPqEH8SSnI/zpU
HJ41gm5TF61GmUev1IjSGtX9R1VYEwF//4THUubVKTfANoAgEGkhUrEtX+EMVFTq
9VJWBCiYVsRtxMhSYmmaer6gfokBa4N9zJzQw0/F+UKd0JktdTJDWUArFbRbaK1E
DVZuOGSQ7uf+zqOfB14yIUKFKRlEwbv4HPIY6o/R4mxpkOnyg5prsc/ylCaI6D08
IgorGbQA7q+7G3n9242R7eM/yWmPitYeSZ6ZqVCpr6nWjfcB+OMsVic07Xhiw+Xd
4tQO+6Yq+3J2jCU77UZeSTcD4eL75BFaPtWFvoFXmGcCtgkzwpv/5TyaAygZ1Biv
O0r4L7HZhjxf1NuZRdV0fBZTmBFBLngf2nNkP8zcIT3TZ93qYxRgmOQDfxK7/M7X
9PBGFAv/alrr1g2SeSrQVStIc/qxccaF4Vn8E7ZvrhkTAkqaZi0jh0SaImyPwDcI
AOcD7aoReeGVb5gTmTjRdSyDmfxu5X8P08EgDDcarjqujtVyxRA0qFmtCY4zboHe
ZCOYWG8A4h/KDd0BAEB20GchHdq05inotUbDeDPcykPUZzmyT6gox3lx0JP82Zle
cyCoYUp2zJ1WXrzTQdmsbzRcmID9vDCmkMm7WLbawgD0wJfuQbbIPukzcpkHtpcH
qH0FwLOOdsNxEpHJSB+5XWkH3UKBQ7KkrsRkMjVopoVDMwYD6gS4UwL6xS8GONy8
RhQ3w9JAPM/QLVuAbgfPraEa1sPu9ficlAF1hh12rDMtoTaovR5IQxgRSm5nCNLg
MzRhqmLxzaCPR/St89E5o/PhCiUC38OcY/8Vll/HoWvPL9QUKayBcXaVctDFyIf3
ARhn0Xos7mjM0ItDWL5iH8sooGKvZF+lr8pispwBVR+w3mqU7WNaCHQcCkNt08MY
3JgWCzgkRi8W9BhkaonKPSz+swnlQCBs+whuP5DMsmkKEDR4ACruwe4UV6+OOPFO
O33lVeEl7b1CZSMaqOyWh7w7UFtPGvT4w6bXtztMD57rZUFkD07XUuJPnw0rXu5d
4DWJ8MMrm3OBTvQROF9xdZhgEPBdzrLfT2vpmg0Mrm1Fm9FM6xjMwJ3M1fXiTl+h
e7WsJXwOKjczduyYClT9ZVqQQVhwajJdyVK9TWxPZc00j3KYWe5pxagCM2LWFpEL
UW5ltYgKiTUsGjESdUOBcIzX0pL/9QgU+k7C+3uZFKw9U6bMaZcDVIIsReWYTEW2
SXyJypK4mKnNjHSHR0MsErUME36CEqIpVhOUn/yMSpluv3tJg0BpK49RM7hR5pQm
hiu+wtKP/HFdnbcmiDkqbLw+MtFMuGpSmJQoUT74RIL7zh90laec1sin3d5oCKB3
eHelcogJ/445blRhto2G/FadfekJ8RgOar/ovDWQikosNhnNpGIm9YShTODmKqAN
iq2wc4WSwdSHK64paF8wPUFHaTupKc/FKLauQTwUHsQWcjKOkntPGO538oQfu5W7
Fg1TY0r5x47Z8sEXJsF+GUAbqplEgJGwS6vgoG+dtxgCLXaY3CTUwBqDzDjVcnVk
LuOzLKYGKO/ntGnJFddQJx8r/XOSU+RNHkNO/VM9+ALnf+iovyGRusBXAQy0KqgH
xw6ChKRio9GYiYrjKIKUlPPWHryIdl0hmeuZQOEdC9DUkc5iH5T9pc6H+5lcCAfa
A3AJHDlvNIBNoHa40tUfL14sMiMV+xNC9HHuFXKMiWL1Zag9MW9wYeo/ryaw1Ygn
jB0IpTF+uKXlZFqWwYxGOKWx7Yux0zMnqt6VwWUVeI4qx75MzJrhrnD0LGyB6c7i
H6520qgv3pg7jzLpNwJl0N30H5a9aWolGZUSbdKzgZqnQTe4+rlKmVsH4HWkArUB
lK4clBfm6havcwA6XX8slpBJexpBT2iFRIMGc4w6xeaee9SjZix8hLnkkG6ZyC2H
nFqUAfruMsmPEr96YzOGe3QT/v/PS0g7SmQQLyvaZ6NKGGTpXwlUeXF6NmsqAwwy
nziWmn1jfBz2+/CDooUeoGN+qmr3yxGqdr7xvZE961kw0PQPULc5wF5J8qG5GzYE
88dW4opRR9LQ+39lGE6Tvqt8SuXHFTCxhk+Wpf0h0iREjW/GuwRJ0EBM00xcdFd2
ntlVxgdS5otDdc97gdOni/bWKFct3rXqbRjV3sAjLfJTtBIQ68u600FwYZIhFqHJ
Mm+TzLEZe2s1uOeQT4OCQWED6ARlUPE9t00OaKPXm6Bu07/pqNlVCxfjtOj+kfe2
VAsjMZ/XA9aJFjxFNZ9nD1qdywvdrlbyESlwi/SJw/ItY72vDgfEo6yRvsAiFBVV
JTzvc997v2Dxp1/wFthL/IBmq01ZNXVXb2eAcVEhANrqexcbQxaN9FQJ6sIcDv+S
pc0+wTurG1m/rYoib/6EhHk3Qxs0veAUXsh0JqdFQ1tEJLB4/876jNo2h3n4FD9x
8PHBZDhnodGM9UfMgc+qcruPWssyfaaAob98vzPr9AspUBcnyTa4Af0XIeIiN6eA
rOOCIfRI4oguqMxolmpMAQfGdwRUt0HMtAIlcCPiFQHFOQQRrBEah/s1juWxq0yl
h2SfpsbZt8WyFTCmU535gnzLbo/SLyzhKq2UhsPdFHpOJn5D9RUwWSc8vxOWLrkI
crxuLk3i8/rZf8cNexIwlqazR9KSYzYWdQUT2krUvlZF6fcQpFQ74+frs1XF7Yi6
DSSJM+UrkUKLgigXhCdkS7+Cnuz6BPOtGeKrTwxoM7cCJugxIHten9jbNccozG2Z
qGQxwlJPTxFRALg7Y610ore9nhZo7OKGuQDCzzMGHzRufZQBdFpk50Pk+3M9qASQ
n2hXgp4bvBoAxhshTuq6p/t+E8o1SX0u7p/tzcwRzcKzdmucRJWglvOUpMPRpE06
0j+mkJLgU+bqRwkr0BjXDQQWtw0g4bkv7oEJg4qVZzT9NKo0Jz3mdPjIDMcEFMVr
3gVEwU6pX2ze74kBo5VAgjUsPYjNz5jm/6lPktgQlUG1zfQ8CGnWtsB0FtKzjPTO
b2NIEgvN5plZH9THCmaz27HalgLLFVlfUFY7CzCqja9ynkJI5AJSSu4uzN2Uzn92
joolC/2BQHjae86fWO6l0dJjs4g9lKoBJFvIZGUMxUAMIxL3pgPt8yyzpbgDhrou
LD3k7+UHEXwDivfbhVoRKonIN2UMrCf52Emqdot12DOIWMhxpdsPka08qz8TMavN
oBbxMqbhEbErQJPeWW4Im88rz+LGQJBxh3zE6f0vX6/IrgJEe7tw29aAGhQMQ5wb
Xqpuwk5kU/rcDN9Xe0aRaIvC6E3Cojn8J+51wAHypYkkQ2rB9UbJe1LFFxMp36Z1
IKiI0UVvKpnRPPV+UPn1wlzFDo/WvvTNYSPi/iLL3LsR/Ct431mkxPYme/xVJN0P
evwcZM5BmrX6igAojDbt7BwbNsSHeL8xL8IAKeMviSz7lCXjNJZnEnCIh7bFxEHJ
xDKYnGDEz/Rx821D9Sgy+u5lReYlvjncUtZQHTXb3ozDN00m7rIsh2lEITP32OpM
8xb3gG61sMKPTNiTV3AsHvQVXVaZpWd66CCTtZ52q3lgZzFUS0SUFJqoaxBa6k5k
sRWJ3q8CwCw22leD5o5uABwC52MzeEUG4Sk4cLRuV7tg7gY/N+E7vukn7V11olzF
eoEKn2ltBhFoGKfP9iujRMK6GY3v+6fZfbvWyRiYwRncEe/+piW+Pf/4HMMO7+Z0
ST2V3YgjvnwKIIwgMu7ruYshm9l7UP0Q9+r0FewoA83rDMEVrDkgARyFBKhCh88/
EqNnnMAxITQ4/enrkYQ3N88d93QvoYdyIM2W+u6s/iiXc6yga6W2mPpnxUxZJo+S
h5Mu177kC7Fu4aKNaLV3gZQHsmQejXdhO+syuc5fo35BQ8P97wtlMixRI46/O1iz
/Nb8K3bBcBY4M8Sz74u8E+HtQA/HFfOhveHUELLVB1A/sjLvNsrtdlDbzuO5FPQ2
RZvZJKN53ojqwELgw+zPE7X6U+VJaDxcTPDY01amITx+a5cJdehjsYQ4kiMCDjL/
bMYBoCdd0DLzGp7JDEi7DVFdqaYxSw9buiwiuklYTkMBnGH3bnY9bPnZqITD1n7v
VwGWA+ABya6mM87Jqsxwi5I1qo90sCoh4ggs3DowVDCmj/5gbmujeJ7a29b3Ou3q
SRgW7azj7MDLFbE10cJoQ2VLNTTUGo176Yl9YYcW/C1OzutDDUT59zNktdRWGXHu
AxMCCJ7lxATyZLyCMG/gsnXLIIwmC20TLV5ZQggjWROU6oIJRzuS7SgV0I3nEH0U
2E1Y+Ih2rP+S60Nz/8N+yDHfesbv361f0pgvbkreV7d1nlYOnaGm4KyW7wU/pEVL
j3wz3qaoVPA4S1Wwt1hKHh7eGg666DhlI5CTqmiLal9BFqn3J/8p5ndXE9Fn4t06
IB1EbBzLt3nODc3xnisodeZEsStHKyDc9Gb6UBgkdMOlhqXPOzJq5NxIvBGrJ6MF
7+LFCV00XxExB3CehCfper2CrN/J0n5l56zTHBynM3nbBjAzIhZtsTZFCXhyp/m4
17bRcIni0+iw62Tld4YZlDijWApHhEczVzmCr+WVc/F+au/smN70eJtGJSC4OFWK
Qd4hEwqe4jyaMxncDlK343c74p6MKD46Vc20y+t63AKe7ucaUCXYkTrJnqfZ72h0
CI5CVK1eAuk6N637iQBtvKyx0Akbvl2U+JJY2znJqMjJroGe3Vhjv7tPJf1dDMDs
DvPz2WcgcT4njLWZBbP4RxJBhPTFsCG+VsAKAmYlGMe1GrCEwRnsSr51YZgywqBt
9o/6nEqedZCJJAqUbDS2G6l6+ATFVaRqdcwnog2SqtvKKtzLgwXjjo6b60bCTnCu
GCxqvSj7ST6U1EgYh1QDjNBCPwXFKrpNo/RlJprkBbaI1KSB95CXr5HJNzbEM0Az
MhbVSYexO8bcaC/JR8k11VcQt2PIAJL4WvLG+bXVLCX6Fxd2SrKWj0S8OunPvGbM
oalOYGxK5ryxTIjkizoJyxC66tpj6M5XM7lfF3URGVax1UwyPTkoSa/elR356ugV
1uv0WISyMySi8Lyathnbf2qYgFllWrILagZL+uS/x6KTZJFJsVkd8PAheWQZvs8N
MBGsqB5faD2lBQs0QhugLlZ+w+S9CfkbH8VFmOnMoKr4wPsQG7r4qwG4yRzp5NQf
dPTLbK2V++x8mQCd83eVmjEu6QNAdtZxK9ijKVwN81pKU/DAwF1d2k3VQdiVYF9G
nCXsrsuIqy0K3jbH1xHmYnLUeN64rEXlltxmr5HockntJaM5R6NR0lkdIniy/yVB
1Ai9EsMY78/f+Q5Ia9V+u3snqfWS9dsdk5Z2QlzQ4M/OragDbY7zBun3PrgeAEFV
FgsN6M9ddVgpPHDaNrJm1qzCYFbCK+EC9uEvHoGN3tQtbD89rbKq6aMoz2bMoeg7
I2HizYT6WdNAEkxHpJJp+ulHkV29crGXOC3NUdJ3yEDlPR2abNIx1p0YT4DMf+rd
JVGS2xW0Yqs4XOp8GY3k1xcbz+2uduv872per/c1lHUapj+B7LGvXX7LrW8h+WAa
iiCKfm3IrrQDi0V/UMQJBfEAu7M5LENcGUkQDD1NwMGYzGIm5mDbhOFhcdAHZ+mA
7d9xSdo0EBB65pbi+lrqXkThaPGPWghUTEBK0xrOjTDXFyvHZPZrdt8trLE6QgS6
Aw4tItDJqSyUMTKTq5bUvBl8dF1LanVMweN1ecuVzfVziRkL5q3azoqUzSjXLYzj
C+La/iRFNmbqOMsxxwFYLAD4ABXsbtjiBOZViosX7x1mYSWXLqlNMfFYJixdc+2f
3R9Q2bvZs8WKceRitHrY8kI56Siy8kCrgq4+jACmUe7ZKdDN0aBKVkOwpWUNDwdj
Yq3eBFCgLYvDP54JuqEHClek2X5us8wyK+zCWVuD+fWkPDpkPzCS3HPGbCJRKx4Y
Eluth6EW7nzFLMXYD3cjgjZV8Dgp4XQbnPRfYWg6IG7qs5XRjQAs07tCIpJj/0jN
vqbOSl1j184isYunU0suszL9Gd4MDfKqRYk0i0V5HJWu7tJAuL/4KmxcYoYbqKg7
1Fzi47Zvar7bcDkTZN8zk5/7kr5uJnioRPhEMEYEFL6yE+Y0gcFa/k41HvKbmVhd
c4W3jq4ZDWil9wMWtSnJVi+WEJuDfyVqIIC/nV6YizbhazaVqhSxLVDrhzGZuxDb
BrFq7FugW+gYDEOiYDwEk3h67fM1SPEen+x4pyPK427gyASZM5uDrG4TPBCj1XG6
0d25cDYX2Q4Swsy7GNps6JVE9v1yaZ17lyBi8cfcgfzzapkI99dAkHdPn7GOZJJx
+t9N1wV4BHshfIacqctrDMaZ0HHkl1sDt+OjdJ6F4fF5CVJbEyHep7JBYIqBbEQW
FC1gcCqsHhcStMXxVS/JnV8fDiobSXuiTlUWHJmZFIj19S5qMlV0I2jJwRw1VZiz
doDnKja98ng8krmoRar6duLLQW6S+RbWMBGgBcl7izsCvigJ4bWwemBynyVxPJI2
cRfhuGAKGulUnZAQI1RxNb6/aA6vAo9Q68/DXVJN3sSq9Mf4e02R/yEPgJX+4vX8
aq2TSpQq971O5+tt0I6qOqDYfQz4u9fNHe0kYhYUuokpuhonS9KnHa6GPFWXTcCs
sGj3/fxKaJorX8AC6ySEyMLTxyFDI4zHW0GfaTAkwdqB0GEUL/sRHJ5ZRmI4hURc
L4kSzamm87yyCTw3hkMiyIH+/5Kl+7h9etOq6Oa4BnGtjtxHi+Yszvw76I2iHYj2
+FMZgtR82qRS/eh+OaHeZvcVmbqfgTRHlXuErrvkRbfQpUEh1rWmyWY9VVunvJAE
w3mFfVe7q7Cqft2dREnWjCasunnM6Nzxp4djLDtjoz2z63YPaQHUBGNAsiIsagj7
43bvCk99B4sG4Twc0wto5Yk6/6xNt6V7fzfkU+U7yyiIouJ+fojNffdN3pguYw8i
qTgaDl2ol5j/3E8mnhMSKk/mP6ZxX2ROLZgtohEMuoNnWw3Q04CEmOr/QjlmjFic
po5dQfoznSgPCz92eiqHLem3nmJuzPFK/u3OlHzc4N/kz062UuRrI2ZQNO9p0Jye
nDoEif4H59Og5B5x7jMvrPMMK4G5Js9gCZCRq5V+PmMoTNawKvNYe290oAeEY2gK
Rc7x5u8yFtqOq4k9Hq7+i9Pi/XJOjWVMnm/euErsfG29XGiVNKEHf955vQd9ybQr
lFFrseIEU5Wu0UaTyhpvGKu6n02Y7/w//ks4QqmmFals5GwrS1obNH9ppc8Lptk8
jkqUU2uLP/9OgohlKbjUWw/a85yA+rFZYvNeWghT5vOvhj6XDB3ScRY0fEZaNeio
HTU1Zo1DMXNzAkGoKUPSEJ/rfERqe7iJDK56HK/ws1jd5hRONMMKAs6SNO1kQxnK
NzJ4paO8v0W5o3xjGAwrM4YlP8nkYL1Hvbf86cwBm6qJ5WaoANfD3ZEJWRnO8oga
XAfmhlKd4uqQLpSC+TUQm84OvrJUf6nB1bo+ZXbuwA0UqAnpvj8COuS9exKY+u9t
g9co05J/yDxoVWfDShqT4RKOaW1SaMHW4p7H5DWjSlDSX0uH2JMyJvUaCEmSmzAk
MVBDUIe0ByrIEZJz7U2LBDbJXwh3YanVBjHZHBZo38E1ywywzzZTo8S3cxHhIeYW
fcNwuO1pe09EsnbVOTU6nFEq28e0VXuLgY9hc/x9wH7LhLV4WHI6h/Cw4tghEpix
ilPplJQ+wL4UsJXsWHobc+yMGy6imOzIxOX7ncPgnLta9PH/A7plYBnII2hW4vbm
Je4EdIH1hQSYZHELw4t/ECeHZazosqgSTxvcZBsMWLWgAbRAkDpEI2izbZKvnkqB
hP8sBCIz4DkGgmhY15G3fFA8m75hXzxBsdw/CkMjVfH+/54aWi6iBMcqD4XnZYGK
7q7AEgo/RjoEZarPyuN31enWbNTNLe8US27Y2Ev9uI4kDxRtkN49rgXIpWbKPUd7
Iwd5fJG7pnQECfQ3wAWqXp9olIkGbmrg2hVKy8lzYTGQNLOaDy69MRqgSWwxFmog
eajmKQmScHPo9WDsTWXSq4/6OX9Ev/NuAHSeP7Bo86WhBcsA3agrtWRbqKRg2oSw
ik804Flbm/QcW+fm9VhQ/kmqImRnWLYMgT5YczPHSkklsJ+if9X1dq69Biv6nW7G
+uoysZ8lOL3WIVumItBMuw1leiDjGUpaYh93xsZK1LNMErdSxv75Nd5MoXOKUlfP
IGvfrnjD3HLYYbACkfPRnuy0MLP4bY9NipzU3t8FmbX94Wjz3etU2ku4PKj4C/NE
FJNNBpUuCUBuYviYqAaBLfEzPbeG1gEsHyal5iBzHMqKUTBVDzSbjpY9THe5inwF
gOAlyUHa0cnZxhXMhm9fc57sU7MlgNymIHiCuBBxvdCVA30CVxCltjhuWxfAGQSK
U37szL0Phx5fwOSlUhDr/cvm2/+dd0vRnLTyenytdy7UdzhunVdSEZu+OwTlM8oZ
am5YsWoph3/OwHUoFaIBiZsy7HxtLICjbz0Ja9KAV8Cb0kBTnMbieB8TqiBV6vHK
m3bwUdjvH2HaPBYCOO102tPDV1hVoTRjulJuxMLcFRVFHPyK0XSzZNgjOaDkW2Z5
UTusOeuudGZmdYfa4SzHmm2Fjnno0PL4pNIGjjuC62zlcw1M3Gzh4ZwMU6fyRgjp
QMeT0xj0Bhs1ykfmfjISHasGdeSyIv1SjgGR3CysBbyLA+cDeKjonGfeBeVxT4Ni
dlaX5tNKje0vV6pQRErN+bEkuJHdfoDnHyqeW8cjZXJa2YYvcUsrm9EF5AST6N18
yRT8Od4ZoSfYjm4H8InbvQk5bjwiyH8AAXYxeN/9FHh3E45oWcvCIzcWEMGTq2uR
MwllZqKnhNJxAInjSYONxExKUiTxHP0ujqxYFQScSbsJlFZ/9ldDFhX0eWFFXhvg
LS6rfKq8dDTYu8Le5WblUTm72WaYIlBGtJuAq+EpLRpUfHcNUOUSurcUILrZkeuo
HYAckJsOZ1EBlal5dBoOR5c18zQuFkF9clrrqfftVFdt1sJ7DupECe0IHOIJ118U
C5mHMUkyOLqf/OAL4o6rqiFna1UeS0kD2qDACjzbi/4eaDFiIMbpMit1DsA3LHbA
tcPlMNCvJ1tRbzIv7CObNWEjlmHho3Rmgv71hvNRsCjQtFY/wTFtjSpHtjz62ld8
swR+Gn55scKzHKPG5ygu0d/l+7RoM4q26v6PKRj5BwbOUfv9Gkghg/3Xe6Dk7uR8
UpL+X6Y77Y8bDUVLMZLr6attZdfhsEtV+b2u5FyaRAaFOXIadeCjCGvP9/WqIeCa
CpZ3SmhhRfCph+zLOJI7TC1yKdrCzaVC4di495Ytiw9mmZdhya8D/PbTpRu+IBn8
iH9AHsmCn+XymU/jgJieGJFIJGj6eJzDRkT89onr7FeQxJZCb3oDX1B8QbUIgnSc
vZ1T++oTbqBY68OzmDgvmIyR+JqPgn2PzYfx/uzBKcFjVALJE+G12pxNgQvWlLbE
CVLZB/GKYhxifKAAxezdxC312WolSeVegjUtxl+KYtCeFlukPEV36LVsVxRQSVEe
CXTd11CJfLHFXDm5LH+yVBkiDzLxEopXwQLJL82hPbii1WpFh3HFfRSCJpYbUakS
fIe/8Bfp+5PmTQlHoacKusR0jJLCISwoD5EJ5IftSbyOGROISvy1fvG9hzxuK2tN
x0T61+zJS5ZIFecbAXlf/U2eUXbhWVKW4m9Wyc3k9GW13IEdzSe8BsyaMFV/1sfl
agqk1SvKqd0zNL1CYA0ol94FQ4Yl4Ju/clF04a7RKoICu/yOp6cNnlJddFWXP1GM
uv1qnAJIb7NY6ideKXRoqkp3MJUkZSp4FIAyk5oKFY64qHN7hFFmcxjPEyXvPiZm
EQ3X2i8o/djk8vCbFGGEgOc2SFUBl92oDR3peom6WKcyamL1R7jkspz2OO3BlNCT
hUMepVJWDY6PVR7atcTQnMldBuAU/IyCVGnBkqRmEZ9/MuQo/QAyTquO8a+MPaBj
ndH+E6PAoLLpW2D70/sIj8U0EccYb2Hutm1kW6/Cask47g/KouFEgtjrnSJAKDZn
1HuJQaWT3YWwBqULAvtxKQDUy/+WRfEYrhP7enjjhQnfzht6jV6txIKrPP/s1XoF
COR8NeroR9H6oElrMPiuiUPTZjh7qWo/jZUPijDnVK1yGkKSbGJWvvhvCTArQqrq
2Hil0UGu50+yzWjrL3FZDviq7yntbpvrWlgPanh7nCMAX7YosyWO7t3DOK8t3Pmp
5IgiVD7QBVncGLl21+55eBZJsrcXvNfp/vy9N7JxIajN+3RZ1Px/apW7eChnWLce
WFI7LDYMNDINDwWIemZzuAOc6XcI1RcJE70YXln+FLXiW8wrjy16o6nwhs/dEJAn
4EKrRu0+edhHMDj76K09Zcm4VMHzpV2FXWWf8kVB32HJv1BVBAfyws8KHyDFNWAD
Gww5fhi7h+myjv/e0YVtEKDfoadAIRwdVG+TA101Md+LE06QDldAAjv4gVkuqV4n
x76RmMpur/Iy11moJVyc3LNC5n32pCA4GCSfODWBIjqtligU6NAxWAYvozI8zd4n
54qLwVhWZVx1eOigu7qcNWgWEca/XK24Hxxp8LpKbVqOpflYu6Ma1KdmL9bzzxH+
iGkStq0vDJwQPpWDzS41Y6HmQZ5Ewi5hWdzbTJZ03BX3GsJCEhK4r7d0HRZ3NRkJ
g1kQsNXKQCnyKATh39SeofSkt823+laS8KikaL169JsTkyrxXwowquq/s1KfA+vE
1aAh1thkw1d17gcGm6iSyw2TBroY6jPqkTtMVo4z4jpkX/PkkAvOhvQzOd9oF+Qy
KWLLi20U1lKQQ2vW1cc1PD7mddITPrq5F33PFWWg9G8zArM7a2GsoaNV2URS2vhw
++qvcwcS/q/gNNYAnNIExN3YKw9Z3NejrTOYKgfpt9UQxbhDtnyYLsvkjUrAhsHj
udU0KQfm5sct7SqugSYAExwv65KlwBSRtpX3Eck0DNL/fTHdPzQaZ161XD2ZNcLb
i9D4qQ8GRAi9QJnp2f1jx0M6P1tf1RlHL9e/saZMIDSelQXHDSbKR49/KxokMmmi
M5LWMJ8nabipLgTr3yFWo8AMrs7O8qFTibiv9tRbIrG3CP+mjkaPjcceS4AmIe/a
a9k03q4zmeXFu0eEy4+DKe4GC8D2UoOQ0NPE5DgU4hg20iZWhmfhd+AONbwqqn/9
xAxNWOj/Fq1vKpbGp4YrClwl5UsYITLhmopeKb2rkoLmK9qHqH7pKxMkKYXGzxcK
wJGPFZYoFGrAggJSJl2yr1ecvlBnTr5V598mqstnXn2D9ay6/TlKF393DgfvfCkU
bGJrF5pFgzoPMePDDlJpeyZ1sm/Hr69fpfI76RT8MMU7my+jkMntO/TvebpySq3Y
Lw9T4FoAEI5cUl3wxKuNQ1Ion+fNqq02RhDjo0RJvrNklIHzSGhW7nEVVuprsypV
KtyJfNqCSnb3+ZDrwIo9ysMai8kfS6J855ncbcwM6u1PIpddJalx5iOqnJR/spLu
dfGLX2laALePYxjYSD2JhXciFi5Ek4HNQWyDb+Pp9x7/X59yEh1sR/np8dJke0OJ
KmviYNZs+OngttLEgt7cOJdlCcqITURtSIGcbX4y6J/XBpU4aUvCMuNaQX1VDzIY
4KnaKdtbLGKRdcsG/TGaAHKdZpHYaRmDzEAwWkiYyiuS5KwpIPYjsb/NePjm8cJm
B9ZkeD8VALPMJ74/ygZuWCDKtJ8CYZDsV/y50B6FmV9367FzG1ckZP0R90Gc9B/x
K57TPlCwaQoPAoS4D/EUx+53S2jIzj9sW54Ug8jtsXvJ/1Gi1oQ2Etv/ZobrPwIX
2WQ38eu4xNzglHkH++8+5P7g1VUGw9LobWa1IMtYtugf2aCSwQtIujzykOD87wh1
t8yb+PQLLTDPk/AD782nJJQFaBcR+WrmibInNITeJm8/kVbv8WxDU/5bkI0e8jL+
GaZXPgSwLmDbF2/telvpad7RZilqgesMuH2elvxTXdTLt6/9cWHnWTzP8z9bPB65
G2Ga9dHn16vV5Vw48WgrcwzSNlTOvcdOoPlr7fHef6kZiUBI3rhILSsLXGwqn0Hr
pT331bQNz2jx8V5vptZSVBulX5qbryPUqS8A7i8QPBAlo3FIFHZrtX5J748hc6/S
ls71N5RjP29f656LaeankCQ3gQ4kuHZp61gwmf69L9Ljold4NcpGuhBNecfo1w3p
Q1DmNylmG5Mw7XFXl3Vi9thPjWCWsM6KA/MnXWRauO/oZNefhTWSs83zUNUL4pPl
R7h8fsQe5Ap6BIzzvV+krO4l8fy8VQAeMyunlOC9h+Qq+qB8R5BfwjVpsp6MJrlK
4t3AY3QsLSVgC0Ns0uw1+4A1lBG2h1XBItwVnaiZE/KOaoemLZPdD8NHJlWoIltL
XFLO8Akr3NoUe93Zye+7bpgieuI5q7plA8dO79QhQmBQPrJfEFntblaJ0XkRcBLj
4+FzihfKQ6Y8Ep1MDvtDRScdAa2POUY4kVFVWOZEg6vfg9hped8X3PAOI1AbGnbf
KzDTfPEImR2+Hbo7rBYEoUEsHFrnrJGNp/pBcsrg1CZpb8eqnNzjCRVC1vaEBt5n
SWna/iq7kdbTvhd58blQpLtp8TeCL2gCirG7WAv+FIvV45jh0/Ih7Vjrj4npF2wN
Kq43OqM8K2Yy0LCZhmnfLZ4+sEwo9z76AuEhfV6i+2Gk6Tlu43+GlfK5y1kvCKfw
Wrg6VZ3ndPWXEClgbDEL4smVAeMv2RA/MwqwmAlv9ofelL36e+mykbH/+DyBY0gM
juItUkWuUSrUCFjw+cpz1WsVSv+SdHGD8xg3ewUW/dc/sGKd0UWdmucHAXhjUUmF
O0pumBO4OypyIsrkZ7niaWfiqrUqX9M5jHiPeVyLF66huqXQS1670ZyCyIxjAgRM
b3LIstQUWLpycA7yFH3quIeGly/ArwDLDIXdiTRpyR986GVQNDyYgRDW7/T0vfcp
eW2nwQ0WItvL3DRVDqTJYZE9kAcImCgu38RKVM1Oejb9mZLE2pbKXPdHf3Yhpa0b
CpfQUoAQIE2iySGXVmTsoNxIYoQgd4YjjNxduFdpg4ibIfGK5ckfD6Pp6fjlt+5E
x8LGWZyl2NEZMmXas1GI1X1ODvGSkwSj2BxT6s7H3c7saRsbj5UjEvxc2EWl1WYe
7bm9fdktZv/kN/gfj9hyS47A74TVkNka5CUo1AybqVmClcuw0OgSI+zl1XsCLaDK
vO2Io8zAfnMvJglXVh8sYp0Ju8GrOxTJzP+K6VBvrqwxRegTI4K/jKyt6Wbxemvo
tv3OhPrNpeUMoCoCnWbhCHCRoYpHqyGHgygskDj1/doD8LWbUSA6oVJ6bVi1dcmn
nXQwMlpRHL5hCTT1aQITHrnR9Gt0mHgWeFp8Nx+Hi2LH+MlZxHbbB7zO7N5ooHKL
Wu8u8Fnc3hToodl1IjnkIUqS8Gpu3Q+G1ApyLbfBD+88JEyvXfdQFAGJFMp9x+b3
szOX5wVQfVKgjyFFQAXo7X/jZSGGNsKa1/JrCUkxZmTa5udwCRl3vIkuwQsXL/eU
Gm/aJn1mpexwyMagney0YAOIlsW8vZzyTIIGtsJrV1kyKweuqNoZMGzYeGqi5MhG
tOH27fDhAFRcNkvdj+0cWA5jiHSUoqbpHOw+yzdPFNpoh6tW6VefZuFcvqm60X95
3QJiVTxGy7yNxAdp94WA8+OnGpBEXxfThKN+z8o8vFXqR4WznlX4eAkneIUmYdIj
udjBJmX/jVhlpCMFGNSbafnSDNYuem185sa4DCLEr7zWOv6G66ng7/TK1wj+AbWf
q81PYGVypPVpXxwmJ6bGaLU+Pt/s4q0zVJRV45cYpTHdvwf/EdspiVho+RA1xa1G
ntdFqQE4TkTjxwxezPjrjD9z6N1gXDTdyn+PqZJeA9lPIA1cdrqHxnIyfyzjW0WI
NUKfFJe3hd0Rh47ZAdi9Y4tgN1veRitB+cjo3YnbJt4sA2hGjjqIn9b7FevYZyam
qbrFkjLlbpW8/N15GGwebcoQLcVbUTXwE9ys2un3II8ridtZu/LbDQLeEr/mB2O7
2MrKVf4M+5s1tmjj58059miZHE2j1UilEjI7abI3NssyZDK2IPtAPwmpomY8JxuF
6hjqvvSBDCOkPuZuMKmmZvQIP+yiz2nUa2V5Ygf9GfGLkXf+AnqvVgAqXCR+CDjO
RMf2kcqELVr4cvSdb2ewRMP60uk8abNjWyZlfIATEllPetXUt6D9ixtkZZGYvOeR
mjB4SJ8A/nCe55yK6hw7K0x6tJeVVf15PoFZYEiV66tGc/HSuY/WozdmJD/AhqQf
uc5HQL7EzluPC8f2zlplU2Y0AoTCrrnD45+Zgygn/QC8l5WoBVwmrFaXLpI2MOtm
g+9A7xjYNyKaeyXNzT5M5EB6XctatTJWgJUkIAGC/l9freZJb3zjBtll0xxAvxzE
jWgR8zsSaSky1rE97Ifg1ksSudArS73DBGrqlNk1Hqw8025OnoYwbT2M0KXDPA2V
c2mkIVNrM/bR/fRJfS1iM1yCjo9QyXFFxgXHBsUrOL7h/yPcon24bDygYKZG8r44
taCaLnwF6sKn3DLB8FwdK4GQD4fksagWJanOqkezNaGPU0KIVylOHCfer5Wk2qj9
t9iTNPcKpd4Edbh4YO/mlRv7Akf3+gLqjcgKKtA85H8RCtmd2SRyJOi8pXwrO59+
SDw2nPi2W9GSflt9Ek3VBPrDK3/egxmi9KqC/HUlPfgjMkN/gLbP0OXHP+Be0Jws
mP6X/nXBsb+ub1CjmMdrdwY47CVFLlWFsH/ygVDuoIyEMY+Qa6wD3iWOUXwE3CTW
vlKvVPoNlRapgNI9oBFAjS/q0FIVE1VmLpDDuH5VXTi7E/fre4+WC14B8IxjH/7d
FXJgyc93LwqKNzV8N2bII1n13M9EJwkXXZtpSjLqjFpTcyvUW1TPeKzRy1cEKcli
KKlM1jsNe4kebhGaRFSnwwpbDy0c9miXh/ErjFw9CB+hY5K0KkO0Gg6BYFHDIMNk
VLf8r29xkUCKI5lnQxRbvx91HjoscKZC64fI2A5Rjy2QSvYlwrzxEE5vOs5khyo0
gY/R/YIdUeAhjNKf+FYpGXSQRfWwxVZYvWYp2GxXTp+68cX+Hy0fBqjHDDRTos9i
tQaHMXT3CdLYS+ErpgDwfrr3x8C/lTlnZjeEWhiH5qz8kiZhH2JAjmkrnamoCKLN
uTzTMPw6QLqiy6sUIdOJe4Jngx3kOipfxLYmjhRgcbkIkhH4YmiXHFA38tJcxtXv
KwHMDGLT7HgtdL5OLLt7Ydjbapw8AQGRnR9evZIzWGbywAd4wY6H8tyzwO8VsZnd
NJdCWS3c+VsaXLN8IlurXOhSgNqfyKYu31Qu7wdFOndBW90YMh4XQOwdeS/hH47y
EmzUyUY5DaZZ3ngzR05L5o9+ig5zGYA6T1CSJpB21M8pkSbnKy+h6RvidJN+7Pqz
SUzmoiuBrKKCM9KMj9P1kxUPrgESCNS+56D6GUEJBu+mlGb48W4NKaUDagFweaiT
2Q1XSvvRE9+eydTYU8RNAbbk6SmT4UUPt/EptN+q2fypO41AuGR9xX0NJ5kEFyuA
00npgLK3luYUzQhxDYaZiwHTT4DT1MkWNvzEtHWIxh3nTxV8z2Hnol10jDbGnxAw
6I4zSftNo/z4UEVrkHf3nkCp8djnktoPImAmU9xrhoaZ+5Mgxe/SapQ9CLhnih6V
LhBdop4QD0CZoxC6xG8c3bYOT3TLviD8xHMPidFs7ssAv/J3QpA0mymY/T6M4YGv
vO9jOHlS4wvf8oc3Xb+cTYmxEuJ5D1w6OHi534kRpGfyJ+jR2oZNkk+0U8frtqXg
4RiGWPg2f8T+0BTmqrJr9pIlToEnDz0V1mfzw74BlDsho9BV9LoPmD5iMcNb9DMh
1++C+IYzPm3mrgLWjtkk2lB4SuyNSHk2QFel7OqMNC69jkqT6gRk31UjogHxl3k8
/ut0eQHVHEVRseGI2kDZV7iOgFsn2YJbpQ1zcwYXU7iyw+VCsGkgunehc2jtVaxJ
C+h2yol2TOSrZPSSk7uE7U6LOerFX1XA1L8/NC8AWmHuVUOdB7abFLgGXzPrZlJm
s92zwBFC5e8NjpJu7+MrFUvb1Gwl3rAoppOBdpzh1yq9cqMiapiDOKIUsLhqCXQR
E/n2LfWv3sj9m4HpEXA/W+gkrpU62yFSUNA9mplSsIBheaXDL474JVbYGQNDD5q7
6UlqBxYXNrbG9leZN3YthSh9n6StYTubSmAY/A8ydz/v+lNA3sF62xObDtwGs8SB
AO5S358INjTMI8OyYSGAUBiKR3ZteP2OSbzMgj62FkRDsm4BB2l0RPXiHE0oKeXL
obvmSqx5dDpVPdZP+WoU+A2W+ZuRTgkVBCb4HYGc3VoGm8uhzWoB5nSD+GSLON/c
PiiFLr0RFVvzN3vIlZAVwV/4615IsGEnR7zW1mgiLHfVh7CyUcrbKUfawhd2upcV
vof3LAwftl0OTLxugoXpDUHzAEyyx8v8jKrLHYTHDyZ0S2+uP9WuRrmyjvHHNq0d
46EASixXYxwrhqP8QPCBz8gkKDK3xDTDQvF/Jh2SAsuMoTuCT6H1b0eeNl9VR0Oi
L9mAjNylC11L14nC6a27nvNvu/5CFiFSPy7kOEsY6S+WuzwLnNsjF5YdnIkHp9iA
vA89l/Qzmm6uOZEelDnKVcSV1ymdvLCPTqJTYxicfMYZE7NKuYS/fh2EMH/I+6z2
qVC+d3qVASCp1v6ANt2ck6z0ykAVCuuivTsRd8Pxkjy+/RckoaxK0lG3LOb7Yb5z
h8r8931nrXoXBmOClVJ4N9FKhqZq5Vy6XEH5mEWfQNLyEUiHuCwhM0tUykprNhqF
4o9tJ93xxrlV1jGkJ6RQqaORbfRqy6G9ELywwWQBZVkohXanhNbSLfdePosWLiAK
86z6ESIv+GP9UFdHR9asL2fqFF0Ez3eKUB7EXcTFj6WQ8wn5kd0s7tvjtJoUK32d
Zi1knNyYTNY7niyqzu1eNWDK2wAbcir4hPx0C55TThI7b9vfqi3Uo3B8PLF2hPpr
NDoCBbr5jJbnhnFUPCqTjIji6vHw2FPc2KlsN7xNahunEN/roAxZBRi/WjzrWwVL
7ADQjmrvK0lqZhvt1nqdQlE5OM3tyvafMJijYz1v2LUBS5XBZZSe7Y9RMJHvtCnS
5KnZpCJ7TACdEGjHsjTpyTgSN143wBHrFTCZAXp9MEhNXZOoD+tGv0GKxBLXvB4l
HouaTMnESxA9nx2He9ScFwAovwg2+Tise1Br6d5sH3LOkksorH5THVji3zClJu20
dPLLuthZugH/KPofot8Tp/Ekv01RYm+cCXGVWg+vHihm9jHAPACfZmn991Mm2wcG
jWl/CTbjfORSt9fXnrkHnsRHAgL8DCxkQ4ojKu4Nmb1aRkMCeSTiaXvDMWE/lRZO
9YQP67mEJlpdE32XzHLbkDPFaDcVCVCGF+FLnZMqQaeJQkOce1Is/xles8IjU4tn
Ez7BJLdkiGBTHGZKDmMVeLGys3PRPtmSlR0Pd6RrFzcbbW2T7heDlBbQdMDEtl7F
2uTF4lPR7ja7+Y2bvKzmo/DrlN/DrvcTS9/xvJnv0E/r3V+0+RAKBP9XcKIfCDn6
PZTjrep34SSScXvDaxlepenM1pS9bzPex3TZ8o5tKjXyOPj5vaKv63f0IRMcEYe9
MfcQDo+cNXrSvJ9WSYTWipKIjbz/Qxmiz19wV4TYPFDNQnCUNgHNzFCoq4d3j0bV
r3ajBrziTNjxTuVZt+oQSytUXSw2id2upPetrcQtPpZXb0nYNzbS1Z+zuM3Pc0h1
C4fq2b+yiBB0VYdfTgiNqwjRmXa23hB5k/UYLiS9gtpij9mkrQCCNazV/MrDd+ed
Biq9CR+Jek9BgZshxpd1X9iNMi+SmGtAGnvuSyfXC8XzJ+V/IaYsOqRxAKzuHvGl
PnNbWsjuqn2vAdDh9HPOhaoGcRz4JNgxy8tzTMydsMmJusy8O94sTbzED+UeGLER
3LoLvAWhUPBvgRD7ZzubTgLaB9IWvg4Ktr4KYTyW1dLp+yYNV46ZnWhrpoizd1nb
/DUOIRO8Ml3OHFvOyvaFGBSLP9BG/d8wySKAZfZPpTDtcNBX+ABxO2Rgvi4n9uZS
tb8ofjFo3Q0K/psdEMEmDd4hUcumSIOuDJ7i+O6zycNVXI6HVDMnDdCaCB5yIq5Z
UjvwgQL4F+QMgm0XuADPQa54HJVnoV3JQCmbmSkmy1N+j8GpwNjtHnVjwKLpnud4
9CKf3CU1J8GD9TIfm0gwrRffSPJVzN+uSZXSp/I9esy4qkUGTP+W9NMd/BAq89qo
hq6H6us5zXwnSPawSOmouS62PJKT8QoWDR5Dxz8tmT5C987fvwatXealLH5/p+X+
ugkQUVbenm+ffeiTJH6u4iG4VDDsw6aIngyxFZjY357eRoU6JY6S4EpTQ29fGgjF
ziYL2LtJoOEzDj6bBOIwG5e5xZTq+xQ6dYjVwhZ2atgIeZ1HYeZeMdoCOM3O/yGd
dexvpn643IGfBsKbD0/HIbA/TF1ZL5Cl9ujbG0ZyUpz95MSv782xWWhJdtGzAEpu
hL7MTUzA7ODkfJiwqFI2vJw2rP0mSCzk9xgxVwWcmMQHtqvMBMLzchv+D6lh/I6d
WCKYjF1vg2yrMv6ScM+7G+PtZqILdjGdQeHI41IkmcQ1M3qSZXIq41Z78w8AD4dS
I3At0TMExu77/yYOea/eHm72FpfN/xNF+20DKl52rxVrVEArVBnV9jgns5oj0kyV
X5xxsFYgh682GeKG0BzH4U3KeOcDK0DacqmdQTGo8FeHaI8WwQPQaHOBEVLzsRO+
TZtq6dvjdIa0drAMj0WyyFHw6MUwQx87cbZ1G8+AITlFbuySXgR+1uHNJgnJo2dl
64Awogb6tZreQo0wS/64KSKLNFkfmzSH55PZOjzmDpQ2NNOaDQ9U2mT4lbLRLC3R
mvyFfprVKaslmfEXRIVSCVdTbawOM580/ZNuW9sdUaU+l/Fmc8oCv+JjWtFN1ekT
qCWlbUxl6xS3zwlzR1pHm+pwW3Ld8Fy88PoAtMNhVNw4dX154bKgwQfpFsTpn7Iu
VEB5tgeUi34o93SZt7J/iM0dLJcvdpvXyzMR8vIhwvGDLDkBGnum+v1u2mohtEbN
ScNvqAte8sO21cEPdBIoLyTRv6EEIEAtg1wx87SHdDmoBoqbT1DlVvwDBCzkEaFJ
1vAEvyWnXrd1afC+NoG2GvuHx8Xvnqc8ZvzmndJ+cpNPMixyQAD3uLneBgmK1P1o
6eKeG1oIA9luHWfyjuDo0gBTqVUqLBvmwMZAXVbmpZB66v1cr0SRx3Re7UBr7rDT
x3H0qVhLAr1nbri0dffCN0qlduLAHbFbtJHQcEGLhZSMpVfxHla6tNy4RtkhOsxE
xpm2NwbjuZ9824U+pxjQzyNhW1MGKcm7Fd6njWMDMbfKDyLbzHJJYYnc3AVyfObu
GZs4kpSh5/Hi34IphkZiOzN/om/xl8AMocA2YABo5YX7SR6UUluQSzpcml0MAmVI
kfz17Ah9h4Otmk8rD+fv6IIPVzesC/qNNy9AWjnxgEoyRUG0yMx+Ls70ZrHx5jDz
ZCXSkfdTRyYd64KR4ZUwzglmrGtKdVgvIOaKd27RbOPNiuFRSt50EFB/n1Z/IXEl
+0bjMeKmAfmJMejox1+z9tXt8cs23pc/QP0kjZnPTuB0n3h7OTPXhn5NDIF7ke+8
q4DAB+hT6wD7Xpqp5DLPVE7IuTm1gxfKSxvJ6/welnXsg31DhCIg+AIPm0JgFsJ1
jp9QWOq8Alc6Gr8F0JHyWBw719rEDc2IEZBASYcdv2IEOAbDlb2jCGB+B8oO9aaj
9ZTPiNwx2TNvq1wzdtKa93XdmwSaqNlJjP+cUYRrqpRUaiQFG60oLZPI7kJYGNMm
qseVQiQK+78sK9pcknnULKCbyBAvZWhkse1UGfTXrov/LsnpQUFUmUnRu8BZ21/5
MjXD/7zuMCzhXi3fY0HrUQxxZD9M7LMh96gLjWfE4p0SHW0UjXqiAfTlUvv3dltz
kzt0Hjig8S9GfFxggLZvf+rBnBmouXHYMryW0YK1SI0kz5a21ZGR9BUpdaB6QeeC
q5rBk79C0pXaDU1qGje/8aumA4dtmEKMAt5evfefl6gBswlAGgeSnSyjNKsfq/Sr
OqQESFAFIK0MyrUfzDpZHVS//RONVZak9D3FVhF56wmQh7xrbDMr5sPdE7Q8XC6C
BtSw430rAa2L77xHz8gjn5901U+obMFXrC0JPbJVjSQ0/fsbpOnhGMV6qyotSpsy
Zi8c9EuFMSS0jo7EnY5fM53quh7LnBMjGPEZ6XDs5/Yv21AYJgwPZu8k/zrEYUjG
WlUHQIVuIeWVVuHSByNvWq0c+PiChcC3PJvz/9G0dGroer7R2GZvy0J64Z5r5Vn9
PmB54eIwfMccYu5SplhfvpcfXNMD4FZkl4Fg0TIleRLGBw05rBm5ohxPrnjsbnta
PVFA1SuzBwG1DELVbIHhTG7P65fzTd5GaTQWCD09cD0FFXu7wuV+VH1NCQisPa0d
jiPs/atl2iK6tFvkJKCMh5m+G3lYuxTKpStCJrbFj2AsBEqWs5HLdoUOjASsV5nx
DmzGOnnUC3bXRnCnFIfQmO0uD9YJP9fLwurrjlQHOwKpNM3ahPW9q2wxJW/Ozwuo
xkwagIN37KOZRT3BVnC350VjJ7zoMlnhy4m3C1AVtkBpUmuWKChKfn8Nl/ABYBex
4ak+UWBKbMa9ctyZugbE/A6+Ibxn1luWTFYjc/+0P1aOwySBKwHUDwPD7TBy3T+G
qXm+vNfplzEvJ01j7UBRVZiMfO+m10VpXpOJIh/sGRvUGTRxGo27uP2zJV6m1871
lk2JQZyDAzfD8qs4Yu1+ugEVky1HQLXHsJL/q7jeVDaB0ZCPK1fRAu3ga4matWy4
iA9U4lrIRzneO8QjQn50RhH4r9LMnk52JENUSxARxp8PZuvVYHdGRq9nUFpK3LEw
7iDa0ighE+6uixt+ivyF65UZv9mKe+mYGQtK3TtiWQgZ6+iBlmV18HTCuw91CGgs
4bhWrvsq17mYSnroDXNmy1SjFnScHhn5PLFEamSe77wAO5k3Q9P8XDptJ3ejJs9l
CUaeBx77syV5JPyMCb5WsjonWW2TuPFj0xHBCZhZHLpXi089vxxhAbPXYkn5GCVr
zC4BbDVbWvRInNlIsgBkG94FuE2LpsARM9uTaWt0LsOHECMs3Q4vBDbSISoqAejN
crXTE5YM5B/tmHs8uR0kpup4TIO+oLqovoVz8UAQTqhk2gov+DQtcQGVKXODi1av
v5PTyiZ2641eFPOsjZ4COR3O2o2I7YbTpP1iHax0LVeZG/KUaRgu7ZGQmf5V1HYE
/QGhug3/xdoiOs4AI4CBnqK3VHRvIN/zzJdxeYrUx2USoZf9nUh7nJbNVtCUp3EN
LxhRGxXCFeo1rUG6VyacaEs6FEy2wnX+RR9gB8ovsffIGhGNTwGw+pEw0qCoBTjs
AhIOwHda262Q4nb3zEBB+tHBRYR2SRoVc7TQ8QCHwrS+bjCLrMrw+OM0U51rP999
s2Kz4dAnX9mg/2680ttCOUQn5ckmYKWp0kntEfgmyWKL5fgeO9dvpay74LsLIBWO
yZ8ZVYutc/qyxbwrlqugfefmlTXaE/e+FF/bQkc8cv6flS41IjtfHWOyoQIFtGVp
7rAxU+nd2y/KURAien9+c36FG4L/TB6DtcRX4rA/9WBa4BbRt6EoaaqQHtiRvMsr
hbltdIKfx2iQPfUwlGDZJ0XjWuAmUeI/j0ItJ/JLQOSzoJbGq8qiL4BfgTA9HL+4
7hCN2McmbbJD+ZT24cy1TDkatpKjwMrh/PAcyqswkxydnIQB8FAokzUzBzo8HLsy
xMry4KORMsULSL9TuzJVOrJObA9u2gCGO/ue2gK1c6XGDyows3KlzcwDVvgIFXM8
x5oEipDs692dvMW1PKStIHINDgJPd23TCiuNxvFsVQQtcANqywRHlBnjzFIeJcC6
ckFgdZBZ3Sorlp61XTcL/RIk/BAW++ILPI7lsnfQvpXN+9YycRW6Woaz4saV1xFY
KFV9VH6L0kDWmgJM04vDJTygZrzCTY2hIM/1W5PGkAVfpJVB4S7oaHU04qF6IGL6
DD4zRkW78DkQme686rCz2SLRmHMS/ML403X48GGqRQ1W3t2qtOqYaVPp0Z8loWFh
R8bcR1+VeLXEB/u7HZEKohAg/pWJmM7Vho/pypw9yiQ1G4aqlxYLwqrRMns9qVC7
bCyrj5wkM5MKEyNWZIhSH5VKIoy6LvxPZF19L4m55ONYKtt5QEOEPp9v+0RcAyah
VzOCi19NGqtBztcMYgVNMbM42+Ton2xGxz+76k6PYvElGmVh8IbkepjDvaay3yEK
wjjCFXK+gAGoqd9chW4BwVLjsGjppc07yyVIQ7a+Tz0WA0ncK8JBf/vP92SuQU+s
PfmDfxVccvDF7K4SvbvwO05T+K2dvxWoqR39f0Z6n0g+joo2mpHhC4lyw2ygz53A
p4bDMsf4rpFn63mrnCYwv4ypsdh6KgirRZwY2drnQxCYCAywORwmvioDP7Lo/LDq
+E41N+JnP/cOUE3VII6tu2TkcbHIXqUFknXvMK5WytyCMWzXeJKFbPeBe7IEmw+x
JJNZ82erreN+aRhqit2KVv4guVN90DfKK23tP/ILAgX78JmX+C7lj7oxQoZukHfC
BxM+bnSpaFJhuViAy3wnSRHCB4mzbjy99Aa3oIoZn2TfUYgykSdv39I33LHn6Ez6
G6C3i3/UuccOy1UPi/wFFaAS3uBMB5M4HvClJvaKXxeO9Gbmobc3+uuuh1SCUxgx
87t+1Qf+ETbRX7aDaGA12BLUYiGhoSY6w8PaldXK6807Sd2bEzHTs6AUII4Kr0R5
KKryzu7fTTRRhTAYUd8fgVRYFk327HxXOdZdHGItk0GGXHPgGNzYn9teCB7+3L8Z
OZ+MdH7Ee+QvoxXnPQpjvezIC8NC2s7de74lA5rxH4v8XXUAtcREld431/sayN0Q
/h3HEa2b5nOHCNlRspL5q+YlVwEh/okvwFiTKaI9UslwI8pI7dlNdLmbYLB7A6Oe
+xdFllB4y/ffcdatlTDOEitlZ+ywGuTwXP/aHJ1OgNzwlpYQ0jDHSiR7bqlA4GM0
5VIGmqLn8ZQqSTMqXq17vlDB8Dl59LJNgpM6AsfAIazYwvR0RheJMqOLgWV9FQus
xvMxZ5WNCXz5sJ5GUKDJBfRcjdbyGe3BS/IGoy0X38hW73VhodOM73MagaqXamk0
FYMoqOSHUH1NFoufQPC1umyqlh0J/4XqW9fOjvO+saZwhdBFwGX5LnsfDgAop28Q
NNN9meEGzXjjTBMqFFJXPn5Y2JINlcBzrom5PaVNFDzWnvFQKF4l8VSMFcDyVMD9
gAWimCYGEcd7KCkD/gDbd9onN3gEiXqxxyeK6mBsFxZtJDnh5+bqnb7yk5VJtORB
aWmRgSsafJa0uRVZBLATPrFeYfpi0XiG3V0Mwj8TZUZW+AA47f/fnvf9NaySapsK
qFTDEDLdaVYoaf/+arrsyyruxvlboRKo4ptMk9pZGIO1gtvtcB5UZ2R9igHfrEwy
dGqtmHF7HP9b0O69dS/hE6BOaFrmX0TF2Bi0YQ7LOZD9fTTB9pPv5I3TRAPTkJ7N
EO84nQZ+sOCf6aVYjG7aIybQudWrQc95+bpMnbeKINqKsK2HRQl5rUzaDqHY6ndO
QDlBc7gSk62lgW7d3uUZH+Vtof9B7UT/qUszWfKCfm/Lvhp2OMziRozVyaZbIBOk
/7HW29q4fzJL2/AC7NuVjTzbAT9jAwz7VHmUW7xE/1ZUn9JGHNBvlzFqj7KKqA9H
YDStZlsuSrLYPO43HbvUQqZetIyEWO2YHznKzhnStspQxzNR3tAisN7iEmzygjJZ
VLCADZSYezxQa37bt4w8uBf9FqgIlryqZxoO+bJO0DiitxFhEHeNrkJ9rphgzk+G
qVs2tNd68NjsOoCoTjtMXdfIb9/EQjQ+WCWXEh1c4xujNjtkHPXlyAZjvYh9rFRB
++ur7ftaIz8eBrbKpCcJJTpqgHy9W8nt7x85jCWfBlcg/N4ltwPEvqLZfeCinhSV
c13/6FK6c6tYrS+Vpk3vh/iph27PZNeWKispjBf6und5hX/CphYgEdYpRsN+e7ml
ditsTz1XZ7bflB9pQhAD6+Q8/An3uaxrS8HCV0H4a4tJAYmVcncLV0lIh3dsbVFw
dHt8wXocKOA4Xmfq9gKxSYkfaZ1lHOE97H/dcdjg8B6UY33rlbYcVvX7GQzEMcJN
tIUXoWqDvg/dsVkYadvdRaWE7r5knzSiXYFiysXHGC99IzBGGe3rInOYTTZZPli8
lQKjtlJeqIbCpi9EHoH+ZsuciW7CGkZ40842VRQUMc6BJi7sNmsfx483IwuETjKd
U5Gp9hJIwbAISEDvzoFV6MzOt8ks7fkCsAOJzAtzDoKj29cT/FVvOPtsv+5Z7Dwt
uNzkuRNyddfKkrKsQD8abT8uSv/VbiIwKM9IXUb1gwVAxd7nO8gzR7lVDpcHBOSb
xaNC6GxCYzL0hUkcbmj3MrsieCsD1RS+Nf0QCS9DZR9S9+uGPqFtBqCt+b43EE6w
MPmE3DCOwGW+HHfoS4tSuNbsnivLXlVHB/broT4W6O3lxqdix+/W1fCpvFRZs9sP
vDg7pJR8qDy1uBJMmT84yl5zGWz9+mCUE9r52bzrQtvJFovfhygiQMtB+q6Vthfk
YS4/2Wv/dWMXkFQnfvjMjRsI350tSJFSmfEnNzth90OdApEl3L2/8pPLmHv/rKtJ
ZXF9eUu0CysvEvs2CcbOD9t+EgqrVEjBas/LF6rFtaYuV3MSryGVWwUh6JYr8mCz
2YQ/J7GHlOdUr+NAHlfI7JtmDDoiJ/jcPvp4X5fQm0FHIDjtPv2aZwnehX1BY1IC
0JFwuXUhDcjv8Tb0O7G2s4nAMpjMDqWafcgbFqRrzVCAaFdzFDSSy4T+W8oJXCR3
7UwV6HkQdPl9pxJnAu63Q4bP9RS8yR0Hgn4DXSLwUqlFZ9YenMPp2SqJZoIba+AD
uYq29pz5NKxoKcAWc00GfDJuD1ZjEtxW8Nf6CbPTC7a6f5zDXUbP0uPg7D5zJfvG
xsXUiJ7jESqHE/rETKWbv7X62UUiIFA1UMhEGA0wNBtkkDZW2q3gTcNvflK2Brjf
nWmexyYrtHR3bm5BHMFuX0Rmtmiw6DSFNNHw6WwvHggrxZiKa2zspY8a6+IX3B8P
9MyBje6QLfXxEVSTLrMmbuqzWwV9J0NNfh612MUUFkfagaIC0lDr5VRnB7gPIMyf
Xd46wJ5gioEom3QwMoTmCCG2kD24kOvHP60tgz6UpP7pqo/5DhMh0FQ0LZjJdoD1
fl46xdYEJoCFb2DQ04htMA+WCjDqI1GmTDdZxCWssl8QxvPwHBQgC5ZXbW60UyO7
GdU6xCuTTlt3HJGVCj8u9PKIFbf/LPM5IGUPP7dUBuPdd+DHqSTaUBrlrUn6V0UF
SU+1GB0ByoYx9LE0QZ7aUjk3lc0UkqyBuSEgmPwrUSXCpUgb8cjWxoELTz6R+uwB
aDlC+mE6xv2vBmVRCpAmhKjoCGjg6h2k2PgeB560YQYWHtC4418v+GwvNsLPDiKO
xWKybDgh6iaqwFxt6Wykukwj0U6yLnQeJwtZeNRphRic7pmED3B5d3wyuBhE1+GR
u6MOqwAGv2NJsn7MuKuQHWnJ8/HLva0KWHLWrYhRPmweqTVZth56IBdAbxD2+LbD
W8TGEriH65aavmUejb/psVEbdKxzqNd+TFcdPmiJmZeLJs/tLeapI40u1HfRzv1x
8MuMx3S1WSlKxHw8k2BkQUztS+ENoSkyCa5Bog7KfhLYX476XuBJel7/al1wUJgj
R0j/RPyWz+KsJOJvOhMHhULpoh8HW+lLkRWQyfzQKK3bqGDSKqXpBQKb6iPwWRMJ
3N1YXZESuox6QTo7Daf9yo84nLNgh84p994nS83AMdjhFl7ijUx0q1WvrEXgArcY
ELlPKYPOl70/vjPnvY19usmvaF12hYvSHupRJ/nuNs2rSjNy8ls2fFk3Yxq+2xir
piF0QiA3bXoLPYI+VPhD/Jrro+egxiAVLgrymgGd5tSYXs/81BxTkQhqPN+yhAec
mScGQJHcjHtvjKLGDjSiglYNxEBLjQJ3pGXTcX4O3kxoUN6HRyW+kAPm4iuEAXNZ
0BIRA+lzcqBLBzw86L5lN2+XQQOtCs8nQIOy5cH0etRY3ig0ZPC5MfA1rPf5QUi4
VRA9qZFE6S1Jsvu/RdGJX9AiOuVKgx7d2tZPlYFATFTQhZRzQL8dMQVVcOZryGJD
w8VLdgWtoIC8dl/GvA3IwzUPEpfURxFmaMCuC9jECNgR059p2O7UL1TSGjcADzM/
jmQ/NTPV8WCyER5CiRccGsk1WEkcBc992Nz5PdASqVqWnebbQhDSTxTo+FzQjaQp
tocwxw4hrs7yFgJUdVB3rSgAbwGLw+9Kybz5rqUlsvaX5mOHmpDLLkppZJ5T3P83
rt0zmh/2WURQ67JgkcSYaOA1oe+MkbBCjxOumMT+CvNHOKXu20yEeg31IRvFfJFd
wSFnooqKDdgfVpiiICVd2JuiDC489B2WndoX7hNt2KbUDEiFj5h5CgDLZ0Ik0Ej0
/WvfXTZ19z/rE5r5UIFY6+j0g+uP9dWX1b/RtByd7HWh1AkA229liIHW/SqUzkfP
SJU2c9MaoXMZRI4keNX+dbGIXcJnshg9Aq/7n7KgIm3JW2bFbjUpzCztgLai0STr
LQ21P+5UqWFovdvSUyjPnA2tfEB3f4/6prmDTfdVxV67vuhZC/RAVAmv862ylEEm
moLo6B4TmxZziIGCDIjYZY8PD7adkd83pA6s/WQq4LKUmMpjhq9KieBRk1uMLqm2
w0U41y2+r6o6/pEEcMGKPOJCgowbPyrkELS6EY+1xTPmeoRmTpFWc3GQe2goCB3s
KDA7uh9pVU9q/+L/BcJaEPRp8h0MGQ8dtYncAwsLGzNxM9THZZhZgMC194Je95Y1
/Q8CujQ4QOIfuntYc20au2c0g9HVSzXy/21u8qAMUkf/4myhNwnljmR9M2EMyH+p
L9DDZBhO4Z0zLEljoxS22MsU/OUq+zYjTfOZkR7ioIKfSs4lXGag3J4tElk1EnFx
LibfCwrkRB80ErJikuONoHNtQGzgBqq5+Xe+dCICFGyBKkNjmq58BTOHXCVUdNhb
96mylBF5dA9wEqBKJ8UJqEu2YCscqSoJTQqdkuzsQZBcPOR2EyUNKFtEpOI7eo8f
lqQrAGpv3PMKDCqXmUN/FgH/cTIN7HFgmscTcglZGgj1UxKiqXbJRhJCP4TVKNkh
tSTJLp5gwZ/Qg2taBsLKk8t4ly4Jux4R39pzgfnpPy5FdYUukWsZUJoxn0jw5hHa
bofZCWZwIQueZ8wOgGYmSuBkRtu7y17L3sbY/yuqmkkc2ZW5Iz3P4A+HJp0tijFD
0Yo/t6sU0tIudsbVFnJ9Q5/TjTyqUaLvJ5SgR6GgcxHa/mnPuQHfp1iK3iUwEjBu
IQL8/XAp4e7m7Z6H1puEp8VvyKnt9NFvQbCFSWtYp5Hn4FynHzKKHbCyvGqTP+Ip
ltzTUkHrU0k+/bMPkrafpLCgzf4Se88cdI91g5Zp3sh9YyMxBhDBANY0V/dx1CmG
RlsXZ5Bjo45yAKQTwj02d6zL2BtCBPW5eekpNNhHWTncNZO47qyD5xaIMJ2TZRgl
3pAyWti1Q+XSUUfYTdIuZXKIt/KB3M8ejtTcXvV5p/MvKw5oWSyYCrIYknh/xbyZ
2EZOu8CdDlsRHRHZkv1iC+Dy753BeDwJM3jfsytfro+m+ShYOEt0pBDcyM+RLfMw
0zBdQB1wqlqsCaxAA8UXKB84QMKbTV1AtrI13bHtXXtipCwuwd4vW+5VRjA24ue2
lUlm4279oA2gWVcPX5Q1J2qATMbNUk/kPMr+rA4bxLIDtMmxTNg3yR0tEevPz5x3
k6v4KEhMFC1egjAX8ujvFY+uiYIZfhlQdZ8LkKT8NdK4aeo5dnqxYdFhHQquzqzd
UsN+37MYmfWIfjf0d+ZlaoA7BzzKXIDXqNlyTxGKP0bRNS9ntxku2/Et8D8Ki7OE
ZaRgmXuKzVEOBEeyl1UAUMOrgi1eig72cp+pqfaKh5YKiTI1YSCCx2tjMKesqW/Y
DM/duIBIOpXgHJtAvExhVUiCaEWcYR1JyfmRzEd4mtxTK8yJDI/8ewPjapfYQm+s
9hNEJTwyrxjQ3tbbRwkBAA+LlItTrDlwcnwymBQrpMvNezXCAgIe+BlMHcP+L07H
qVzduO3WTmMOol6ewrqqrM3n9E4iadTpzCvkPbAt3YOn5Fa/+ezv9g4GOKXjAent
N4ZUFKsr4NbuwXaxsCgqpxSftaoyfi8m6DK11qCMhGvb+MLtsVEXrSaGysezTOgG
DEFbSFnSJUSVBvLCAgSNkDnBluT77I+HgV2VrN4+39MMbHUvEjlhbwJiT81wG/ki
FCR87O2z4KeUhfGKWuJRBtjm8bVx5JwSyILQHexRlhVuu5oVA7I3kssaZxCy7xY8
wQfYfICbrTELSn4M8KusjEXrbjzltz+ioV2Sb1n3Ad/bLCKAjwvNUpoLWIeRkyRJ
PtSML66Qrzx0V8b4WCdz7o86ljMoeywA+MqUsUVaY/jih2EizaLDQMKrnWwq4EgS
Ox2ZV8+LU5w0irCKiJinus8dFSoKH+HDGaonNZsM0FfVSYW9nrqtX95lGAscKURE
pw+EXp7kyikz5kJZ1v3LR6y0nJq9M+kUbitPs1ZokxlSz6gB28RKXEC4FkPeipAF
CAEt15UBgsoOmwMeFroiFIqkPKPhBSt3LCKmKprRb6V29Q48Uw2Mz8/Y9NsB/eRc
Uz61V1unggFJNxhW8HeLsO181yPhrqkarS5e59R0RmTTWZ1z2+yxDTbhOXKoNtkx
dR/vPgJQG226/xl/vp/i1dfl0lABbPriI/vvxtPIzk+wduh67aDXZoBe+OM8taer
+ssjygk3eYk6UmsRWHfnllu87t6BfxwUoSYemJ6rlf/IdtHhsmzhtrhklrUzCBWD
IiD/j57GVRjFgosR9QGEjToEimeKDGUOHbeSNGewtydy7Sr9zNz1aKsGjmvND/6i
zmYZCvQoOLRC/Ysl5HCr9dtHpPEnMZZ3OzlO/+naYexyp96rScj5dOMonN0YfUsV
JAsOFcv7a+gVnTTbSRRJELRXnjl35HyloivoKRpU7YxQ6QYpCRRqG72jW9VIXY3C
6dl0aygVlrq7w7RXhBB2R4Iu8Zy63xuIxVN9gEeznQUBgIb4zbb4zn+BGqm8YNJN
ZNFWgjNd/8ueT/+xF1jMKXT8e74Ot1ndkDCBpD0AqkRSPiNSQ/OIJtcDHMHBt6sl
AuOlUfgJOIimVVM0IWeK6bkg2qbviVUvKavaj4Gxuyjqio78dUxql2KLxu/XqQQM
ttMGkhjFyqh8sUzxZWAiqEBaBxIbUf7EY5cYhl+2qRvxYkvl3aP2K0BgoGFHfKc5
OaXuPWxe9CuGdyn8cRS+4Hfs7FF5z43VLGfuJic0XNPLMjzjvQadF3os/U2p9cBM
SaeXGMa9IARslOCIQBBQ8LcsxQc8Z45OgOHH1KOfUtybecbDaDKEhWChGHGFv2uc
Njk1CVUQhBH8F57D5q3WPsLj/IyGn/cukaceEGBB6qAS8h480r9iDhjAGnC5Xbgg
kKcEmZBUdSauBxqvPeEgn8P4IE7bHASAhT4gpaVVyoISeOCckL8RrdSiwvgFOVBH
6O2RgOmaXJ5eWse7xhFMOSOEkP42Oi4AywTjYO2dGyNuS16t46zbkzlaCd9f5ZDe
DOZgtdHmDsU9IjQ7Pb+ki23Y7NvNhJQ9EXB9M9b7uHWwe5I5qKVjUyLKvJtYjXJl
XT6EmXXApBQB5y6Hl4vnRFNpKS/tpxd9ynZyNZvl3QZZtyAwtu0ufeEqig/EZ6Vu
OK0Wp5Q1Ftyr350FU0cI5McXlFyM4nN6DmHgOBgnh9yxfDD4cOUVeTI4egggxAqv
z6Y+2hPydpgtHROFWNzCM9qRsWxktAi9mLuTYp3PtFNJc99cXRfezheFtFoKO6Vm
ymFnz80SJaOLhH7crWGspciE48XsciSgoQXjCPiPOygZGN30fxTrc00X/bVD2JmV
TDcxQ2gi0TbnpnbVTLl9VUkoPcPfJQWnTAShEkbpucdQbuG5iTXLf9NxaUOxpcb6
WmGanrR8vIwztkyUktq4Cazf3Yovnf5lH3XObz5xuH1wxQyV71x9WhGXQXlZvmTU
tRlWcLVlUPeUwiudmBx+IYWjHC0XaUXj5VVDwApcm0RgIHTETtjiCq/PPro5n6qK
x9Q56NbUS7+C0OYpyuRjH8Fjyc5SpjzQzYybI9Fyy19YZgIGpyA7Fmpadoo8V9lX
5xdyS3BYTO1ZcMAer6l8RVkAl+81k9a0x4UZn8uWac8lmWhSj6mwV1oyXZJ1INgo
LLLoQc8vZPGnuS1XEiW0iHgh0HAW0H0vKr9iwVmWkPJkcGRmKrCMZ/74XFrLzwnK
w0oCCMoNR0AELmNBm5YaeuVsaOBWVEAHbmDmAzN5blQDWYL9HN39WoYOWUG/+A0a
inZYiT+vRld0sa8lkmTDGCx2AMquhB+0EnAX6xDL8f06b66iwigLYU04jabPizj9
X3qXcoW7TZDZzSwhz2WOfydZFJOdY7tSw7juTlOvgWx4OG231nYZl6CwmNqdVf5Y
OEgmKcSBY7pzSCn1CD28nErFdOA8PXXNiitBjYerwjWXkSBfHWyNl1yxCCB06io2
W7svHwBodq02maGXp6gpoNosOqlF05MnCm15+VqSKKiuIEDwvnn4YgEAOwfaE17q
JCBOo39rZthQtjraIBOluKSo5+1nKobdlQ21snYSCrUh/CRsmQ6lHp5mASFiqqhk
8b8gHiLcq4flzdIT8CAZ9G0UqTqR0o3sSq4pmnJyVxczASxx9Md11GDKwy6Ar1TB
IngLGh/W1Da/4ckmBTRsakhqLkt3IdU4p44ytmWhXsjHdshJGu+9XXdSnnuv5HX8
IkMbdeTy/U2OD1Svu08jHjFH7oIk4IceEjCzYo5YqkeJA3OireYREPSdUS9RBMyy
M9EU+q351I/8fFdzbykYskiXOMc/xqyiw1Tg5IbE9CEAgiC+l9mgkirjVHNHizA0
nyFbWSGYXD77d8p3q7ZM1tarTnjWn0T0vmD0Vb13/Hmqo8ROJigMfDaVJCVCE+X7
WYhZfGKM9bjXZY4PgMw0B/M/NkUIjv4NNt4ebx4Xg5Om39G85gcdDWPdnReyC+z2
MWYTTEsmwh1fC2PsU2CdaFR+k4cw+4Pq3Fl3NwJZru6Wnc4q9khKDx5h6C0n1dq4
2k34xDIWFVF7jbGDv6y3TnmSxaoOqtASaBGKLKo2wknaDRdS7i5J4DRLFg+dmSYh
qc10wYNK7VvhnyjMaWdrKKKGFLbpc9rW5EtGadwS3hPc8R21mAeOr7BJ8zThY7p/
HTRCsgcqp97dCXkFbZOw3W+X/AdpO1P3y/sTV7D1WJ5KDFO61OJQGIrZL50HBDSP
vAoYAjruLGBR/gagYJ2JCdtu+ZU02wLAYchM79I0z3zBfnn77e7NJ81zg3jwlc1E
TSU/+6AAHyVvWKATA1DaQqBKNtwzTAwFnYmUDRARZjIufUv/k3g7qHotziPOn4Jj
iaPTjogOF7pXUS5wcahBKwYrU64iqCE08UshL6PeIjIWZKn55ieoW031Nh+vvRbH
yHx27jt8Jqkk3mTOPGf1ErAbVfEQ1p/EEfh41eJfE69Sam3Xt86OxWbxKG1jueZn
4usneyxlYCOLTvjNWOmEJjZOaLQ4t2knQDBZ/YobOMzWQCkQVN23H8GrVHvbaSkL
7720gPPFszZPjlVYidjUpDudbQXpnwOs+sCXyeyK4PCZ4o/OpggTJYB85jsmN4TK
tIS/9dWThav9Ws+YbJVH0JnGCV/HKndEaULPtQZiwvrLyt+ETltuLN6ASTmTpjB0
J/e6hmECbPoQcOXsMM7ITQTPf9kAWb0s++AsT8UTGmLZ+ni+lvu/ScMKAxHVOypf
lh36n6VylYFw9eknafm21VTNwMtxGBTNoUV1KSoR3xufkSuDuFsot7dk1cvJQ4o6
/qJg1YTYishPx/Tuw+JQEQGw1QEjGjNLivhFMlaNlStgpKcxYV9SgvgbFrOlxMN1
SN1eor32ZrQY4tHR/RM2vzFcn4QudmOjxmQ5n9r/j/Mf0+WbowVnYy7/py7NLzG6
m7amCjhZrZrEXVvrx1GP2BniYzgWer1mYew3qJgP4DYNA/l8GawvlPY442sjNzl4
YhF02x6XL2TtllF6mRqoJemgrBdYcGsL2xlYx0JEy2gYofbydeaFzXLXnibRxq6g
jEQ9orEA1FjW7vqTGjTHr7jAl1Y3e0GnAoXRfx5DvFS5FitQ4HMzduLuMTyVHkCd
/EfWS7IZiDUsk0ZIGtGYfVkIz6oAiTCnfWtOoWSbM+OjXKnwhAcRhNcmNMCxXQOf
AjCYVzIAkpAEyXi7n10d13517wI2v9GenvHIOqSsTf2+9mf50CdaoC7d/0cNG4SG
AgjmKSYxgPfK+Iri9dTpjrafCr7jA0+8USDEjHX5stQck1a8Us2E8xL39Rvxj565
W9Td3ZYEtQ5jiJARi1QdCkbMxERjIr2P5apri0JffSZyGuNLSeHIw5/djyIngJka
Segmn/Iue/AcY20n09Hpjmo/5/EhY2ah0vmnhWEYQSbfhFCAQD7HLH/B4r6UI5gR
2t5wWXeQQkGtO/ZF+z+FQ3mNlN9rUcWFT8hvVsRIvP0lOy0ddKeJwlccwWoIknIy
Qyc/+df1IjrWv5sHHsfYNoN1suIxACX3LpHeCZXUjWRo0xy6wKxd0mGDz5B/i0fm
6k+S+DPsX6BF4B1AQr2CCETo28BYUSsM9uWkrGKlPV5GRkWDaRDdDUMyGagJznQE
TvQGKJV9Do24Wtnuu2IgU/cVBbTYCEzOS99YVXO4PzhmDD66tCqQ370gy9sMl4cq
5L4t8dQwpB5f89HJkACAWaOuI/N+ERpqKIRFcI0R4NdgV5NeipvU240ou3QuiYCc
DfiOiaUdcy+BCqF0jPU52lp62f7pBQhMpCouk5xnwLGFSdtN5XMH4pXoMhOlrnrn
Dht6Y0yj8JqFeuEDs40qnQSlpmIqcVzBjewUI98/z+iOUnJPdemOjZ7r94PeHJum
CUa59jCYbkL1rvKKj89BvqzVzsdVywLvtNK2X6QqYxjtH+Q8bOrQz9pIOoC1OO27
eeF6HP+fUlBX+GA+vTRdF3qs2IE7DwLcesPqZVtLAlRBHZpOd9RMWvsHlC71qLDg
XLF1kTd+UZ3jLfW7UjrPqB9J9HgxIGpGHa0jT4NFglDls7AduEufYMklMvj+yKGE
OMyw5QPAPn1Fl78+Jp3AF823VEqMmUdqWiN5sJ82fjT+mSpwsZLl3vrJFkvRER9H
TwRtVaJsamxVQaq0ktAHuCYNIsBCp4873ziXNno7aMelKxHQiKO/rHKdLOv92hX/
lZdZtV1n3vEuwOGhANu/oeHK3FT0SWRU5uCTc/LdmghlGiyoLFfToP5WrzTnLOXE
0JMcg6gVLVeeQnwcY7wrGrWnEnH5i3raP7Rp/cEZPhl2KI3btPQ6vpxgchNqVuAj
KtWH30ieV/o0a29eeGTVf3RWHNr5Xt+YySDhO5EsYzu4grN8XMdS7/NI13et/IDc
qXVfkxN4Jg/kyJ3PoLlfDum1ZNvK067Mt2FqFgSpVNef/QNpyDRE3CiW94keAx4X
2RMKaBNHGJGmv0yDCQ6RrZzoTCANjsOu9CVvUKIq3PPa1pVveMX/iqnwlFCJakOq
SythXW97PpsWYqEDiIm3KAb3DVMmJfBqJe/7Okb2i608qkZwS5wXMMIG9PvISrmP
YDgL/i9T0ihcqu6M3cL6/Cu8G46iTjpFJsMjz9NsbZvkLEou6GgEsjhra8ZlxbFF
afe6oTK8xYu3un5KxuGzfHfRdsIXF53/Vb1bDrqDU9LfuaqFAn3h8jBtZ7h7kk/h
4MdZ73u0KkXw6kYihhJ6OYs3ZRKxBxl4bH+ayiWbyhnEMRN+nYpJNJ2kLy4VGu3s
tbgdzHhVLw6fhPYQdxYv3mxRmOa8BnevMisDbubEvrlzSZwr8ef44scjzsivQfsD
RUNnZl9ijDd6WUaOnUYvxPjHlAk+0pVCbp0KNKU5nwsGZyPKJj+s3CEVlf2+qNty
Xr9oEeOOSlIwOHwQP/QJ5KNQh/tCxIZjk2w/fWK9OTh/Gt7SoIpL3crdBm88cMWA
Jjl1j63uMG2mVLf9hqg2Y2lMGUDDB/quB+Ix9vHfCod7M6KFLwQSYBFAsfVCghMU
4rW820BdX1iI7dMIrpq+FlYtTje63Ss71sFX/hmipW1Qc4AP9QFRsK4RiVM02Dq3
Sa1iZEMRw5xBU8BzaANvy03cl5mZMQe/OdiYgu10eZoI14WFET8GftoYAEakBbLp
vaZY8g0r3RCdNeqxm+vUxbFpsNIKPJaelV97Ab2lHC2LsbX9xca+DO72z+ya0U5z
+0GGz0HEpViOIlDBW9Ha9DvmvDhVH/yYqS+xAmpJh6mrR0mSsDog/eGPbScrYKdM
huUIFXp9mdAG73NOi/mt9f6mJVMNC+99KFEsytuomaoLIMjNodmZY41Rdg2kXhLk
61bleook4U4424NWfXrzYc/09L1QUY6EssaHs7P3ztjmoNu9Bjqj4r5hXsLGYpBr
JDErm08OKM/RR1u782oo2SSa9j0Sq2DItFnO7LG6NrA6RWpntOr6wROXweHDCAnK
kIlxrMSMIFSNZCq596TsZ366ssseneV8fGp6NwBzZDjMe0ZQkVlBLlmFQ3bUhowh
XIqpIOh0SBCbPgY9e6K2njq+zmlaC/gYD7m+M7nbib+l7WryIehy/9w/HYIMJV+9
zW2iJQU0UWJ8uYAZv7j1PWbsKp4Qq1WifTthsZCnIQEDVVpZFlvK6Qekf/czNPUB
+heLaxSpnOtqE5ZT5XfqLcOxxgjRVV6BFd++g9twCCyMVJ893vGW+FPcSVL8vj2I
XoDjPvLrP3ZQ0/FUgZXUF/qiLo6jladEVt0kocSCLkI8nsunGa0bkQW3H/kt7ZwT
17aKOfv4b4po7m6IsIfOP00o8YNbrx2l6bDf4yZrsSwJk1GSYWc+nyrXy9nKoP5m
CAiWM6Xp83MPPe0kmPWXvaWwbjMohKunsOlCK6pfy2/K9zr7FhfNdQ6MoZHdpEU6
m6DvhHvaUqjp3f4mlevz4seIjvv9fBgLd8xoMBdQRn1PzMTSHd7vyFvWmrqvksU9
yJexNZWS/L5IlfJiG6G6Z014kUIT0aKXTKJ9nxU4wEjLXzpnXIwYEplFRjolww8P
EZpQU3KhwzX5LfT6HVUzXmd2Rj2/korlFwYIIVARRQEQr5QAReWykQF1APdzhqPt
KO8MAARBhskHX1Ciq7Gng7ZsP2mXm8CDfp2XlElcB7FW144yuUz9SiSwjAmT9WVk
LNfyf+4rIBrIJRI2eUoEWeXK55/yyH10N9FP8Zpvx8+yrIc8cFE4MXynQGzMuvSw
h7Eh+c9PIQzs+bNWTsgRDtIYFPqUaaZle1eWBG9INQRGF3M5KQw1N15kHn91ewxC
AdPGJxLopvW5nWZpqYpbxgdLavXLd4Yp/BYI2Mxs0ZAJnZBYj5NMFsRIQrWQAwn2
yBmOflYfJLQSfQKEwD3IN8nJu5aRLc/bty80lZjatyj64VhDBbYcMh03utKPfNE7
IcLl6bwE46/rdTFz/ekX+NVEfJiHVrKQn+9VawEJ3dsY2I74xRzVhe7c3Krq8xjG
Sl1KWuj5AlcWS4nADnxq72xWFwMbwUnBS1eQN6RZZ11ZJpymzwFHok3esOG5FSaI
5IyGHYAhsk43akU3txiaUTfjzu69aKq3W9ZpB5UahllTuckOnVfBw/70iUBjliyG
+/8nwPIOmwPwDxDC6XRWw6zTGTkAKGVOgRJ5i63kcTGjrInUqlAYrxwtEnAkpG6D
lehME6qNC+zf38tnt0+yONVYyUetYU840FjVb9zMapHX4IqRgA13KlDZztfOafSh
y7hPm+8WL0BVehdcbdZSYbQYA28wvdeLY4H3qf+TooOnhhWOf/YTu8hut7I6shc+
RrWGmAkSIW/Q4yKgyU2Co6ldXNnfDe3xsWFldKcAZFhEaYbmjHu3Xg9L+1MhpUOV
i1hTwecg3nkOngF4F5joUZWFbwZF5veQiCtwmIh5O/x3uQ1NoWj0Zc1qn1Ag34QI
y2yifR1Iyf3uG9G4EAws8mjVc+aCwMYsxZqJfI0h56Y+HWmR3w6SyOamy42tQ8/h
j92orDqUfqsus/YTOH1Bb3CMcus2ZIuCUptRh4UZijdODNoCsisbmDgh1mnMBgxS
lpc30qFfZoVDmd0UVgCz6jTIU6R6fVxCVhO2e7IlHAgkk+VOkQlAxRYQu6dGtaid
ZT0lypBP4mLvix9bytDBEOCwWRfloe7HtPhuCtCluKhRQz5RMdxuz6zmzKwwGJP6
RtS2nxrlYueftCdIVCS/PO7YJyEdMxjVt8aJIDzKfOsrDnKRJmMt14+/FvfGmelt
UhypRvPNxQjHu1PbclNb7wcukCMODjecFMwNLdNer5+e0056AgndOVNiZ1OCC3wE
CUTMbjCEnMBXAcF0LlfILLtmVH4xnqbi8KKcvHmgCpCL3B+yqeJ9vDG/Mzly9IJx
KaqXJPfJi0sTTR7wCdfmNX1+H8r8/WQnWIURdSUDOwcYFce/aYSR/N59G/eX7Uyh
1ynB6i8ZpFdFsJZw6dTb5H9QZ2tOmkNTsEub0vZvM1m366lO5laCYHlw4nOZH0TT
EYVd1iY0XdhsxdNS2/cS/iMpN7KcJcslaAmW1DVL8ft//TyB4ImfygwHCNRY0O7z
3wzePmiVi+GzKnTw7MwVJ8GJAdiZ5pJXV77dE8SiFNFPDOcKWeegd6rmv+lDe71v
WGt6Cu50m+rGR2QlW/6rHNTRbNvmRN2j5TkHM03GDfLTW/XqTCbThE8sbDQ1IoDX
662+O9LZdAwCUF81ZwkbPpuodf7TUcFB4Z7gy6MmqiAIHzS9hvplIwUhdZQt2jQ3
03h8HAeQ1s1/WgDFQbLOtYYNtqeI1bWv0MCvfvcLuHK4Xwd1Jp5gLnfVT/E/2Z5k
KQ3ogP73QUcFws82C2n0jA2wPGj58/gFcQ+w4cT33sT/xM3dBDM/bkA2F+1byKF1
IddvnvD3NgjQlAM5ef1wykDN30f/2Xg5NepIe7gAhJmKXCJEYbNi7olE8li5SZiO
tCXJESMLEThDx7pBQUmEM5mKk7lkbusJaHlnTXz0bYTGiSvM1CkL8dcCx1pW9oxw
P7plyPLAi/YiL1jb76aqbll0oDavUy8guYROeunpTktXS8sgCPXNax/USR9PPssE
CCGeScUb+3+pRfCKy0unyQWL6SRWcztpWpqXeRpTWV5toIvgr6Q6rnBRKFJ88Hni
qM6O+zECHzY3szuF2qdMQGzRWHr9G++rr62zmZz+CNIpRkFsCUAKK37m6tLinf37
TLKCcXxzxukBYtbANgO4ZmIf14l+w3IhS+Uj/GKZWW2gClZJACsI5d9Q2ifexNKI
U4a+/VHT4WPLl+/o9R3X3zpv9muCXGrkrUyvw9vtEGXhjcYjNPmakgaWeDDSk1Xl
3YQi/5GqIYBM+pn+9IN7L7ufaM9TNsj0m72htOYsiFBoGckYvwkFKcb+JxHQRdZg
9ZU8STNdrg+3ThMqOrWqEHouVFRDnFl8TG6TptBHShB5ntjhODqK5EyLIjlgdNzf
Mpazu6ihVP6gYzWxIJdhthlSi30OJRbzW9MOzwzc+G+EpovXDYoygU/dVp/N1G5u
gdh4pF38QVShe9zn+ZtFuhyng8syNyIsuJZ10gtty3pHid7+xJzb/xCUowislxCk
epeRqasd7wlp6G6gUixq3sGHEeG0xVbhlB82R/6moRaL6uFZWiZK4na878BFghSl
d+Q6tvL5hiO0xl26TOVsiDE7wSzeOF0PQ4R1ynCQ8Q4UCn5eQTJ3NmicGj4XgWI/
WfF48Vfk8DvzgY+yjTsZMiMHiC8MID4H5idfP4yP40xQHbgRFnoiAOhIeTN4XujH
+1f06wPPsNFRRlZopUqXAPn3MUQHzKN2SWcya+aMmtdfcJH6c/oss6E9Drj77PXu
ZMfUzLZE+AN5l/9p/fBn9ZC/RPdZmPu/w85aOaFyvGn60U735daNAUEddzPCOjri
fpqegFlR9K20I0/UKfyhUK9FArbmPslyF9Ni5h/dtEpbkB8XIWKR7VnA+Uqnxb2q
+9jEAQd0GEFgSV22y+wFsJh3AaskA923fUXdwbPB1SxWNZ7Q98I5suGTe1EtQi7J
cd///lApnbzDU6BJYWYmShWXyZY2bp6SfFbaoUDkXDnWKEN9y8WyDEffhP8AemZ0
en4MHz7M5jvcxZsGnz73QTFg6V32gKR7h/vBl4D/DJeyUSDB6adspRdiof6ddcxz
+3KAh9qFIcQqkoFWL2kIGqRFCukZfiM6//Q3mqYGHHBwH4K6bMfQoQhhNnwItLG2
TCq9Eup2pAMUkJHzc+lT26ms6HBNpr0uHKYKTOjqMKk5j3I5wwRjo0Ak/0+xfD6j
OTfrwD4uCWqocXxVUxCs5U7FwPT/nQ8OYHsM1KULA3whukqIEfPsMs0S80mWiAO/
eG5HWga+Y5zIzf1Kj68wWw4w19juBUzca3dBvp58pKZaziklVVF4K4oYeh4zWkB7
WLk07vJk3/GTsiq7qQQzB8sEvreXKpqMtTNeV/JV8GLlXxuEs6cyeHlgK/H1lCFg
BZ0u56eFX2GgUG2UIfKoVPmNHBJoMmutz955wldemGfSzHP+ZgFbWGAz559A/Xb/
lhLI3y2XMV2EyaBQtkc4jj/Lz84wjNQVCSbX6VC07UrH/7wZsRThLH4UbB3W2+Dd
hkeq3mDRd9ZqZUyk3A/0uNMaIQEIoH1ctJAIctB4aGRjA5vbaOSjPHYZR37c/Yi0
kZ4MKF88BvoquqWgX6MC/bSsp9Je1GSXT8MQG7BgYYoykNY7zP+s/74AkcUdPA8Z
ybvJ2arOnrMDC/qs1w98hN5zOr1Ra6fdOMP6IkliS64VPReOp7+QkpqjFZecWVWM
SJrKs3mRUrlypCAGcRViRaunyhHjTYkYeU87XOtyRFaEcROw9sT2YLiPzzc4lK68
ThV66nVAPJGfmj1aia4S0pE5UhrEOdf1QGVv/Orz7bmv2/uqsExfPFV8sy9nCnwX
efnChB3FQWuGEBEBZ626qhmlMDroKHBkQXq0ELqQFw4CPAOAfO7fwOldbTKB4DVi
mGkvwiWlZVU4TF6cRKLR6GtIiNxqfpj+n6GaQKiBwzjdvfQXDubwFAozZVvnsbPl
Z5lZ6KkG4/M1xs3jX9FG4fLjfbLm3A32Tj/I59SaBFyKphtHGGgBEb1AH2y3Kp4j
nAHOkczjHSy0G9p6EKxbfXUgctwmBhtNV2Ib+6Cr2PtU+tPQPP3b5IfNNF+TSATH
2ZnDPV75U2RGbkw4wR75tHdjaNUTBwl+ifn754BtA5LZJ/eXpzBBo2hEz3mO2++h
APUhP+FZOLx80JVSMz7k8EkLnI0XZ/2h8NsnbDRZ5QhcIf9Dr8ujswLKdtcC+pMK
gSgLYyG+nbRylLPuUyDzdFdZcBL5V/oVUENZZTen/9sBxxdhYZYamHvcyc96n8Fk
NuBTv9qt+WQ4KKK37K4hjSkt/lweTofyEhAnbNr1biLz4XBtoaNwvyjjIborevlR
1wsYuF4bwuHcF58LvHvi8vPhRwevLPCw6HMbiUaT3sEvqzL0HvDm10AEbvsYhSSH
QPT/fttWaxIK/tsxNLHIrWNMapkysDkI/zVl59IgHojeL4zsYWf6dY5UYDcMIQxN
PQd/CrZ8FtTs4BBSyQuiztoj5CTSQ1kV0UJvcK27+kOEsFMHUKh1ceF/hNHaSFzE
GOWE6oFpE8H4kJO/7UAG0nwKE+4wMF8QZ8qr/6W+10c1tywcwENWD1T+GZoxSjpj
SKqXblapZPl8ZxUyvW7cmPOKhkHno2cJmUELWI2j9BaUB+E7tabMpT1qey0YOhXZ
hYeYDJUGA5OBmA1U0rqV43MbxdGPwP364y2OhxcnGeJ/W2LTH+q9/7HlD4M8nv00
vdSEpdJO6DFBs1jAQ1IZoJYUvZNCkhairYlkYPzC2qy589boH6u5AObOShmbipE7
AAa4+R6XVU3NuJP7O4YYai0aOr68mUlGtoYKPlMNSV6plvtIuBIdxggqh274OVCm
ulHnXuub35U8HQ+MJqD1lVgxuLYt1wqh8mmj4SUMWdfK/BvgwmfJBdgR/WZpEa/z
BqmGPTkKzzR31piu4r+7V0UhYkE8LX6HHrljVbafF5QDSfLMnaC+vdAe30lrJW2r
r7UybMzx9VLM1Ke5twmdISZUasagrnjI4EtA4b2xeWCymB1QceUN4mjvgwNJs9Hg
0F1Q7NiDmmnfG6CwKtAZ+dv3+W8VlhIHg1Y5kvbk8nAfbPayPgB8aVHVNXEJm4eR
uFg9tDEVnG1BeU4P/rQynxJ5ys5rXUE0LJP8hl64rr81nMlQikRk5kW6X5vclZNq
1fSwQkVMLAoQ3/861A6BRDt6J85VPZY6YDTIlWEFvIW7hdmgtnSW4YnHcenPF/lz
shOJupl87IRuZk4eY9MBQOexvQWUoCE+Xv5N4ID/0WVy6Lih82lAUOqOwtJhx1i9
EN12f9yNSTVViIrbTyc9bDakvHq4bet1xf5q1YkeToKPLXusHpthmQLQexi7LagL
cmG1EqmgkgnIZ/s4FxAJhsqk8bgiYWJcV3g+SNmTu31ZGJqk8tFuOTa/I8Ls1M3G
wZwIlgwbPkMrW4pF4k97usSAKFTtG9Ll/BOmP9ZJB4bUBAQvHj/jtyGXBDrSkn/b
TJMYlLFHd/tDTtruHs9o+NmJnO07ryTq8OZT2oAHK19N8Jnm7JZCgajAeZZg7Kks
l+lhqOydtO56Vjq8sSZksgDJJDbhGVNs3pPQR1L0cOvVfyfifcE+H2FcQtAvcbYg
uPhFxCq1rNXVDGqrE6vky9bHpH7A0EDw43m7J5ju/vc/l2nW3OvikoDbGWqPn/vw
WBM2zZ3TD7mowvI+hXoKKRbIMRaRyPS4icqTo4f/Ud0K+31PCjfsu8hdBE5PVfyV
JFarJdJ+H9JlI9Xbpo0q5ni+UkT0p03xaWImuRn/LUdNhZF+OCzRgabApbeRVZ4D
cdKnLsi/Df2CAPwapM2G1yBz7Km05vWt91/7X/5anM+sf67I462rdwm0xVHgQ9bi
lgMF1WiKzULv+Duflh3uDYuIj5M3ktQICLV0oqR4OKppiQMpOPaeriYP8AnFQ9pf
hQi2sQu+0zV2qxfq/Z8JTM4npHQL+y7VUeXdBb2GjAiNC3NjCCN1OcZ/5qV16dP7
bx6oubypwL12qJaADq+MKnv7IydN1UM2GIl5Usk2VWRmv97aXpnUehe4x97IsHcC
mixI4N6pAwrgDtPZWoQeR3UCm8xYRT1hrS4FMWpIt0/SPOpARGL0HUIwerAGRrwR
AZsZbW+waR5AM3c2/Rk9AbqmgWmaAe+NDgS+ci4jHkK/ODki9fT+nEd9DpVKMxcJ
adgnzgGllhTBY/S2bVdL2SwixacQN7EwfjfHrKAaMDvHSBN1WaFYMR5/uu05GknK
zhlhsqSTMq0OszVTor2K8bEzqQFkupwqDCP9DyWD/QUnuJNiWm3r+bjrijUF+lqh
61xZtnZ5G54gKLheRTzW9sdxfprvuKQuh0Vb81OWt2XBr0dxnw0NE9FTRznFlwTq
3ubVvdAFozH+oAnFGHY1iQr8jPVamErVfnQ6KXNTD0IR71/s56K71YKcCP7Vsq1t
8FTQFUPvmfZJOcxtaB5MluiHpBDHPvYg/sAS1ec7dHR4oKEzL0CSxDgd4SudLqKk
WZOPOKM7n53Ss2RKFYgWOHRdJF21Bk7hxU7FxI/as0UNAD+sOXTw+jwu2+oCry3N
SXtoIRpBoaEci8BkeJuA8oXyOT1UGsqGdLm8SQyxGRftcmReoTdteBXUgxcKub9l
z9+UMZdb2nCMebMztHPYV3+jwcp8AkyrhRutKo8EaQXqXbBkbaiF4VegBkGEhn4N
piWw2AT+6s7xJ/lqg1BS6FnSREc11u+ZD8AgXmdkIOOWUGgXaH2WiNjfcQ4cPjjh
DlADSWsjryN2Q0R8R+EOtlVn7xehTVZZeU9iIYvoyA/Uog7z4wkdSEF2wvX3Wios
gwdeK0eza7EzSTQPSdurWfCxu8087drYIChc+RIs2kl6TcI+RLebm+gbdau1cRoF
FMbeqo4k5HPYN+sajYKYpfKc+3fAwrIUeqPdAlYLsvFzAXVP2JlAuGABU70c3/fV
7Mq+q/5UjB/EASUmzuwzVGSX+a27AqL6GCavGekdl98UTxUDBYGByYW9+wJTlFiu
dzKkZCnLgai9PBxEuEmfZPNZCQx9IHUYhetsC1HYvT8ZqHeliRFx5JzSilX5o+Dn
r6UIOA34ff5Uc4SM5b7AWP3irCDQYaLTdBJfiAoAe6TECf3AbcpkxFmQOXUDZnhA
ZmGtvrPDRJSV/E00oZJUVryK3NMz2Lj+AMS8xyAZKYiKWXoZMjYvLkEUOHXwiF7Q
vwxJNvNdBtz1H25kv8AiAZluP2cgo30AMrtoUldMV8tnz8V3j0pJp/LfMfpzmktB
08YJ6CgKIT0o5X6r6qFePywAp3VO1TYXt0Wc7aylcETJBKeGW4bVMJ2kNQLMPzcN
la7UjHdfplztRD1zv4cHPsaekjObaKTKwv+OXSwiYt4JowQDCVqyLEJOlJ2jLDAx
pI/ukV9lVFndpQxAY8ExF+jo7/Ke3PpMCO59rG4o9kVXU+lwMAjA0uJZgqbcuJ+u
SVtVJf/061Ooc0LmFM2n/yArTmJRtiDn6JYeFWb0wwQbIqqv65zpIhrCm4dRUozq
EMOEu9tG1dhzpb2mdcPRosIbBkGr+gY5fL1xbMycSnSsmMzRlgk2e0EOLhQ4sMLc
iBKR1RXEG6RamOdNFZrlacMoVFP+3IX4U4b5Hl3ui2xM6avTtyVEHZ9aByr560Mn
+OLlI/IBBJIUkVB5tQR0iLZcOoBwNWiW8PNSazY6b68hQmw9gsGd3U8/bnEnRsQ0
l8Luf5nnrpvEii3OwoGLsfTPuVxqbslxK7chzDUDeiXft6CZ/LMwLuL2Bf557QoB
GrdkN9bxAKHuBBM83NNuQCd1BpkSU2EjifKx8iW5rBYVwV5uaSTexuVgN+p2hE0x
jgt8PLtQpqe1oz+ADdTxUdZ1kUzQVXaDaSDSMOpPCT08qzlBKrlUVu1/nErXCyp9
Z7aJere0/feqSeMv+F51JX410oYQUm89ivNK6MPcaAc9dHGonJsOV+HH+IzjC5wf
pjNdJZWtOks8GBmdeT6im7w30MUQlmAPaQP3aljayEKZSM/V6JfMlwCF0qOBRbB+
/yctvbuV9Pbwk/v6BOqohzxoXfmQdvXweAz2ADjIbyOqSMZ4USQnV6raoI433CPQ
Vkjro513yGTSUv12dKKRvUxXdUVcnDgcE9V5wRA++t/V++2g9eck0IbCg8GEFDxP
dNTINfS1JOqhoiSxfy/ZjfE2ODK7voGzxidNL0gVR4iO5I54v5MJP364+oyIgSmt
qbf80niqqjAq5B6QBshNT5AtNrfeBdQ6jqND0kRKH0CR+MwGvwDfXXy5zS/cR9U9
4+qQ2QXscI2R3fIdm4GI/ZqbyyW23Pb6WnecI1zcWVraWeoP2Ky6j0UW5r7RlZIY
I/rR5zm/nIi1JBvzakTWGOm+p4b8sbSU9zIXhNLJVXsl/ZXvZA3KUIdpvZkedOUK
rTS2T9TGMTcuAAFeVo5zRKhL19ZheGym6ax//wcdBlndBMHVu1yj4Vuyay7FfOfZ
ElYSQE/il0VfgRrR/OpqbQOlE/6+MdhJsIc7zGX0J4j7CBLHrWeM8+dfH9OiiKae
IvTQRHUHXRBYjcE0K7ZajmJFjr1+AJ3ClRmY2L6F2A1E09uUIEYgzEjfktJGW0qA
zGwR8v1uOjFXQxj9/JpWtY+RvYeBg5za4a9UOUnF2+C8XqIyxdm18sRobBrK+vZF
e5AHq7hGwMdqLe/hJfge5vfb2/RYMRhuLdjMw6tLZbbalNXi8gl/FtmrBg5wEUwD
lY/gPt3jd8uGCzn4ck+sMqFQbIMFp0a6QNn7ph1p7Q1wuNCJCasKi87VHNF+bN95
xS+pURdRX8acob5pNWgHwoW2McfEvRxiqYGxdinVzVYl/QkFzOPYNQiDKbkos7e3
OzVNQrtpkxfuT3wzhJ/U7IykMmVCX222e9u+XFV0BagverNEnnJKeWM5w+t3CaMo
xEZqpvdMpkfuTA4sewVMvttMRaOJZ5c3iw0MmhOFRqtotpSo95zM90ccxFuAYlBt
r7pXCiGvwKGLlkLUaQTDPfgSeS+I1wE+xyVPZGv9FY1+KNt6yqwPuR9hnMzpUoSa
QjvOsw2Qb1IXmiGS+HQZtNN2z2QCTY9vQV2HqAoA1aanamOU8ApLOnBnYNmeZ2HU
ozusktjAcWR0ZD0eUrjA1VRb8ydD5HKYW3Z31f/rNY/SE4wUYHvhjIjehb5kPRWs
PxvY7Pp3LXw9sVvL+ifnMgptDesAyGy3mkElIsyen5rK0LDjiCA7CTFtHjXH18vH
z94K1P8+VS4Fw6z1YI5+jj/OkeAWqCmjRnz+XEquOBwPeHFg45npaVRoJ3vXi0w2
ybMH1y/xuU2p48tBcfXCdH42UJh1g26zV+zj4sfbjvxjDEbayLTwzJvRdBZzM/0K
gZnLZGElQGmEX5xP9sMhdARCPv4W+ZbCsGXAWSYnVf/yzJCE88Wtg/GPqBcgW+qU
CXXxywiPxTVKMnnrKOH+8GCz5SBcjoOLR07Xd7Hivm25LaeNc3LJ4oklOHvYVI62
8nyMYh/ksPWBVR0zNihdTZ7kODsffy/AXXmOduCT8gjeTrIF2f5AhfYDae0qCKT+
5io6Kkp53Q83LtO9u+HQIArbRSccqlJnVf4xIqIWJ84zxLmlHtJLzuCGiDO1a2sj
5okGY98dHwdrk8/+pmj09MH768BsR7vl6SCzrkZwSAaeG2n++WwrnV/thEU3+nqg
1oUQsDE+bVPIXkq+lmQjxtXPL76ZtW924U594cUsliqseeyeVM6KgQ/+zIukzXc1
9THPaLaec0hP/yfDEM/by8TVtl3ezohO6zyHHcy41gJFCAxN0VHcJUI2lSZ9ztYu
P828dGN94GLW02W4BUduu8e5ylWKdmuUENW0rhCCFDeE0zE/AAubRHo0NWdQoc4D
lJxXJzJAyDKxlb7vZgSX6W+w7c7bBj1DPiRkLBPpAWRS2zRZs2hBKaJugJ57rNpa
CUcubz5/eqqwgZ9MmUEDh/oWMSWeo/eXfaTzrEjjkb0gciWzFG77sSowZ15Opfn8
FO7RkuFplQrHXop/EovWDRG2w0rZ+VMA2gaWIHHpZlXZrFbHutd7SyzSV4vEdns3
7bYg7Yi14ap+/rdk8FH/PksVzwUpn4yEQ/WnvJPg/BNAD7xz+EnOB4Xbjj8PgViL
s7nAD5QaX1NFkj052DdIc7YDuqWfvNifax2bMNFQ6bteDWVQjNBY6HrKiZcz8Sxu
BDDkw+9nbAToLQfBBO0g0E/qT0DyHVYCmv9bfvr8yFc316X7OKaML2xW6xrg1lf4
8u4ruYzQFfi9XOi+13jrQbaDF6N+RvAu0KJkSPIzlTvv0xKJw+QZOEut5BX68K4O
0wFR7b9bW2mtHIIqe0hCnfKTdWgDuIQNbfRHwfVKgGimpmALAjrORRLIEJ5wLmaC
Ve8cw2n0QX3vw44tTPj+/C131Yw7veCNc0UvePlBMXac7H0kJgjfhy/igNlsBmYO
39UORVCbKLS2yJJxvPRW//0CqtpDGDhPpg4/MrzdNbkLJKVfZV+H5bvN5SIgfqqy
Pk428uzEWlGrb3SMvtJt8VQ/QnPZCQPWsB7D6EBjZ0cZ5DjyD+YgAr5banYi2EZ5
XL7AL90Tm14RlVSnOoxYflWVq4ol03ZZWdtxeMEeaOSWzVgfDaIAZ9a26+wKHgAk
neVySfZEgGrvfvaSJaUjb/Iskvr/aF4LocQTMtG+iYlz3SABIpvktM6ntRi8yFbN
Y0iv+U/QOOUYHyZuytZ0h1omhviLeEC536c3vJDS9dRpC0pRHO9POUh/pkLCalaf
wgf92QYqKGiRTPsKPwqxBoHFDIVW9JIkxWgVEsw9hof1LKYBN9MfHoeb51ChW7Vn
4APgb+BMUG6hAw7MqzClf1U2ojC/aqbX0Ly/ZLGxt8DEz7JrlP2EskZApeAlOOxi
TkXyWs8vJkUiihQtaDCEXa6MY8+x0nLIfgUQVp3YtmVYZYlJ/FBFyzwZmGSPco0z
mLbZEwoCjQ2OPeLObeZfOfj/FjYQs1su10ABOK7pP4PygYBQQ7eUvB2KJDfYusTm
dgNL5c3oSkqHgatwPcnSvJYPiiPnpwkd6LyqqZ/xFO6YWkm7fwe6Y6pxc7RjCjZT
CzV3p+gZMQn6dQRi1RVetfDufbTIiESOhODZC4Vu5is0+b0kpXceC9/iVwtGMA8v
+jnjp7rPb+k6BTuSUrOCGh0QgNxTyVxhYA7GOK3rJh8qpRmv7DL/Ql6VbN11mIwg
DErxgLDn4eV25I63Le22f0cCw79Vr4xRrYBbchPznWFzOAoy1BRE05nnHf7/NHud
TEeuwzxcWO5tg+kZZk/JO0hxG2fZ6kQa/GRaMJQ2o7rRDwmkXL6i5C42LrHJ1MiC
Y/WL8fjEOu+AVbDzMIoMyDYH7H+rs6EJCjjFi0dIrT+1EaXdfo0/bZ+T7wN43AB8
7zFmNVGy5LiIplZUVp5HLqaj8uf/tzVpM/xDFRkPsI5VnQyTGcWxqTg/4GB9x0Z2
vJNtXC2Dvm5sDMVk/VuK5wwnOJZKU8sD4zG0C/bj2K+LPCDQfo5zHo0ceWUS8GfK
YgYzgipAP5hGVVHbcjBxxL1usAmvlHYBmi1jyu0tBmz52WW4P2xGBW2BOYPjLCzt
BS/7mKOxReVDkzSVxX0zdL4uAljB3l4F25/MHk3oG46pYz0l+B8putw9+HyEvnj5
uLV8vmvqydN1/Zguj1DhkG2+YGRw3k+Tb34kXlIBXqrOP0FlmVuDS6g37WL0U8p+
reVSAYD0NxXUg9RyFZPw52625xyH1d6zjzojnLTXTu+B4INwJPXgJLaTGaHKQzC4
5m00EkgzJ3cOwhwF/7yXe8jc+Hlr/DlcFmvdeyilt21TqFAGapN11v4p0KqzHfrM
VtrD3IqKC89CziyNYpCVN0qqu680JzXCuL/Vcx1o5GPFuPtV/ZTEkwuvK+a47Kq0
GjeuuzkhpyIUEiBc0BOQwour/aWOGOXAsIl6bPSQn6BSBIRgXWalXHpCXZ0Tvi72
lXCm3qyAILuDn8Q4TQqLpf6YIZwAXHmidQMJ5uBQEc3RrC0huhPw7bbLiPH/U9tQ
p73shFjFK4nRpKpP74REaTna4uLpR2EuzNy9/PkhpIETcFy9aDSBYvg/1dl4f1wV
mXzUGCa/2yORXxPiKwVY/ritQOQ3lk+b/2nf6CdU0zp8H0k0TyHd0KfmGx0W0MM+
ghDr7HuEHpEkSe/ERI5RT9C7570VpNA1SVJlX5Ca7L+Vtm+2kyU9hSZUGjyTvwMg
xWuWIN+BnTg+ngVWtg1YV2PJpOZg3BuWhlgDvulf7oJN8pxaYyuO7YEFPJK9qKvX
UWlYJjvvt3KlSRF96jT0b3bGrc0K/Di8u9upt6XrIeCR0DRZDvaRpnqI3KH3+O0g
rqPzz6tXMqh1xL1PZ1Dtj3WdWugCBrJJ0EB9yXhu4L6XQwz5WAAKN1G4UU1iDS9b
Vntd7EuyNs3Dolwv8dw8CEG55wMpLNmLM+LlYWxp1WJnTD1+BUJ9z2+wKVI38rnd
my6TQzVbr7lYUurktwAO4Pgmu+3HQhz4JF6RuUAOtw86GyyjNWjgOy2/qvU/xpCn
yWvQyQjWLRKEVd7ytKptqZ0sd7S1rT+UZfmZcT7bkNur2Nf+TwdSpBBu8wELMjc1
q6k1jt7mHTjwUQ2jLnTBJK4WSpkKGO3J/mMGcfCceJskoTl6pEp8jKufAVHpqMwd
Eh7LUPl5K2GJ3gS9D/P0G6rFVCnBDH1E0aUZoIVfwQIXtKL3wgBQFJTqczuJTKWU
9JQBe3DQ2+v6apE/bWboflsUNnbaXfTCCjQfu4uH49P5g2LkjIzmR08KCzE8eP0H
O83jKmPcN2wBheSfg3l1Y7O6h/+jkr1zM9tInxfUg7RQMDpvTk1E7p5vBpVRErb2
eiupN66wqxJ46D1h0eL3bkia/xQ6glVc1ie0zAymVjsPPge2tMouloHBqeY9O85d
P4t6sZGkasq7r2M87Yg4GsBQOnxXhyrWnP1Qx7Rv56/Bnat2bSpz53WZLXmnZ2Ed
j0UNt9NjKtL0cU+cf4Xkf+sA8dKbKubKNS3Z36C+vs0yb9ODBoXSBy+JRhZDpa3X
BZuPAUrocz80MP14/dnDp2NBUQbqDkeIxViilMNwrdJ98nAQV+B1Je3YGqmaVcwY
o7NmHhPq2xTGIhNgTq1mgCCx6ZqLN+5zPAnOUlHYIN4kMFab+jPp7p2fkOFitYD7
WeuibtAgDhG4hf8Ah9JrOGW1fxAk21izNAaHQojjtHEzrYqqqEadSIMRJIZRRZwg
Vn12qxNR/21xyCBgirSQhz+l/JSRdB8SiLScvr4BjZ6juiWL99by3ktQkz3dv9s7
h7YQrfOLQBK7077PCxaQvretpkfAKFA0Btjb735bPnBH5kJ0CFT4iI1MKb3EmjuB
tmsgYyoN2W91tgtCxxsuKGrVJBpXFG9tcjcUtIwNTPVwgRAEveKqU1Jk+e+D2BDI
PZLFspuiXuwD3mWWGcGXooFY8urNdiLjj89Mq3eWPmYFPZB6L+9BEKgyZd9GR9nn
FHhECCuQnWWpYPsRHnLzVq3OiGSQNZqi6rvYGSU70KA+JORXKkKBTrgKKRnNCV/f
pN8IgovanRJ7bcI4X5x5sz/d0J6l/Rg/L1i+b43A03CMPpc/UYs8n4sCMePA2veq
C9+G2KzHZwrJ03/XwgarWBBRoaq+q5wH3cwSwhFmreCXqmREVr3t5CvIg+OwNzK2
SrrgWNB+W1zf0O7+kHms0jAZN7MWiplms0BdqlJSmAjFa4XzOKW5AYUZoiad6rQe
BkW4tK1k4KG7vlNeqDrz0XBT9iDVhojFdmg+/IJk2XTPEFxiMfpzIEENYLAUNv2f
OqHgCeGLP0ITEO5pXL6tEMhrnT9Nb7Q4tfMlCOrpSdQD2M5ZQLf7kK9ToT8XxcLb
BsTIm5VmzAzyX5hwgUzB3VLgpUcqMnsTSwprHNh0NpDH8lqE780LDbpcsn6yhQG+
jUPweIJOW3pbndoRAD8eRCBubSVLf6joIBB4o6sK2HwcNz2Pp4oiovbPCfk8f5d4
tCUKpg4CdB5OsROC9KdViwlgEIXbwGf9xGMRmhPApE+I0dRBjJz1hi5vppaq+4O5
YDQk78Ki9E2wLHv8QdUaZQs6seQ1P1uwWz5K8tS5DG7xmrBupCuigqJITGnhiZd3
jRClzaP927g2YzDTTqUMO1QxuCmMm3Ag5ud0uk6Jj17WOXVE6Fff904lrC3NHHFK
yXjqK3rp7ZQ534I7RlA85LL3yjpUv0Vd7+janQ1hwiLlp5rZLcpNsoEIPeI2a196
4jGIL5N02NoTKEfgSxlH6CXpMsDeXW9sw7L1WNy3yyoUICiJN5QfKhCcG0gP7d9U
suZNG5lr/ZxlgFLte+6XQNBrYbQcNlWEZ977fisSNVwEtPu0AQQu+VPjxuwxf8Oe
V6UzM9/9CwaoW4dBYf9DUyRRDiy04ejYZTnkqWB95EDBJoqA7+l+i9VeW5nCT9os
GB85UnZrTr5Dk+3Rv8D/N+HAuw5ECFLUkluKlBDK//KfbH9kWwE/D8NDiW2hXRUZ
S0gW1kX7qkeIIsSFt+y1BrA3U5QodggwwwZvgYsF/DPCqfkUeD+7Zosa+uDFU4DI
aIU69TkcOuIUEZUJpzitCGh9gEEf5URKRt8cLHECrEgjlohMvTPdom7Bo9KcvgjH
Mo6m4ZHSN1klIW0mzjXUNWuflVkRR7IP08f3oJqXK2DvVc5BvW5Y2HXKJINQTUSV
5R8o4magcmh/wvxeNxO4Yz0m7Gc26gR125f+q/6yMj0QOJsxw++6v9vTJPPvA3NI
TQBiiVMagAvrmPZvZBERk3kxeu7mMrAOhGh7dw2LzeRo+/470iL8Bpn14N6GAA8q
SzoLtU3RnCYZGOBniSCCrNzsPpX6AXjZQRChOiWycwcvd0shVYRJ8s2s1zN13N9M
eVEoZPoogjgHBdDN8TcCGz5P0LLUCUGlPxxMvzUk8tnjbAc9G1GFH4uYN/9jpliv
Njs+a9iOeTNnZkBwFWKZplOFx3l5odT7WMWSH7Je+qpCBxZZr9GY+eNXx3t/T9xL
el8kc4Ozp73JFJ+9s3TekVn9MjkjvYQnXpCq+eYPlrg9umjFBASm02lLMQgX5j7G
7M19HzpvlbMEhOhkRmKCKRJktzOery9khyGBXPN3JqTWUqsRTELjgNfg3VKzYWrb
atW4o8DaYhKkcXNWjGEiDnDOjp0LbJeniKddvHFBoNnqUkqrMU5woLamEVM7UYOD
cyFOaH5BX9HIJNh/n2IIPim4e1UHU2V0Go6KTpTaRPp/hE71M4eDHryY+hhJLCrU
8Qd5lBEkRw8+05+dHbDu6qQPM6UYb5f6LV8ctgrOQesSr4U3mk4e7aCi+qLrIThz
YpcT3DrQPzMoVuffyEUrToaDINMA9eG+0edOHr5Y3Lyme7G4VQ97cI+QhCZvAkAU
4eO0pHLLcadV0XRJ3MNjn2xtWcjj0bVgFvEYklqyb9JVb4fFVWlx17McQIYP4GX0
ymvH1fMPJC/TNun60PnFSMWiwTkpff/V38kcHDt1V+Et/e1jo2omcLF763c7AvaG
WVAUV0L9KlAlrkVxGcOlTxr53FAmXWU3zzJ9f59tRGdJfV5B5sXqCovA6RGU9kHm
dDPR6XmV1+Qh6AREyHpz8UGLxTnvTMRZYTmH9SSoH4V09DDNBiVJKGtn8V1sLlG8
Gimv0LQDLhEQhKiwFUYAxcssBdUWs2DsFmcNuhdF0pl3ecIkKMgOoUIx1DlBP+Tb
GU8V6Rj2yGiXeZzMTe46tDzMP+Cdl5PKcsp+Ir01HtvdILC2FFs+TWmAMPYLArdU
eOVPejKe+VAHVOYyN3YqSvVARjx01Ciu2SOKpGxDyoc9xHFtLbrLtLfH1ScdAJln
n2hVa9SM5MXalPKxK9kL1wSuJdf74IXcZtlMmtXdqJdcjWN1b7XhKM800HvdgOr3
+1HYUxb0JIF7L6bZE9eAvIqO/dFRFSV4/Z6ZAnz1qI8/fr/NLrMKC3wPdCnPriiU
vVnZCD2apu7WwrQ7h1wLly0+SUt5y2bi/wgal/SIYlljYTwlYvRrlPCbI1NP5L28
xJUf57kMc6w7xF2Ts4AaU0nOKwj/BA5BDKK8OCluk1p4PNcwRuwOmVzJOF3ijriN
OHLOGoICjyNBKL4ZiAf3TzpHFx9XmtztzQ39xhKrOoRTv1YV/Acdxd22Gooit95t
giv+V3yqumgRv0tPhmYjEjyyRrqyQniJHNLMgsgr92awakjUYhAEyKOWA4ru+rFv
stVDE8RBTfApnB29uTqtVoX8kdu03zGtTwE9TMokPSfXIqVWpYvUt5XDL8GNUeAI
bXo/y2WdhAgAmvzEO3hNe2EK7EJ2c0n7Frp+WM3pHSXFTHYcKtHvCSTD0G8cWC8f
Gytt7f5DCN5gF4hRo9EIHSQRjQl+3eMRwF2b6xNmg3y9Cs5Qh3CQTn1OsQCIp3uP
AWedksySVQA1R/OJr8jSRFeTbHC9yBb92mKnHfLNfm907NtI4KbdTEoozvNQbF6I
3sn2oS9uQAbSifQ+AzoKn2cGRG/yxAKqss3crubpDJaQ1ZWRC8YJzNhU6uMx1/Cl
r/Js4sBXlmLUKwybaXzijXuoTV+x97jephtYXrbIi/JjZ9ei7YRczJKWsIV2YrF4
S1QuDW5hz0yS0wOJ5r4YssjIZvmGTQHAkcL2PQi8Dl6y/ByfAXIF5QuIpptay+xi
77E421VnMar/6SNXvR2hl8vEBfW3r8R9cKbCAcosqRZUwDebIMf38QQ2UFxPN5tf
54aQfX0pzzZeYSto7kiMTqrDU6EKFgsNGj/UlFgp/dOVgoUKg+IIQOyiS/VF2qZv
JX7eOkSP3PJin32pt9MMa8j/DnNLsYeXFGvGJBl3x69DhJQ0wISplJkHXlTNllfl
cAST8EE/U09DC/TZ3MV7kCCo3Ox2/PPdTdBcBXXnUj3WrMlxZqnkqhX8V5vriEiV
21Ts+8FOqGTpCoWmNde9x1Q60wuEGyVl82lvuFsDeI343F0PAzUzZFMwCT6lsfo4
A6FY+zHkCQkRoKEuvoqRgfz4Bxatx7G2wxm92vbPwUbonCcUaycoITRptd9U/W/4
tniYiFlSAjxaHYeq61EyUwyvrjIajs2vXlguPWv63rY3iU3GNeh8v5jNaK2LGN6E
VSJceuWxRJEWVhFNVth3PmQSPyi+l2vu8E1trr2jkO8AaqrFY0jNLXcP2kMEcEQT
zRYOz+soG5VP9K6BoZ3bvVmEeuvmGUZ7+2hZBaK0/uxY5G6i0WJtY69pLaydQkJc
o4y4agFcmp1BdEzKKM5b7xt48gxs64HU0SbJ9tggjsec1sJUjImjdluRlFdbpB8Q
YOircBp0iMr+iUWkIPtZZC6kg6idk8HDAVGZQTyPQX+dlpHv1gZ3vojWW3gi7bgz
FhopMjvpt9JF2floJeR7ajqYYXCCDAd8+sGWYn179K+HakmKNckRJ34BXpexasIP
pyakqQ+tL3zdnXdplOu2BZZWVO6SNusR49fHDYnBkATuS8CAp7FB4gk0HUL3Ct7a
IgwleLmXYTa7saMSDaa8c4AMFLhls/WrD2QlMJh9MX4WD4c0sNX2akByMV7nHxJ9
Z3dknMmjdVCrKuH+uYYItp/zc9f6audNmQzNksHWUMkXfZ+fqpCjike2WmIvsxtn
1p6xrHm5rdZjEIJYVR1YE0asAoK4mwNt8mtMZWsESdPdW82Fy8B3Fs3hnpi/cXqm
fsuyG1Q5isAnfOP7dX5pgC4fki7KFqH9kuzpBJYJQXN46AIehteZvdL6Zbe1w5dt
67uO3RFNbcmv/iwEUscAb2VmvHbZbJuGEGW5wdJDVe3jI4dmZ0ahc9VYpFiFUztx
5CvGRZTKEtI+mgq5DFaEASqX7/hy5gR00Z/gohQzgcfhFnDsDuwj4zGBYe34o0jX
4chdFjBFvte+9TRCeaOXu9FmjTzD7BSMShmGGrONYStlhD9yW4j+7JdL5V/xFe9o
dYBCY/KgIim1iOE/VxNoeWJkPfKJ3ydEgpb3Rhh8PGv2pJWhKopMittKi9NEVsKh
hrZj1ajDClfOwdzpA7fCRuLI/dcoMENLUxBkRJ6BqLfq2eMCZqI2k/QLaMrVeOJO
v4iB/6q21z9Z1WEuQBmEFws+QkLW3qiFT10u1UVQIJBmtOOzUyuVT5leYoIJ4sVg
e75j6NDMeFFHUBRv2NXVbCEFed/7DOxOhSKUKCaRVI8jR4G1XOX4WJYVfsmE6X/9
6PdCoKnxFbkm29smQAKbm7VzOqbC3ibEQX2eIhPw+ix2rXFawOsFIU3DSv23d9U7
MeksvMhceuWzMCrAOitMmS0Ow57j5wiF6GXm6vCo8eit59x0OkC/pLF1jMHkCbUa
fHAWkA5XawHjjSeyAfKJpFVfutoKoqXLbMbqxl+01B7AqYcL8LXZxMNpm0QlU0bH
S8UTQnPQElaaKmBfDMZUEFYqHxCfNjtBjTHJX8pPyYpYcWBPeDkoUtnCzYRlZR2e
DPUlHLbcgtmd3krHWJfuWcw5SB1F1MwRdk5GOLxLHk3RYQW9RbLslVfyWQb4aP1x
fC229/hGpuwT/zMvzdiaAS1Bw9L80GyYEpANJT3sbMjRR2CKVVCDKCwI1DIXLmV+
h311uQ0mC8RCqRVAPfi4Mu62IKi6VLQodvuycm7zFazq8qlqZpNRTdEryJd8cnpA
Cm6rCU3PnZBRHYKPsnP494wZoPOrGNM6zzjmrME+x7+I08JT9SC80yydfZ93YTP4
9tf8FB3XDhrQRHbLsT276UDwgoY69orQgPXun/Oc+mgM5Q818L4wo/K0i75xxhkC
wNg4FNJDM22IYrrcxrDJ+n0vNHFIatNcI0aDoXmLeJ8IuwKRkrUFAQBGZ54N5Qnj
7CrvcjXbltIzV04JJPvwZQvEYCYrCUtuY8bfrN7wPEqteUp3HPyudHOYnplMaznZ
SBSHE+4AbO8qIVN5ssspnZ5p3Lvv4usJPazrkTh8w63upujEkVjrfwVyjaOYhx7J
yokX4cHmozyGZxNWBxoO+bKyNOWLJchhdsSMIra0B0+cFaeYOP0bW1joBIMqQ1e6
GQlbz70yZStaQWR49OKvj2ewn764LF9g0UZdFF130unOjZ3n2cjcOheOcyu5sWcs
6FRUATJmycGXSXxL4xEIv0GzotOlCTkzByf+r2/17en8ZO7lD8AXC9PuhuX0c6KE
Lc7/aJj4gJ3rCYdVBQwr0zQDbiIVq1TLCQl4ofr57w/KMMJnZSa6KhBV2A2ZFqrg
b2rsORIf1GUIsBfCFk3eHUNTSwAT2tXJ5g5f2TPvxrw5g7BhJvdrOVl+afJrQ328
tzuWfzj7aI4Gcm0g4/R2Nua7ueowEXK1/cZuxskeHjFGkZFHRrMpHcQ0REmJNuMa
tl+3wAs2jEe2zK5HMqnNGf+DYRQ6XqoGDPHK9HtJ6lVBR5ON3V6Vqg4U5W9tngxO
9ViyS+aCiHhvslHkKuD8ILNhj63UCio3YpfNnVQJGoXs0LV0eMDFiLtlBDNa76MB
ugyy2enHP7lMKRRqw8KQV6FtNKxQWOXwNa6B+bA3Kum9/kUM0CUmakCucRJzpUGn
844R4tMzwTyPYsvM0ZjKdJp+DLvtNUgJV7K6RHV3wi1ageBdqpPVrLoDPpqiTf8k
hP/Um/BzeRI8MKL0QKYV9+wOkxMADCjGum+jZLqFS8DxVPzQhXvgHQ2dIV218hN5
e5SPsR+O1XaLO3aJcPLyxCgTEZcIa/XxeK9RI54Ne4oZJlUK5o6a80Ler76PtVTG
9ZzjNp7dnjCiFS96SRnkqPhXEpwvz221cr/S9QDscXW64fSlURXuFPqYw8daILiK
XyEFy8HjkROMFKFTRENQoS+k2NqwzWNQjFTzvwehEa80385EMZP3vPC5GzJouYUZ
ntAMc9mPXQVJKpI6KHUi+2rVd1a6uY9GAFI49mBDKp6N9Y/sp+Zlbr5jhDWReCxQ
R1w3pI/4qgRLAiDdij54pT/q9oDSNV74xzmbMijaxLZWn/QqLLa4WPySb0wAlW7o
ah8f0zDNdnoEu6OSVDysXtLjBEVKBzC0E/WoRpNut7B3AcoVyHBemAQ17wQ4g90k
FqNGXwPH6w0uenQz8RDMTKJuxyGviJrZhGcx9DT+I3GOr8HsqFZ1vzAtz9jfOrCD
qA3KzvQwgHHruyz8pcihH4Ax0mTi7UEs2ki0mvV/cMl1C8dcVct9goOWlOuA1KLV
nycAmCvFVCh+AIK2dNDAGBbE1LlwXKaqzd+YGk0vBb21S7RdZd6hykRRkSJ0UWc7
2VHlbTFOGLhrs0KLmWl5z6iHKBxldSZ1jS7ngeJHD4e8PLqT2tcyQ5zre/j5HDju
rvXWgPIjxr5nF/rEmmd5UVrfPHrMdYXZIAFLhMczN2nidoEulnypr0elUFGCTFSj
piHCrzzQFSFnruX9VxbT+RbX1mrG6qdL2OxIApB3OPpKrLFToMs0DZzSyjLd1Zb4
WThXAb8imTrZFk4sqhcjY+SyxSm41lh4R+YgaedTm2NgaaRQh2F4MMP3jDBEr0pb
MW5PjGOgya/SG28f8nX/r3beM75CmHrpbM1WCcrAC82AJ0iPLhBk86nSxsAWYISd
3skM4tAGGRTMduGK95zjLAwi60YrHw4nieFsPY3VyUW2SprX/Uxqdr02F0gzwFn4
WWFyfCqDiAjSHciT5IoBdDmDIDnPfmazDIhc6PalPY5Mvlb921ggRJ5U9pjYlmlG
1VXVd/1AOW1xx7CLNczY57jpP1cf6ta3CquoSZFMM1vHmX0f4uHmygRdtY5fkcOT
tbKy+uAekI7DPkN8Ji3EmCJdPPqUGLxq4fE6tNtel0mbxIe+tTp98xTSWGbo4y4n
yyTRRdcfHIGDO11QykBO658plJStdeAtUDXonCM2M228VZOD4vnLPn+9LAxJHkQP
MUyMw0mbfsBMxIo6mHQD5qbrt62nRMMVJIq0lPv2HUcqSpDoY95+YI0hDpOmcW6k
t8YZFAVWdnaj59fs8x5xU1Ovkm5b0aTYpczR56yqoJlWLWcWTuJdpojkTEKlQAt8
yDQDnYlZeLyR6ffM0/5KbDQFuwO6RFvVaIVI1+LPXHs3Q+PiBoVI0TkpmCeN857a
cqNZyOWJTXAW4jT6PHJ0MWdrgaSpPAVUwXtZX8uKez9VcQHOs/r0w1EweXVWTBwA
B34ac5Zg8OeJ3r+JCRIMRGhXPRsb/wg3bp5FIRGEt8IBKuaZnSNnP80bo+NIzDCP
Jx6MIdpDG22xf0DVCNTgf34AVxh7te9TMmB1ITx3qrsCHlUIRHzPRJ1XjmWJ/A8Z
uiwnV7+5mdToiWxBtatHVmSAFeUA77/g771e2pL7b4iKJLjriTj0W4pnti0X47Xy
AjJtwJiu0RxdGdjbmVjKlyqSZdDblHKbllP86cBImRHrMdV4ap3OskRwD44tOxY4
cXybFGIgYhq5t69lsVFd8QKhMjARnJBx5eFCElkCoe1zMwsG7xH5mus9MT7FNEFx
wOjWYXJRFB2DoPQAEH7YQYX0t7R3M9n1qC84W8+4bRS/WPpGUu7HD3JSy87n3+Qq
ceZKhkG4LiwcQ1rwypXVsiohSfvgV4mrQY8O+pBDN1kPyYOCqFJFwj3zhYCYSTJ3
b5/5nUcCM8QxpvAIBjai3vPA+8vS89Nmtcp3nw8RZHaZXqaDmjArhIB0JCPB5AtH
xcf1lX3c/W4IEAaOgFxSfMNsfE3bPOAcOyriXUJeb2OmH4EgZajZWi4r2z1e+FHg
w3A/rIUs3EofXAXmmPPhm9nlqaj5Z9mTIgdRzNfNZzJuzT3bBQBrqKNbHQG4zmcW
8tbPgS1/PDHsWIefJG6lv6UKYMsPa/TcEdy9pcZM1wwAYDjjSOZ/1yFsOVB4Kfzh
a/L6mLxiSu5cuj12XXKvpOLg3PRITly/CT0rU3UXOSINKT4Mv+jaH5qasRx95RXK
zuz3geskw0X6nl0AKHpSFBAReJx7sj+9TwKuA1RTTUgEWMrOeeOhWzabfJq8a9vp
5MgQ09lv050WPcJYeDHhejtTMGc6PCyTO1jQuni7Dd5NvYcv3bwAftKzyok7p0D5
JeSeJGMdeFUcmJ84Y6iBWGXMaGxYDLTJLqqb5+LcC46hmEqwHIOuA8+zJM7PWUls
25/egj4Ev2UkyUxiyGxApeUR3dgJXAZYJD/FMbgSs43eLiyg/6jT9JF+RZJN5TyK
BQE4lUYVpS8qaX/jqgHYBb7mSYtOjRmS3Qc6jIEHMXabHp6iA4aw6yoHPWCkJKFr
0dMuRnqo+LIe0UBMumEVjtPscmBU3yB3R/68t1+xW94IieJJ+jXS7NUUAeCFYVH9
Tv3vFZBiV7McKSX44zeaG5UHQYPEyYoEQ4kOWbzzXNrv1irAHuid2UeenCVrYPC3
B17Zyfaq3rhAnEYR+KJ6o6angCgXxf9p0rPVq+fKq+PLpcZ82hfZbQInZWpIKDDS
gGJ7ZI/8x9jJHj+KyI7UGqjAsoZFATHX/WF19GXjJiU/A3MjYYP5kYW7zcELIM2m
2rvDS9JJM5Q+QMNGf0JTIC0tKR3lIrsjiPGOSVkDwuj7DPkIUPRksZUtqliqSI8t
srhxC8HaJEwXH1mpPqSwmfxttgw1sWBdd7U13P1Mrdt9qAwA68ACJsZpFGjpmF+K
1bmudoSuqdsEGgV+2mh1hj8GkdqBhbsgVl8o0SCHotsEoaneU9Kx25UHSlVyMjjP
PLBpC/J1FY1Ko6u1sJ5nADrTNNk+3UEt/yG9zZMm9HoIG8TjIB8wACz1RvfmYL2Z
n+O47aJ4/E0IBDCh++rwTJj/+KFbPPBP6u4BUwhiBIII6jgPYqN22WyZypu20HFY
S9s6vaJoC+VLyrqcJkRwQixAnlb0B8GPrUMwPP9DhNYh+U4eOcLOsAvo78ylHGZj
HzpCkFATJweKDdLq3mtl4s0BVg+Q+7qmgfKGAk3a4E8aKvgbqPHLA6/GygekbHzM
VpVJCxHx023z8kIlV+VAmhdx/MZLNDknMnsSgrQLE/PvWs42lTp35/IXanUTXVPW
o/UvATGbPrQ0TYsJEpMX9+zdtUjnUWVBvhujYS/5IMAP8EgoNlZbvHUymTSWZGMR
u8rizqatM6Z5+OrPImKkF0/zslL8nxj/eakhQE1gkqRmlfqmTR1TeOMagtpaCSO5
lYQefiKuv80lKIGDeEU5fVXXwq14DAgqJjzu8/r4IWY/yM+gRLHjgea5B1BuE79A
P0fKxmTGctqjHfTf2618NZSOmTsrNnrYG954pNJxll8DlqF1rteeROU51uf7WF7Y
5U3s7EAQVYuRkieArf3vmzSLbpG9QNNh3Wp3yMbY8qiu5kpHJdq3YfOzaqpfP3v/
aK28h+QaKFsLfLXVb8lXuY9miAq1JHSMUGlBRv2ccTUxTMVf/cpQw1UbFiS0yRjQ
CzK5Ew0+rKo6POs4S4cUi0pZDiabbLwGKfubQTPp2R7vka2xSkOEEdEc2Qo8ZkLn
G6PZoZ1nd72++P/Cu8KX7hTbsaqebh5Iaps3ifL1w6ybasXDRbPZLmSBLdZvbKBm
GD6AC8oW812haL+LfxAc2Jh59dB3SBU2KstMnthXD79WG18YfFrLfBrWItkBESgZ
udrLFYHoJQJnTXZ4QboAv14XH+N4uL+6imGIb7v6IMUiZ56/krMSFHiL+Zi+lcEm
7saAwg2m156Fg80pApimRVIL8Iyn8D5XIQIQ0vzL+80gAOI6PaWDHgMYMiJzlLSo
EKNz4IRQSvfDNmdIYMOArV+xUE57MclSRI6hn3N3omqyOTP7nhL7ghx5s7Rb2z0C
/Js1kD/Fbl6HwAZ3wKAQ2vYEKIQZRcnWoI8sLNuh08MF8Sfuv4Alg1iuPw7LrkiH
A6N0qvIREuJV7B1t0OTZIrym3K6Jdrlor7c7X3RGxGMpqd8WWHdJKbUezrVfTnwo
kZ/GBbd8uF6/gqUKfNcyjqvYtxTvYplcmhGG2C7k9/3dd7r+qVQXPvsH8ZC6++4s
dd+Zf3S8V/ttna1XU/n8gcqKlf8HP+WfVuk61TxZxtSfQLaGvEFZ4AaiilexwPgr
PtjUr3vRfTDiOlGTNr2oKfyGGyS2hh4j3EyGu9KeFfcEHFSL7k4UAH5YfN03AvTP
I3HQ77K0Umnnh8bO18JG32C1S+CYfFP1tcMg2grv6GNv6wPYZzCqMgWCc0iFDLKC
lM63jc6eGOUvf6sqSMhkqvHhYRoqdvvjmo4nO0FacH5SYxaaIVvSd323gqIla/i+
JM/p+XZIpfu6IWIp/h3YJVp5+F6dobX1YX0ydGM5qupJR4trw/gL8KGdWY0S7zhN
KIzernHuUSS+k1RjefbTozyGGb56vUTbGGWTjeaMQSX5oV3grdEP80B5ho3MNHgH
V5sYNylkyZWFoy0fj2N8mOdwTPzzfKTpL4JXhhQcsHKhNVaM0c47vBOx59pvgtYX
1Y7JhVAbGIDhufE5xrVZfwy4PYbn88xYJt4NN1PiFQbFtXbXqkYrwVPMP4zbpTKK
zeaGwz/qskrD0+x8xXYQU9nI+nOY3jn7At98+jlt/xud1N/ZYfljdZAlfsqZti3p
vlJpXQMI59NSnvKmDvrRwLocnMiezNtNpjuEjXrHnDn9zP0FvPJ768+vbDvYRzvW
RHWlSaaWt71Aeuk5JqB3RmnyNBpo72aWKvuZfPt8q6zKovhYGudkGmv7fJE4N+Yr
2D2GBh1K60O3Rue0eiPw7m2wsgPkER08+zonLhOTOMUoYDp/FfBEeS2cMyxI3Pgr
YZ/VmtvaptgSE14QsfZ5rXJ1pOt13cqirv9+tCAGkJd/3SJl5PEY/FBFyn8GIyv/
RZ7bR6oBBNVZv9so6Z2mqn6r9VJ99d85jQQ+d3YMbhe1Gt5+gu5OwPLAteaCCQJs
p08cQovvVutH1PvZbLkCRykBcxLpVWn0+3Go5JMlnOotIbof0EcK3wZXCaivqEAO
ftWwoLY9NZ605FxkH01DTP5zmxTSxE7PjEz1zv11kT9D/wcu0y9mEX8+5xaJ9veg
/LJUmJIzdgefUmtP1ezaPmi4feYHGA65uX8Xaoq8y5Iv8/CNaqNcfOC73oQ2t/dy
U3wRJrznnd5/NTZXRiCC2dFgk8qH30z9/N3SAOCv+MuLAYhW/y529jynLtqizhc8
GgcUcfATwl7lZN/HD4QdDIA8EvmBWPMGe2OXDqBRHyqRaF68CTujhJrdFZAb5gI4
nrIyIDSyuVZAGYHZ+BYOkayPrqW1vU1Ynt5FE1zVJ85yk5rVIltBuN7sfDBn4G0o
tYX/1/AwKey5M4hSwqzfEk4MhmEUEAkN4qAPsAJ312/CzSejFKeMvzRt8s6SI7BY
KV7u2o5koLCNfLSrOpEEsDi/Qpyd0SMDJbFNpEhdLSxcBdJEpqEJVcldCCnjzhfr
9ls0sFu8qAjG9YjkcN6w9Ccc+rMX70xYXH8FwlUXxoNe6LL/NPmZFxZ8TTWasMtZ
JeXzYmHiThTB2UmvXN7wZrj5cdXYNUmUp5wTddw5X8Q0ICcJq37N3LR7v569U6TG
JtD0wpCNo2UtipluIPUBVwJg/5mvJskySVMlGfVtqfBqCTy/IzH+WPuDtvEF2qHC
9sc1znNG1N4TDeQ9QB8PHJf+F3TF2PHImV5YR7ZSnlsYz1fm5wZhm+uCNqL2a5K9
keas3oIxD2NGzbmGaKaIXA2j4lhzhQQuOtUnl2FTafZ9MkbGbQ8JyEMcVQdQiW3m
/hw+17eI25CdZMy0X+O1A3/G6649ECxo6Ryr8f2Fx9R+4CCtBUiuYlYl4rzNBIv7
mp20cCM7GiHm+/xtZkO2oXquCkb+oRvR7sCIRzqD5R+OB6UiBTcd1Bbaws96WLz7
xlAefm1zU1xdQ6JQ33nMRpqxscBNpE08b2f0K1XwXTkFahx090NVe6/Jz1v4DVD4
MQumlokLnM9f+JB85+IuZR/igROiNcI/BFBoLOdDbXTG7+FQFByXIuwULvM9/EHu
9lZp5AnZOVXDOFXjkgLbIlqrD46CVNV36aZfaaxNjQzliks0tLuGQ/DaED0ztFWn
LE31DSCWXvKwKlO81fCM/447SX1VK4807v7KHq4gqYbAKj0Wac/XJwWEFJ29DLQW
DheM+CFxJrq81So/Pdy7u/qpctK6NZFbQJVDVCKcS2CPhEKWBqfB+v0Gx7SuA6d0
IiV5xR/AWFfa+csi2gcvowkbD532kgkInLKGJOxKyO94aSmrHUNTvt0jRv4hlXL0
56xuyQ/AqmFseNx4TYGL/f3clQmCoRJAZzu6B92RVxxfmpvfMHAtz8FskWM4mbIo
yCB1LOPBoNZP2Gqw2XDr5xMK8CcRZt8ZB2xyROcyDgqGie558IWcin5ikpNQJtxP
H2kbI8UkK4xkILg2ncwZq77wnZ3Uy5OxXorL6Ifet4EINWM3CmrozP7mVoYkNHln
4cdtdV7nzGIHp4X1/lLyyK/PNSukQ5nVKbcDSRv6H036vMMLNrIBYk8iXoJEyKiS
ubW2AaMR3vXfZleiWoj3/toiOQI4gxBvNvYN9Jjj030qfVfO6Mdl6LhNZG7xFI8m
SGEMDI1Iv+C8Ulj8FiU/NTNhfrjM4wX2ZEW0jxPsOhRJDvYH2tihFbSN86i17Ula
QhKiyM5ClIQqWVPdz8o4VQ8D+F0/yPKhshaqSh3cO878282MUER8edT8hoNIiL8n
jNzWIw3PnNXEHXvO6LMYhpmcpWzFYg4LYFmeqMGcD2l7sFTa3n4W0PaVJXYsPtWt
x7N9WMymO/BJ9nqcIM3MvzlvXzb6bOKXV4szwtDDoaj3oUK3gpgpflwRS1fyB31/
22QO6877h4thTgMA1GII4H1Vd7eisIWDy459QFHuYLYviCGmU4kvLXM7Vy8z+v71
eJNAWkuoQn+/34YMPrjUEEmSc6TT/5hrmSvx1i+6rusao3O5KK7GA5MxIhRDFIKy
XG8ACcWjjrgA/qEM1Cep3XpNoClSuWh2a0FnjE58wKQk/mVb5X1miysncBT2+orl
MrMYFqPQ5rrgmDN1Od47cyBs+LUtqy7zlI7YZa/ZxBngw1xtTFMQYKjY2r4FkLB5
NCKtk+6bmiOz38tMYe08GKOcYHUtWwHAKVu8xvD9p+F2h260jKLnU0779fr4hH2z
UWpL4i/4Hm/f69vnS7403XfJCHZPPi7sOckoh8e7qhbtsUIfOElCMO1COliNk7V4
wIpffCq3SBKpCtDav7iQbZH9azJ3C/Tp1O8+ppF/7Wvcq/0ZPAObq8eh2+NIf0TV
L5NDTiYgU8Q0x2DYv5p+L40HNQ5mupAy+tm7UdOG/u6VLIwjrCPtPIBnRh1T2mEq
M8hGXwXbrOg5Aokt5UREN1rXx7+SLXv4q86340C0EwxOssAfjCyo/hwUfSgRj4Yf
WShvwJppGZp4C6EbGM1Rtj0GS9GxgJvgYUNuyBoY4yNrJu66ci6z/HT++mlS7jV0
cmaqKhU90WWPw5rdhs03khnxZ7Om8m7180oT2DdAQNvX3/h7zogatdeoca9MWxem
gmeHqdm2TD459SfQV3TsNeqaam0YN6mO4RSn06PkVQ99K+3Lm4YO4I9B/S6ehNPd
sQRQh0FEGrLhYv3tU/zSfvk4GW4xBy9n8N6VjQljBi/wJTMXKBtlRVI8385MthKu
XimPg73DCU1QhCOApVI7yKfXtVY3t1JW4RaT7+xdwDGTuX7bsfZ9tEfkJBC/WYeE
Q3L11lE1DywTD2XnYiqiRIOVD1AJbfTC2TN7wa57QPhQrqSwSGGJitmzEbcoGZ8G
z62VY/BU59neFSNUIo2SdDpk5BghBmjc7GWgyeo/43srQ+tnhNVObiNVLojZL14u
rz16ZeH9eSfqLRfWHyIxtqvmMb0c3H1wfNa/ma5D+IsORHwQl/4VlPtIroW5lwFY
Rq/4BaaubGPQ5NRq+ldWAnH6SYsYwz7xsRApax6r9fnuHAkRy8yeYmyEGwczygvf
1zmQdoWEiiqfvuRv6TepkF7knnP/P9KmyaNDmp6ifuZLVhIiFXhz2M5CztSqhVnd
zx+pLaMPjc4ldOGRvIMjIIgUW0xq2WaMxTLpNj7OYMgDTZaeGvwWzoATFQjtAGWJ
Xzv+FcmQFLKn+IHiqiz7gX7xEUnMpFe13tv7uLWbUBRYGk23c/NKxS7Mxh6sPcJJ
aBSte9uo+6F+5/wo6Qyi7fkfv1oxNxLL1wN6KohG/TsJ5X4JleWjdOLe+Vz0m6tr
K3yOGbpHHqjvpOKzkrh+yTp0xSHV4tp6M2EFE4uMmSoew0MRVgUxmNp/2z8rmTGC
bDvzgCDqILT+5KpNwr5R21EaUvRyXnuFi0YgNioJqRA00pDK5gEQb7sgEHRXWshR
6xGuQMe0DvHZ7YTHGZRdjTM8Ui2Rz+XtxOB0hHhYRM8OZnCCUTcbcsbTIeRno7ot
yylcYeljc+0T/qgwj/OMCv3Fo/pRzLebbfALloJh4thNnkC8+ho5/bLqMP2PQ54Y
bLobRM7gCK8Acvy8MZAXke4lslUj8k+Ev7LRHwh7MQvKWcCIN/b719JyyIwxOM2W
9XRP57aOgu70sUQg38lfFJn81bWePj25MUGHuoFmaWYIsAtGWT1VYsYZ0Ig0RWm+
/M0UO7XMTIp8LIKjFpMe+XAP0aSxeXUZ0k2VqQloKq0+BeoDqTkzoqPmRTVo/x/Y
pq++sTOU72UqPu67G28rgkOKEK9VC4sZsSaieVKVz1j7v55GvY91jezxicki+dVn
VuSjz0VLPwY3Zc1w1QDdC0dH0r6SRrTTMsCFyn9MLrMANU5ezcfvgMgYWFITUtot
andgwSPq/tX6WvdK33RqlEUDKZ8fA5OgFWiHVZh9U8/u/S4Dgs7sgucNrQvoeNwB
sARjsrFydZ/vJ067OrfAa0Ija7SzQh9SNKekuzYYcfw6FnU9R6KysM0ySRXTEBAg
N5emJt67hMnZuS3lt6341cvg2DfcKm/afBWPZ2aG2xY3xHJAfAi0j7tTe54oAlfY
yU+uGQM6eGAh2BdVJP8el0fwJf9W9qTbbhh1Dkj7dRL0DKp2wrAJEeTHmCjcTWXr
Ys68/Q6SZ4rLihbR9j/V/cAdC20Yn0uHij1F9rbZ17kAeBRxbVUADzyyLBF0wlRq
ZCNBTe2tzu9mzUoOti/CfnfSBM5bf7Fi0oCUR19Ofxv52vG9H0DPv1CniACp1Pm9
JV5KRuVZLa5ovxHW8HqsF++P2wZR/zcspBrN9inb8sxmi7g8LBkIjHTO8SAs/N1p
E4VAwmgplXLv2Z1IYXnIInGV/lx9Mr9w8zUTcCvyGAnOWZUYdqaqht3WWQsrVAQ0
I/U9PYSEV2yDDGqjM4kGQOOrDPC+WNCEGLcDUSM+M3xXsWpEvqiWawtKjD4itm8K
X/BTsVMt2nrJDnUkfFgV9AyleWfcHlsw6NnaFnHOqMD2pNHUtaUiunyX2TfVbr4l
6X8JR6XGfBL65bZqNfinBcjLktxeh2f1ojHwmTaKA/tu+dMYL1E54B3D410lsvQI
y/vLs17T8G8AUkN2MMtr5AgiySdtnNN7Q+Q4WIoBgR5swVjwNVBeakghimoM3gG2
yG/Vx+qWfPO4XFUl0kljtzZ8Qto31q28uuj0P4MFc32yPWZ7NKzBABfHFOryJwHC
oH7gWBArCvJHvtjfVtzBFa8EzpbHxzTc9vchu0dTsGwrdxwPgUF+SmaFhi5+y9Wf
D1sFUhfIkP4UfW48MpGpU+k+HQChnvN4n6eB+96UUKdjxDuXYJanXtiPY8nRRx7z
PPY0AcWf3mxE3MkYJm+KQzVBE0YgobfJKvMz1uScUNgbwv5JaoYiqBaYmAzycJCi
k6Vl21u5VtRvIrUstc3M7x61ScrvUG/ho25bGXHOq6koCp16lqWbHuy9CEquHLnr
Gv3194trktDTMUhy6aUxkH+KoJj7C4IEHbgoRp+J0OO3iy0KO49sT2Q/QxNUoScX
WQ49rjGcQdbAZD+FwSDsgAZLppvVmw8UDvxgUi+H7oUDs7k5kRzqLeUWuAxZ0HzM
tD2GcBQqb0pPjt3XhyRcBCe2CcqWszC10AQArxI3lHvYUSPJpLVSM+NZEwAsT4/o
X0syF8AE/2JDNRA7YwiebhOzRyMM3iOeGs4X1JV52/jRuwJ24DiGDQR66hFeRwVk
GN8ebI8KEwsj1AQhAkfc/bxm11T9LSho9Rpa2otyIP2NhrUQ0x7bD+FOOIb5w+e9
811UYT5JYYy0snnqCHSx+ZuIH54lfcoPV0ahrulsgZODZ2Dx5GIO+Bne4x4ajdvO
ueJwt/oh3yiyFM+DQFgASNjohFTFOVqE1FOkS86EsoGbno7O2X9uruFAx9rGcXH5
s1AFCrO982kiFrZpAaTAGyC+WtR6oq3LdOD2GpOQwxKu/f+TJz59IRk7re4BoMIg
jiGB1YmvqTDWarYRxxgF1X3HooqJu9zrLLHNe3fjxIzhYgC8dXNFGA+lZEyWPWzj
NzkiRdcAj90YNQGF1qQXm2QN9Q7F3ZHcWIgo+uYBuLNHKEweyBHlk3LVsDOlx0Db
IZnDBSk5ikGnZQrNGoFilyg8gUxewPbnGZJcVgaouJzWL1NOaTyjC4rvqdo/SmPi
8wztk4/hgAhkh81TUdlDaJenxgLgN28cyqPS91rbKhy1qP40jCAotIjv/QCGBPyI
BILKutReZgEJmL9MIPbeFHTS4V8/G3hArG6VJ0EkRoXs13rSedp/1HjQhnWfownC
iVwmU2u7xkm/WKewVnNPDR0rJIsoS783gw1sKQxmgbwcPGi5wYVD6jS+t+qwAFUx
4siAFm64hetrorKke+PHEhOx8rsbhFLp7kh66kVgafzxlrI2Q6yQRFTFfoFBaxbY
9eOvbFkNUUBebW/H7mN9p99nCIBNbXT5bN61Viqy2rjVkUZjoJhzMDc/xCzmrHH0
TdVNDJpa0LpM0kOVLgV7LBaVo6/lkNak1kbPO02U+xLCAX8D5LmHYx+Us+F3Eoew
alzOnqFYTWp6oJua3nTa0B/vKRzG8KjeUtyMTfp6X5G60CV9g4dinS259aRn4LgF
dudhFhETq6+ificCMnLyzzEw57Cb6HBTXMO0VaF6uJE6JQ6aD+aX4R2S/wDw9Ln+
OhHARWJRDTjAlCpS9Qqhtqt1JTIPJsuuVEdWcArjT3IHU99PpZjz1NfM05QqnDtq
h+pB6f/ogDARYjyZ5ZEJt4ese9zgxf8B4ikCqtXF6E0ZUZXFxsT6pNJOYvFpA2mK
jyR/vmuAq4K4KuFs5WF85fD2FZX9+WLye8GpI57/0Ml9Fmw++v8Cyudo/GlCCBlm
RTS2sRPPtAjhY2iycBjbpZeQ6GbxGCGC9XaGjAnkocrLaX/BO/YTRjjt5zxHAQrv
ctpfXsp0SuKOWnYDgeWeJCYeBDoW93XUDyisjq8uljG1kZ5oiGXPma9tw9sfaexf
Kr22O7HWCTxzzn7fPGGVMvFFkvnML8n4+ZaSVfGnt2AXqqQ4GdldTkFufxX0O5RJ
iXxDrndLFhuwucaSBxCuNE97S29e01DK+d+LQki7VFaJQkPF690odoNI0nv12j5W
mjb5ScvjUQfMQAmgTstbpuc3+Ev/S8lujoWdZ47CT34d6JnxObhEiJsSDQysHDse
a4QDGX+iDhe3qoRYF5Hh543NrrxVHre361abYHcG99vTR+Req6fx4xWJjInJ3FQG
YCswFjC+oZL1nnMcLYn4NcB27xJWT4/hx/yFfsFGdxNbXifQcUf7klNoxt81HmsQ
LAEO0zM+mbjKEGdpbgxye6Akmrb6QWPbIlrvs45viAMhh5d1GbpWBbe774QN4y3U
e9ErBTOCgcoYWV7XHDZJHk+PLxzlFi4e9tAcD/eACo7hcgUD/wIDNrH+viEShCEb
NtjIylpr3fdz173rlvPyl/ElyfUxDcV4xFJQ+BuUDIpe5W/0UmukKunyfTmGrq72
XgmLW4nycuzITxBF55VdnBENWax2V5J8Nvgk0kGE6bCICwxvXN1sA/Px6xcdo0cH
HV6tLnl65H0VhO8DOmJMOYTG/GpXt442hb3EcY+2otoZ6gSkQyjCB4V7a2ge66pY
hgkO6ElVR0nAI+hN9QzyXOq/jea1oyeV4ByeUgNTGSvPf4CNjWBe0amyGlulEwX5
c5Czyx9Bymaeyd+T8qS0dUmOwzUdjaNhlY9/SX0c7VCe0BKW8W6hkCKPz7seXcZI
WrgkV0Gs9Go0TuyEJ7wGq+zXNSO/SIcUSDX41wiMZ+thiKcBNi1VcXOJjW8mjgXb
X4EZFQ4uBIHupsM05d/Pzf2G2ow8FqK73PmhFV33MkcF+jN3LzY768KMthywog8k
exNOYtqGJrY93e7R00cI2m/SxnodLd7H5EzC6GlEDTIvXu2sT4xcZh206r2eS+lF
sHyuyMzduyQqk0mYl+tBueZsgdmaoLjy6UybFyV7Vbwlkulf2ejxiziYSFUmN5p3
c6spN5vK+l+DtDgInjcTF6y1Qs3EZw7rwD27MYO8C2yKp7s3w5NQJMtJT/I7MTR5
g+ffKW9lgr7/IKYxqsiQjcqXywsC8Kqcy8BUKOJp5NShCDdQuaZFjN+tMwcq+95a
Y1A7+/ne5H6BDwH81buOUfi+DW6KtSfyh6NUi/1q+vHM5pyYMdPD5oQJeidOc6OS
f/aByfDOqmscRnB5hoLvdvajySoyCfBtdZ0una/9EW1HGm+aC7YhObUjtUpu49mh
mabz7LB80mwNKDaSJzx2dul3l1jTprtWQHiCaLwF7sQIpsrGl5CG7eXtlZGjGs2p
BmyxyBgKveez7flXmQ3nWWMBxnT+EIe1NV3RSSyiLml/xZoyPFtB6P37fiVmtJNB
VFrWIqVpXcHEz1t/F8fGHy3KoxctZ1P31J6ZjQiOG2dz9WpWLCLZvC274s9rkqd5
Lwj3dNaz5hZBf1s2lCAs8tFfUbTIojVe99KNPuqtUUpo1SwhbOxQy/rufsWjhqya
/l3nRtoGr5u2+N1yNUUzhFE04YlQ4tT82zRi6TSzTbhLN+ZR1l0tkjznLXQZoeey
Uz/PmbPyj7RrToX0eQkzVHzlJnuB21FQmgTA6lH7SFdwSN8ojhb16etJcbAi3Dgt
W3dqtOVk0ZBSa1brmO41+m6MRUjV9f8o3OWEQMNu5x+eeQG5OwOOF3TBx11YHtmU
xYeCfXW5bk0PCP6gfjmKQnVoy2zODyzQjONXGMPZ+/n6w8P2LF3aWdXaPFAfvmft
ybOtKVI/EbAuRfrKSSGDvUJjxKrcZA0+xAs2aYz+tzsUVB+YDsiPoe2DKyZnLym2
wQpwHROrIuoD56NR5VArCiHsX1LfqJQc76uPAQEK/hnUZR1bARv0wDOBlhW1xBwF
A//rqfQ0xpibxqJeRAbXDkjhi8+0JlPtKNQV1rxZmBCplQijiFU+vIXsTw/Lq8Df
WrCsStfIG5Imu/gLCcVQdWnCfO+elKnon+d6ZfRcVaOhkdgfW2VicjSQa9MTAoiO
bRpk5XSU+GxywrtM/4jXg7vDv4hqvOXzqi9IbF3cxjUWQZ+cawTU/tl3fQX229yx
NHrJS5CJ7QC0ZpskUEIuUebq+CWrVRUZ0twLbRoELyzs1BmvNC+taI5nJraKN/wc
PR5SwYHEtqF0AU0Enxf5afiLNUqHS0Zrzyzcq9YkDu1KYl3WLBEwzZTKM7CRRztV
WNUIf4Ihi8SHgi5F9G+rBHCtH++OW7fcU09IgV8innt3cWJSv6QdEBD/yHFf11aF
blXqHh2D2Ng3Xm6qq4O3ivCnjM04U/gqPzNDOfALOS6u4bzYmsBYal4OKKDKB45g
dpyxcVVg/DpzpHatwACjELBrHIVZIZlquF5kVQXuC0cZ1Bmu8fK8+SB/ARUfGeqL
iresWr5bSTbAYHDD8zZk536R06bf75sF6BXJC5wg1AheIrgmNlvzy9eE69MZvSmS
JSPCldzGyaCmHrJisLRbkvR12w/kyhP8oTmc2+8V3TIm7UuHehoTPLFfJgvhi95J
cjVe6ZQ6Yj0LXc5um+gNAPU4hGValwv+c9ldj5UPGXzuTW7RuoFgkVOQ/+1bqJzy
S3AMkdHfV7rLbxlagZC4TZa4w+jWPj7Stvz7s10AVz/d6amx2hq7BvmeA3hU88B3
kWo64JaNNxsOJ1+PX04NIKAvlT8asGy+47KtL+IEcLL5RW6/UdPn3B1JxW4bnjBO
FIo64RU3R5QIeJie9+A5IlSZiHOpoYOR9Zab0jyBENMhJ3NmybUKC21Txfp5lMJ1
bI6+TO2RzpsHmjCcxOo01LppeYO5zRk7p5n3l2CF0ppK0F6cPNGOFJZ3PQtsLTDE
uT6K7XyF+mqVXon2QPCAC4U+G4pI4K9pBTynvOrHyE7XqHsqYmqurdUGiYuBCcqW
ay73Qu0y0EEBnXci/JDoZ8ExVBRSKuQIp0vslfM60ZUCw+zLpT7yAlQ8Tovvz1Fg
ABIz9EFCuuuPptNSBJGKz+vK86Kfn5o0Yo91vVk9kTKmsWx81aT46R2e8Ti3+uXd
0V8RJOfXoIHaQ9N0VtESq/cAjkytjC/gb1KlPC5PxfKz+X4kKXpsJtFXneZyXyQs
6MtSbGfcwkT8R5jw/mo0MJPAPghhUpCqYrmf26P+CkSfXUvwCB36zPwDIzOqhfA3
MmuCA+fAb1gceOH+ZMf1HbqcUH3ny4oGB2ouu+kZK7ZfDALURUqNzCRjWSV6lEW2
UpvEiUmdyprQtuVuWa1lOI+0VwM4ILUsRAXazWzyI07PiJ++K75QYpZ9R37jFSh+
/k0TyEEfDblCvCS4Ly88LbwfIohQgRqb3KOmLXb6OFdwjM/PYFy0YF1E/YUdEfuI
8Zi9yrrpwz4X7jmJeyhBjGBJDVVvrnbCPD2yyS07liFw3g85ihs/mgv7f2xPjQTJ
DkauRiwVAN3AVBq7UtNuuXpaBW9HtkX77cY5HMMVTx8tmMtCsyCSGuV+hrGzytOz
3/L2mWLRn+OvKP4id1u7eGii/nadFQB8PPTH9yiuwsh46aEPnIJEeW81F++xkioK
GeaALTZaXWkmDXhp/khTaClv8wLAeXHq+s7ekiVjeGYNN1C3b3W98qG2B2HzzuMz
zliQnXWvNgPy4JoiJwhFKGbwRbXrcVYoAjnhrrCfE1LX4FzV+f+Jk0Daos7bo3Mu
d6u5lQmT2s5G0zpXXHa/FSd4ufPdtXbj5HDJlG9sK238lXfro0fK2o7DSMDG2qOp
dnztkyV9XJbMhsXIaWHBlNfw3XQNxYC5AKt7RluxGkrecneA0tU0SRi73uK2KiRk
axYgXgL4Lum275OzNehRhkzOZoFq3DKZwGjkkfvkGHuDAsJO8yXUtCACrYGZ8JAZ
6d8Ek4WkXuWNH3gP5l6BGE4UAtBwAI4BVz3Cos4STdQm29PxxV5FwZlrGUTMZ/9L
ytLyuRWIatdijojC5ymvrOuaqAiXH3cKnvQ4FeQt9NPfo/9d9Wcoo+v7NcobqLJZ
ltEyAfGXI3rfqccRP0JSQyj1g8zRPk0rTr6CI77/3n2iAMe5Qes3LtJ59AFur96z
FnzvaOd+nOaOUrl81ll9uCqRsPt/rMCuyWv7/KOTzW6++Dc5+AbWWFhtcxQ9ROUC
W6H7Ufpub7ZlRxycEKn0zjgIva60Dss8pnvshWMrimQGDFeCRPHuo+aMwjYfFkCg
PU5P9b9lfGiDMpo0a21so1aVQ9XSTZgF2/em8UqjHsE4P8N77ZfjOeIHPsh4zAzN
FXxDyjedy0AwnJTwTiMkMOZEfHYWU7Ke/O/bmu98WL9t23yurEWkhcJu+kwpGoGx
/eqA1xSmFEnDequjUd7EkF9Me7Bm+loyyMdgBHLyIWbMdWy3DL+RKdEWW45+g6O0
d5QlwX7tmvp5JHUL74XIUSswaL6gWeNIdAJnnTjVDwjVqcV0gCkE78Z0ZtJUtRgW
w/cLjSG/3B+MNXc39d8E+PRYP9ptizeC1vJfhGbFew9EorKyzRajKgAuZUb+aU6k
EGWXluX92SXl0fB4m8OR+yHQe6dC09M1coUFdYFeKNXQzxFd1p9rT3+I9CiQWKk2
Dg8vQichaNUtLJM0Ld5lrUgOLNi7qNAtdP1uZSroV41goRyIcWtA6odcmj1/WH+6
Gy96jnJooERUcJ9qE13rne4uWK8/GM9hLIBbmo76VYzHQLPbVaXgvXmVzjBGxpLn
eaztyzQs70qauPkWwJ7MZH+suZlo8EO0knhsxRvHQZCQIf6GIS9d5w6B1+7dDqfR
oq0pg01OzL05EWnPqPRqVsVN2dzgA/EHXkod1g5zgu6YpHaMhz0HpPFSUXfH/fc5
/LN0ZQTXOzvGdp1koS2wExeuZMH074pFK43XssYTLiARU2EUN52CO647yanvwRyv
i/FPPoCIq2kfWbGyZiVeoubx8cQpIZw6voF49eP+xrpqMvXAG5lj9w0qXKgcvg+2
udZHu7wrkINxrFMlwxmJWqPwN6MNQKGZvMWqhQ+u3BPsfIYlOmhl+wD2yPapYoxl
dDn5lXjG35nHp2mSpqzUp1dhlkFl6DQ7lFE0FDHZSB93I4wpAdTqVRnvJWSdsYVj
UQWk/AG3sKtKm38XVAm2Fw6ortbFTO4jDoTHq4/j+QKfiE0+5xPBefBeSRjeCe4d
9Nnft9at4y4zyeNQnIFrjRsq8Q6gbMcLBo5px0FjV32fb7GsiH6M8RCTw0kjxuf8
Z8DGaZVYlNTVuAjvxdamVL4SN+cNcAkDNHEzvvoiv9mkxmhMUPXPyFslWJsRRfJY
svzd2+c/VKdDgF+FUQJu6m0rt5d8xXBOn34WX1dhfu9pq9BKtYlK+ezxsLWOJ2Wo
XSUEs3L8p4rXvQJYn2nGyHrAFLu4lD/hVzrWgHhT25252ZBIcYVDHHZuIZ1w6o+o
D+YjrW4jwZX0L+bgx+Dvxl/dDffkIRo6RzapP5prvT4zIL/DTcCqQMP+uX1nlhOA
NUt0LauYLSLC/kPYAZjBhtUOYV/oVjPglV3Fn/3XOyBdTG24DZKUlBV7Fb36Gxca
H4meNTVMo6Ab41S8HepMe3hvbnb9YTAfp+VFyXHgPlDB+QMY0j6qOwoqgbOZODJj
IUoQvfURqojk+yRShpwXAiHusCLOx7OgYrZYEYOFjs3Svr7Mur5jwpr3qhj9PnVg
VJ5ubsxWMJzmlvn1yfhCz9NJHT4oITU7hf2zGpA5hgmteMvz+wUh2/hI0gsFV5Ee
RuEP5WjmS1P6zKTupRn1R48C6tMNU1XBj5vr+AtBQ8RbmF4cWEdFf7AuvWbu28Wp
O9MYRW3QKShF38tAmX75jk87xBj7igxw92aumiSsxMI/O3hLN10cRNBZ2SHFF6Li
QpFR/NC3ixECBmHsUtgjsjJIv6b66TvKNfah0+hTtJKgIBnCBBTmLg2HWKtS1JdP
6EEeGRNE2wZ/yQC/0Xz0p4PqkluQGA1jzp6dCeH70kM6mLTe6zp561LJuFiyddl9
AcbXrYrjEHIowd26Jj/WRIoXsdGeTvcRBjjSdg9+3WTKNlIae8XX3Nyszh2TUhDT
XMnAmUuEGZqHmZ9peYMzp5sobbpYixjy9GVkQCYh3v1st7D7wxBAc2JqBqFBKiHN
GJ8CHcaEVgwNDaapxlPFLor+dZR2rb6xvvuZdvXvJ8WN3OZSI9+RDex90twO99nP
J9gvmEPIuocmCj1wSUgtIHtQKKCAc76+MJteklx/iOtrmI+UgUGLUoA8926oKpGs
+TwluXVsUWJMpQCGq6PekTaEMd5ab10TOnHoCdJOapJ4ev00HK+9KXPLGHFCYdo/
jjzb3W3N3kvswxNkALaZlRjYD7TBoVDZDTrZHujduVbKXecMQQw7TMOw8le25B0K
5h/RYTroTQIBt83v8/8+SOAOpv0thFYSOInwH/U6NFdGyo2zrwcOZ9d8v5mptoGG
yCeXtyM9awCs3GdN3PH1j1yU2vuGQqHWzFDtRBIthzlIarvYRohuI7GvJW++cOBD
mJilaDpTcm+nbqKxBbvqewGf9L6GF98L+V5Y9rgbSwUX7zIZ5HKJqtpc2/U5uELn
5ZHWrURyTcFad2dyovQ5XJku82bsgsRLgKB1FF/gV+VBO0Kgst0uoOsqijmXZBR4
7WNaDUwnv6+cNODDoaVmL5CDDQqAejpl2q5lFD9HLCcEovAFJ9Vz2k9uTuFpY21M
g0KkK7PwzL7zRite2xU/gR5wBQB3Ay1X9y+ptsTztGRiZqtbnFVroyL8vV2jQc73
Cg9AEox1o4id0Fi3ulvoiDwo4oscTMkSeCV8GhR2B4rRwQweOEMBacCn4/HaVfwu
VrCo0aL8EQxtrChH+lR1h6rK5e+6CnXny9ENfnzopv5yWZtcAIlsFBg/E9s946tj
lkpKAO3aGdnCHEfNn6IaCYZNd5u3KPBrLouD4DaLHBF++a7qNG/nMOuSBnXjKcNQ
zJ9UFUzf9O8lsNkQ3bhRElqPkrt2OkhX7a1JCHNvgHkrXhXe7yjXOIKq+WhuFNjn
yxNb30wlz2V5df3VCIp77jADxAmrrKIvBXWXsXk51gktZ778NMrXh0RYpglpmww0
bmfGPyX5ETRIbogwAzJJGmGIaIGAiDpSuMAMYpoYvWS8WssrTk5mTXndjVi6qOit
8WZV6EudiFhR5ttu7f4EW2PAw7YXUQAh6II6Wt5KOHupksMWicLJ2K8heKok+3u4
zsigOJ6k190+9PLAzSmlKtoMgAzKSpfcGYUcdssZ6x1HCn40+hIAC+Jzp0Txqnj0
qkqN/PG0PCjGq2JZxUMazCTnvvViz/bT6/gzuzgJVr1ZljFTpvnVNFJw8URjADuI
BzBYtXlYLtm6dizNsiEzWYCOYBvkwF5a1lh02sye5HiKBOR2Qw62weT8TpGEZwEq
O3xdXSt6LMz4eFnfhnWhfDtOTcg90Gg0Y70QRfdSnU6eG33wZ8SMNNA2uCpvEzKN
KvdMY7Ki5VGz+tE68eca+J6RyRuEknlVM6TSltBoYFRXAzTlTfpCaGHE05dlyZkD
BbdqDgt2yLRkAdDyxyta6rUnKYzLR+eYNky+X49yoB9OwcrdpkYECfJcIblWxhRj
AH4++zRiI+Jqhz2YGe4w2exFEoUabdV9mkBGtYDH0dGWOssOFo/1l8RQfBVZz6fY
yXHOtw6Cx+1Sxh+FBimqx04TesTVZjyctGnWPt8RwARGpDoPsQmlRBJ32D4Gobg+
uPpWZWo01q9QQsp9evmwh3AVJk+KHMv6++63FGDWe5qndkE0NaqfOSP2xC9yepD+
MM6PXIISkOQ4vhu7mpc15BTiFag5quFppqYNnNVG8GJWLkg6k/1vrbd+9Ma/1xGb
f5bu9iHGNbB+Gw5NvTsCgZvn189hAv3IQzJAiH7bxMfg+qIQqpp2vpRfj07eNi5o
aolN+vJNszNvRKZPcCP9unjiOnzZNmWOGfAPXhYYKq5zFtBKZwHpVz+ne7Mtf055
HlSm0gaEa7EchSac5cS09HbgrXMV/M0fwiLYho4w25Hs1PN1Knti0osZ+n/q3o8l
JRntu08yLyKGOGQIAqzcFR/Cs5V4n6bmRNJ3bq6xab9ouNZ4d0x2kV5ls33N07WM
s2oq0k8hsiVZkc8rVcE6gtJEv/RS7cSHbDGIj7GXtIIojZWram5RLr8d4sNsGmbW
bJt7G3HMXj03TiLr8sHLaiAKPQOwl/4Lu0y9U1nG6HW47Gws1aeNbSpaDKcW/9zp
F1I07PaLfAC9uz1WvMW3rINPyh+6kAoKlGAO+s4w9VBIvWMh60kpIzd0CEnEIui5
JEtN9iW6c31lMbJGTgkX2zkiJ8VWYNsuPnbwcxnVFke1mZ9UkZQeaf9eO99ZKjZG
nG7AJP3OUGQk5k6PpE6GVpf+RsJzZtmii7CkIApucVxYsgHjmt6z2z4UZhpTjGUu
NQ50u70W+cZOuUtUp1gXQdS7YkSsekcFOw55kkkRo6KofkE+Go8FQzKpQkY3ZWFb
xg4Cn/MQzFCi6iUctKV9zs++3LnmpvQsJPkLv+vkGcP4uVTo+/wSe1nY9imqTOYe
RTC6MF0QKzEVT7Ip1zLqtFu4I+3gLlVXEul9lPg2CiYa1KR2SbNytPl7EhCfaTbx
O9b/DyxS5yE2GCSgmzs+mFILXt5tDzxbMOt+xMJyg11yjkpT3Xpuo/ioC9ORzKMh
4Efc2FXDjF5hJEWuA1kd4mJUnvbmfiW06B7amS1qpAKdIL+g8+56xfpyEqyQ0gEf
iUL6NQUapimarli8W80p7DOsLvYbNdqjCJjOLusPb1sEtS6RuQGcqIFHwc58bRGw
yGE6+kbSI5ZDDY2R8G6svsY4HCNF+kcxklXgjikyrf2eW0y3o8qraJ4E+K/ZfWBE
z1A8K8W+Td8jABqiJOM6axptODEOhrYyKeegJW3yW4YdOyDCXtdIsh6XfTB1AjVG
3gret+DIa+hUFjlgLAFUj7Iin9A8c/8xB7J8/21zBwyc6BHz5/mOH2aLFxycsCoz
9hQuqxzEwnYfvy4XVccffstYG4Nq7mVcgRSksrWsR+zSkXa04NOWlS9pw95VO/Iv
ANhyqLgTmDCimiqr+I59ijLVgnH1qbQOjY2kTkA/Zbk6T1RCyrKO4clhsknlCm8f
KECi3955sHV9BRiD1pSDuHSEhEyys5z98zNSh8QtsMeoIRK7Tqav+YVnQFNmvSiP
YIuxAWlT5F1aem30M043rmcCOJcffh9U+dAPPV4dnOpq+j0AGEUE9Ej94yPS4lG4
r41U6M569/bHBIdVd2pYPoEQg1Y3HA7ltQepo/Giycv5DRU3dPU2QehmzmPbOn43
eIUf15U/2DxEWrlQnTYSKlXUlMmGACBePebTvIQNEIEl6NPjYHT3idPqHrIEpTuR
VMTf4JoE07/T3NWPOo+9me8xuYHsG24B5OhIKZKzQA06FFKl678hzcxBIzIYt2Tw
GL+i2zyisw9VoOlmGDuvWLb+MuEv6hySbtRftkTgh2USgEBQ4diSrF+lzatz+daM
5WAUfbIwFUj7alKl349HDrYIon6UJAKYfvJsoOFH/a4KPZJK3KZHrocUtzMieoNc
vKIEjnyDgUIB5BAE7UZzpCx6QkHrgakp+hFIXKR21GaINQgAODRg3bcl3B9Z/2QF
YdUBgwQ7xt27p/QYjcMsekWRqO23/m6uK0eQl7eKqsxrugkFjz3pXDfyKcTsehQr
ifir7PqjXybMToyoIqspP9+Mdf3p/Iw18zn/UZCSDzPeH3lhQdnSgbWaGiz8HlA6
OAVSey6gNAjESi2R1z9/Qw6KN3RWcRUEQN2rzZy3/WNRCLxtpoER8LjNHSV1ZcfY
q8j+hvoIfhR/WLpseTEZGY/RtCIZUYov7agOaZRzP6dvQcx86VFYOwYKsZd3LElF
tU0gFNAWWxCOOD9gHBnBGxz3er+1qkG20nlHFeLgyK3OEuPizH/QmtORKgqOv36n
pyrH+7LVbACoY9SkHm+x1trSF47fZxkPTbEyX9IRDyqFj0xZ0avq53ZcLiW2OZse
CmubK7Tv00aeBxGQjEAJ2iB2VmJyGYV8RVij1fPKAXE4/1F8ffY4zw7mUTUep+6I
0q2jNfEHRSkmfRCPnqsXKjmXbXtBqjusQGW3mEojZFH5kaRhhFW6SXMi9q/yBG4X
qiz7DbFQn41TSUiJHqbPBJKM0FNirp5VNVPz01xd8PBAurx3ln8CqzbybF3XWlkl
ZVb34KGKlhWF7QsOZsWl1Xb/gwbvRaY0xP0qZNkzsXszd0ehqVqFZBqzK+yo9/qn
/OeaAcQWG6K4ynGo1qMiB6URKX8R3PtxztPzuaIIAiZTgx9VoTNXhBS+76BK2/Nu
DVTYjMLAZ7nnuWITi8KYUVTx0WwZKwCS32jJA8Ka4F/M1F6w4pTt7wuSZ5W/Blt7
HQ8crGUZ2wJaNm6q5UBXCsMsYDeR+tu8Vj2sJ3oXSO54otBMI+9F49Zu4nOxHFLc
vQm+tP23KztD9fmueLGGWB/bG2LahtTd5xAqt7+9UsWfqSm6HogI9NeZ2Z9sLiuc
JbDRvipObXpsxqQWpZ9LRBaLQJhzxNSJVo/ya63xXoUHNYn+jUrJcRIjcuboYJMJ
eGQbkXj7UC3Axx+MzJUXAL+RwbZctzcSj+Dh/utdM3S3mraAs0Vnl2U8Z6vzYHfW
hplabLFF8usd7Meks5GFOM8ZHtHG5Ol8XtfMEURn17OA4MsZP5IHSBHcqaiwIsov
jDNdA7r4+TiDKo4JPe/jUP8ZtV4ote8E4r7ZARV/ZsSkq2ktPaZqYp54X7tSO9Qn
75m1hiBVtIjicQ5+dUIEe3nYJrBfmzEYnPSkLv8fsPRLkPlw4BW+rG5xQye4+VTj
5xvPte1vBASlwVGKsqZ/2rO1d9dDQsLnGR3EJsebZ3ZvTe1YJRMbGqn7wuTP82As
IfYPWP7fPdy6YszJKGq7BRxWaO3/urk703bm8YoaVbo4zNyBweGG11oZnGYh+wKb
8SdnzUIX0NwNddPYTpwMgpGJfj+kbnqI3OVm5W7rx7NsUXZYmTaIAq//zkw5VP/j
R3nO7hbOt5b33WXNTdFKo00IyFW0dcJB1jwUrIIQ5lsc42Oz3UGwKsdQ8/JGT9fP
HQiIu760Y9q75W4ZTB5FYVkp2oOR6XUAlt0JP5hXA34VR28LBmhK8hN+BJpJBX2T
hTDU/Ll67PUD5b3fqYR64LCf6AqhPqWC6kQ3MWWkEA4DRgwinbcQSu7CBg1uJ9H3
6AxSvLaQ3IBkeP8WomOynimoCj9Cw7z7TVO5SQR7jsfJAWTUHpZ9Nrti0Iv1Ronk
kd8Lsg2ADWHoE0W/+tE864A2dQUornyuXQ+lKFWiqX0aBhMKfYYj8R9i3WfQOnbU
zVgJSrXGuxTvMsqpmvyx7d/pFKajytYiahV3/PWdNdAcQY753SaxzpE7ugRpq5gb
3fycmpBqbVYFgC0bpcLmheha9JXskID9+PJ4SLLaS0gQmE79dOhamKmdqjxpyDZa
kWOyIllbXoAc6zL2rsLjxVOgvDlnNe792yQD0dOIpb26w2T2BTChkOAg1caj3ITl
AT5bWE0vh/FOTmXsB+iYC2lGzZC9pojjm2+GVXwlQRzIahwb9XdRNJv8RhLnEhjp
x4YkkihtOvcw1ti28MZOOJPEwAFFToqgyiDp24YBoA2hfHoclliZFSLZThzVJ3Lo
KIKIKGKPwqauur/o1gYlEV3n65irh4mtH/wiIQnhnVKeYJe4F0KU8KC7+CTcwi+s
/GvilULEXwpq88rFksO7YFtPnRwMYjT3Vh/Zg9/AGjCW/roxUQUM+vYiLhjI9vw6
a7SpBmQApqdVnv8Vy6KTO0LFg5yfqm30G20PqYF3ckL6y+2SJ9YWAl6iwaPepATU
EsozURdZowRVkfUzlO+0KYYGxbM5z4xVPiBK5MQzjC4Ysbqb23lqgC1M5B7WE7HB
N7T3Xm0xchGM/EKS1ilMTP1P+RrFJFjWMKl2H6MZstOfPsXjLtmQZ0ebOsUNqYmK
hnR4DsMfXWMFUB4KPdSZn5O2wPke+O+mZhn5Zs9y+sKlRHNw9t+/mVnwqA1qSbq9
KstKFPGAlz2CGco/i+6waUy8zFCyejagKeq4AGSI2Oh+u/+mdNB+Bsk5SEDZZcLA
4FT3t5DLoUZB7rFT/6J+F+xRTT+GRVvTCXPMLgaumIZoO7V51VUU1TXxF2I6x/U5
sIuILUOIWMJS3dPv1l/U/n7g8DM81zjAX+47saVvJTlcLXDVS0YL0ni67+W/2/DC
pfJsTykmNcUrN2BfM/JGh+Prw4AY4iibAbqASTMw6cmygHxf0cwTul6DaXy0D9Zv
Z5zLHNDYy9cEaQjTUX7sfJVQgYGzRAnKG3CtMhBupil6O43nggVxJ5KFiUNjO925
aABRPodF+ACeVmrwLOCCw7x07wNGQ6Dqirg5TYd/aDG1cx1LosJ+bhbw2qdx7bq6
M1UWs6dPxSYKed+by+fJxkwQGJ3S7lJE1OhnYGuqrpl/N0//aBDb1zgKehI6mOeU
aAnooyKPQSuZpGcEcLWGJ5GJbKqShG+1CrkZELeaKHc2TtOCzvcS/hTBkMOzD0ND
qaQ2sfKDHZ0zTMQANa41JFTVYccRjrdF5Xn7I5GYq6Syecft+dmKDAD2vQHJl8Re
H13NunPXZWdDk95hisbhFBhQ0fKQxi2tJbp7tWY8MOacofmzlUlaZojTmz9riQqV
EENqBSgfYlVGlgQFfcCQHNQqBxdnnxnKs28yrHr13c4tIS5L4t2S9SqbXkEM6lEs
cW9AkETaDVQFWXIVlTtRvpoITfeseNeYTxpCy0FOFiqBmNV9hagO3/CoeMR/a35a
Yx++0bVFzbNpzaQUqHvuCoP5D7KMdEpcr5sqtUIOwvF89x52ovTWbLGhvL/j4fEC
M1/WfEo+E1mfzF9B0lMC0xjT3sxukLUjyOKaeKfjkBJblin1wom1+tCzOb5GM2vl
gYxmZErN+HFa4fpjl+vN8KKgnVmCK/jOlsH7rkrxGdcaaXghoTBjcMHt0L/lvuPF
kGgwZd0i3HPJtRJwEdrWYHXETgIMKkK7T8nMFvThWdI3qaN5EXar3T4R/RyhZFZV
hZp0pGmhukbBKSCFq57bhwGjOGuUhWu9tl/IVVo5YPIdt5sZraapZmAZZsyprCEy
s27Ehfj8jtUKgknAgLEdJlilFX185E4fWDtytRP+I05P7/aJtX0L1BRdZh4/vZq9
595x1pZqtJgTyrpFzdCG/0qEWGIjz1tV9pj7dj4RUuwLJkXEm8XDOc3HMBxl/k3U
JrApGAK6M+VPraF2dsZ7zMOqQjQYRo44qwuB1KEkb1lBYWZvH8UDYqfJHw4RXpKR
io0468pXTXf+Nixo2Q+7jitAuL4ouC8jtEJqoUBgVrE6QL410m/zKAreGqHCtEVo
PvRjBAH1XzuLJFfvR850zZEnM/JaYinGji400ztZW5g3I7gGGU3A1GOj+pdYiEJB
1qpTny71qy9cTezo8hw8FN3enOhljP2khZmWdHA1HyKyjJFSI8qovZSZ2fji+Zmj
xqqxk+xT9LIomTiCaloOSE45D3Gh8+T6G3g5uWfutIqnv2/1/zj2yG/GQsFS8qsf
5jtBDVU2sDXUxMF/wioZ0UXPWJ6yKkzfhLQvdThufuuNkmfIBeCjaDEqvwyiqsEy
SBk/3FqkEHlGFdof0HfYY7bGeySp3msxIF5GFWZh5TSx76bKrbuo4N8xcN+gQ4eV
JJlnYBeO/+/CRyZlFnjsJZYMw94pW5fS5BHcqkJ04y3sTbMyMJbQ2muttOY4RAUU
FilIGFWYpAfTuctpjZGi06wSKnfynsQQscIOG6uTst2pDlLHvHw7gwVrHCDFR6U3
MIJy6zGQQWaQPzFpZQ5I7IxpS94XHNhCJPwIUsqwfaLeuxsCaTgwDI0DJQFN3o3s
AkfXr5QmYVsTq7HPNzPyksFB9lVDpxsXTMIGrbtTilP75dti4ruOSKf5LHeCnK68
hT2rNrUawUVN1ZpmwdKlRZkNrIKi1eXCReo14b5YY6wLhSiRzOwR9GgN9nJuF84h
HdLPfYB2yPFMPU6eiM7U18VSkWhdp5GReUBsB02YuqdD09auvzaOeJaxkrB9NnCU
ccTyHRKr/oDY6R2X+DRBFU1ZO8ejf2CDi30ZHBYiB6JkaNTdEb9tfLKwuLSMBR2Z
RCPB+dLQJwkn5G7bmOZ4CBGCWSgm22Gmo2Xh8h9XC8jNNUFJFp9eRJg2SB6C6W7w
n3s/ZcVbs6C+SfKW+lr5rX2CwyWkJZWEY8RZVwtmnzEEsPdOpjGjI46p+rbfVGwr
rdY3z8GLjTfoqgNRIFQrljb72LsETay7ofkzFem15Rnc6dxOBV9D7rlYl61qUebQ
4buxyIiMsluCRHSdsKLpcGJsbXJF0IjudQ2D1HxdKlLiC+XNSIbFQ5/Wdm2uFOBD
9InV7K3hlg8COxb0m2XdAI39MrOXbDM4pubnDg4T/8JThEz2MP4OMx1Ta+QtTyKf
KAIEXqYKIVO/3GMIXiFfH8jfNmFm4eSyP5wrVPlth07pwKpyBWwCYCmM9h3B0BFX
ShrdwEGg52g4jy832T5I47KPlAeWCIxn5Zqrj3Up9QDE3bQzwsibS3VS1m6lirwy
0R0mrH8jztmj1VxZUAUmcsucn53TIsq42trPvBwSglz5O0tKLvnC05WoUCjbVoEU
kgTdmlJAET5sFI+Iv9psPrX/LRgtchtgaI9wtmgz5CK51IbXxNIs2BdmtGNndkEd
eM0nTKJl6LlzgEz82Q5100xtOalxKNGfXAKDCwCvGG/pzBZDJdoPFlY8wLXHMaJY
/pfU4LgdMzscYgvVGmM2/yaJAGuVinHIm9xipHFyYezlo1oMVetFyQJszuXUzqwU
OD2Y+5cit+iOtluLdWbg7tr0aSXqJILzUEt1WdmVqCdzi5QPWY3WNXQSQusCF0qK
cG9b9FlIxp8PCHGSSS2GTwnHdqTtRjIF5DKqcoq8icC0/moneMTO6lpcL/vF3+ru
oEVCXaOqvpGHGlS5V4SVDbeHiEdpCSNdXO3h2W4WrUFBm3mN51eeFGxCpME3lxW0
WlvBd1i8fzNox2fza5KtjjA5mrMaAY+e9t4HJL5ohPxUEC3/Bxm2+75eOtlsi1Wz
Jvlt/3NbwPwjULGexT/kyh2i4JH7T3qkrO67T8ha0RhOU1+AoBVXIsc1J91TkYLt
rq5jzGSOW3WC7VXDus8DVKU3ntVxJCJHz1opuluDFl6DtIMd55nP7HukzU2hutHX
hm1ZGomqggA8qkJ5VbQr/hq7m3tY7Df1UT2b+gSxgRALlKpBs9pGjKmRhdbGL+Tw
A6rz8L0T0692VA0pVp/ifE4jsV1HM+Cre7N3cztQPSIVbY371xumG2P6AXRy2WGD
KTXuATBC5IB5/poO/o2g5moCdKr4ZS23alR7pAA3BKPeeGCI2rIBYLCQDXErOU1M
3Anh6nBcGASZgjcOpw30hJmAvriO2rU5DZo1OBo4n7PYxbthOjpFJ+akeUl+/k/K
Mt87lBxDaFXYU1w+jTTp9zbRYchbSfLTMQzDbRaXSPOchY+ssrGjp0gpNeO1YXYv
zcPKThEDoivnnahbmR1d5P3t9pYctWL7tL8u2ZssadH6llYVyxlfkNZtwrzaNZKr
anC3Y+Sm/dKewqTyaNIeR8VJCbZGh4fyIQPJ+UB550VfzLWJhEp9JIa874xcw6ZP
xMKx8Vz7DTYJbo2Z4iMBtnqoNuz4RPqiSSLN8QMvWeHWJ3PfF/rNWjnHhda9nA9n
ASeWE/qKj/Ec0LLx70CHGGuzmq6+PeHV6D5UbLl84qjB+2timBEan5eDDEXWRbQF
mOSuSFhebm0lgRrlVpvqzkig7K3vbAfXzCo4egdE5XgpGkHbzio3ItVJ6RAQXBva
Ja9I8QCYRAlTkM9YNmDUlDcZfEDWFooXyJPIQZQkFaZmw5eN9WK4p802PuetHgBS
x2/D3Yl1VGpo35OdnSQlyUWHkLgi/tccMpY7yIoyevGR+Sww0/f9rFNyrsWbiPSJ
BXrrA0mEQTZGUfb5eW7rS8BBIer9hHhx0Umx5per2V/WYbeK8Gyevx64z5aF/z3W
1esWicJxsxpmxuPq9kdjv6fHRlZ1jnKmLZQAafVWAV88vu5njDVnpGCSQ2Ti0yVh
8SN0lneuBGZ4DutZBxvEMvH8X8hJZB/z1dcmh9a/6dIbYjMBrkc+9cMe6forJtLh
97P1w295/XIGvPUUuxRLNrpg9Uz5tDYZVMsBElSAqMb+0e3PpBMBhlV5n6Dys+q/
QCIZgmFOKNB+wuXpK/vVCnfhquGfBqGQIvO24zl+BRAXctNXlpvMlsmz7qLD6mn1
EMry6aJIgU0qgh54ZWMxtnAQrmDst0yJqEwISE9Iyfz2qFOZ2ptwVNp1LYIZV4eR
2te86aPY0tvmvmsB6g13KxL/FTNYT/R3kRLOIMy7qCXMxNG+gY9HTbTLrqt8llb1
ddwMsthwwAkOVadBubGKEerM/Rd6NQXCE79n0zf+fZvBAeNOX5Jf2dNqg3k+cphR
eRvsKHQrnYk0p/1/nkUroTdsaglm+2vn4M2/SSylX/ICRiWMrrXMyI1Wt6LY34LR
8C7aqI2mTep7Jk7R6f9ZlRi1OjrIFX9IUdMKhyneF33IkszZcM2tCwHfgasBg8IW
psim3KI+RCjFr6VWofwA5C//QFucCRi5WDs9J+YsV6pzA/tSk7CJ/h0U9cP5K43/
AhDFwcik/2LacFxepMyEEnVksV7uAW1Km/wAOSgGacv0z7VxsRd84JW4O2H+7BEZ
Kj5MaC0mVtpEu6djkTxb6vWzud2ZOlak0joTV8XnlOlXvoQ75Y7M77JTVTFDmIB/
RnSXhgux2RwzmyxkVEG6cGDSYfMmhrIsYCs1NZzq4WQiNA7Xajt6uaOBtAx8Muy+
y5H7tdnf3TLxSBylUFAmtMNblsepnEa5BzvU5dcyd8YqfO/hPHSe8Uf8pXqW1OB7
8V5U+S9DrFQxvXTuAIdrqATg9fiK3lgOc/Wi8IZdp+g7rp4AnwRfLfK94hjn6z06
WTeOgvv4o4JNG7Spqw2Xdh3g3jypCUAxRzymLn2o6cRLjyl3k/8Pn8+r3uVbdbfv
teY7wqPc/CTYXSuuUHinH3jGx8+tKJw42TiAd7/f3dzkFGJE6q9l/mgxpBfyGWd+
sdxbWKNME+DThnB9nVQFptoDiNqMXyNEPJ4lhsGBIiaqxZSOeKArgQm1DXh9lpy+
65gV3F6vcAiKm35J7Wv5Gag8+xuoqSLj1eZgAix1oeFQaBiu0G1ddIjQfgLmeEv2
PKjm4qRttoCj6YmS6/gsn6y+JHTqfr5tf2hfMdmM805P5xwCtob6PQVSTbIfkQRT
0H9tXIvrkbOJJ8ht8PIX8RkEAD2qrWu/gsV67Jteg/7Z85wxvkOOV/QBkTOCoY2B
MVKctf5NVnMnkOO6vICVYPjZ0v5Rz+hTacCkEvpsMBZ0a7eqFNxWe4ZBg5zXoYwv
GRsgS/SKbp2U4a4RIJE5vCkqJnrB8WxGIQqJzbs2cqWG5FZiTUcT4z84zwLbXTUt
ZDHMfiT/DoafOMyXy9pwm4bovK6UB2RCQNv+AXPuAl6SKtKVkWBExcb3tC32bWLO
A5Auf7X4BFSC7oZGV5ysn/tjjAnge/76Wb9p7A9ejSYgA9TVFOq93z+ud3WDjEPp
odH+9IOv6JqsE4YWo0bryvQoMqLogY1Cm/znftIV8cZKEc+b8WtpKOJCO/Q0/KmI
sgdXYD15QgOauqJOldTz3AtQdVQfHOP+9QgfSXQjKRKCrOcy9q2yQzSKmhAMWqQk
7Hax3t0z+kVoFZNZNOrWObc64YH3mKXPL47ftOqYJEaAighMzxZP5VFG/qGErZS7
5ZMQO+/P6SdHOlPMU+xy6U/uMxf9U0/eKn5EaNQUdVSBCtXuo6g3XlKPWYRf0jqT
ma7nOY0xUiB48M/xWbfkQ2faeggPV5jUf/buhmxIvR7RgyAnOlEg0PjPwBEemRIJ
5P15jneIUBh1TGj7ot0meYOe+Yq1urJoIejYmYsvljpX4j4Vo/zXyHaGDx1ouozj
rDnlqiiKpzLhUrxneH3Wz9q7LphuywJURW/zlu9fjEAnkUofRfOrzdeRyU5Sa3ne
BAIfIFtt4UKLJk+w6K2UZJIPoqhYD++RknIgZ2Iy87CdLVpCzEt1vOn05TI8/RYC
qaIxOoRrf6OfnFZ9dzUD0wUcYc2jiG46hiun+l37GQojXq2mh/ppFf3JUfhQcZZz
cJIT82BiIjw1TD06DCEXYxpECM23g2DFy7nVwMXFoPegtoRu8thgZfalIHjYTDHZ
mtOF4L3Q1YR4nB/7tkNWffaeFtnLGTcxDrN2jKl3zPselkN7VXaN7+b0rom6vkMu
rWa/N9+tuAP+Phs5ImHolU3uNwNpQP27B6015DWbZaGhIjJlYpEU5rpZX4ZzRnG3
CJLCLk5OHPzzMc5sEPzNQcjXcRPJK2P8OH+zY2DrPJbEGlqVAt9KzjNEh854Yuz5
oeewggIOA7iansuZRIcmYIe73lME+urt7CZvoA7HrhlQXkxuCQ4uZJn8Qg61DjF6
+qgGDWIAN6rIudcbg8P/qWY1Gvf4wa0b028SESRCql9a+KT3/yHJ6Q7RZ1pbUdS9
qIwZqU9gq+QLaDPItl4kw52hvpLfZJRxDJwplJsfNR5KmPXNdqWgIeTbzGFG2A57
Lu6zATxoIE9ebHrykSezFTodLR13mpEavpxZn+K1Ul1V2RMbyEKjnhTrvyDH9RJc
IvSnUywQyLtVlrP/7UnbFojuKIY9YuMBGv6AQaQz3p2XhVa/ApSDoT5CgPIKzdY+
1GLQHgQ2FMaqGXw7OdzmHa8dK7AtXX13/D2rXOfq4PlpxEi9ddiKGwgzkM+H7u8G
bIxQsX78yNC4i5xkJ/jeI7BdoYgXjugowRWo6pXYvsef1VKm7nbe+zlD9e+ik4GX
inKR8ytKcdSCC11mS2MK+xodIXQSVWlVZ0kVZfPBbAB5drPRrF2ypZm3Ib6f7jQL
RoU5IfM19eUsbEJ572AnIMQXRyf/4YPZc8tA9QwWgxWQsWed9mv6a/NpbN1NpOu2
Rp5w613ToM5XFDjXjm/+eNW6xI1eqAaKky73YyvfhyiEzwE5apUUKFL3qWUSBaXY
Ho/xGXHFLC0tH18pXWbJHtoJDNnXAQG88jxWUZ5TukZKypk0q3xsd+IvUk1G2Q0w
5p/UGHkcHUT08of9eg0IwlassHyaPKvEbiDZTuvtOv4a81VM2DsHmooTPxFg86/F
Xf8KkREJoMx8sfT30i/nNlmv7GFwthcHrxA9H/OvYfw9L9xXg2Kz5UZO7RRW5Qju
J5lkhMekfB+DUqaf1CDrWDDJA7/pY7CJrPHKNzZuSXGR5qNxqPar73TYADWBo+k0
66RdddwOnn4jN6i903veGKvHHviQB0C86D4e5+XkTXtt7JytuMH0BracbSSf9Jg9
p6hxtn3TAluKFiOAKD7NHNCHMgQXT3iYee7RiwBu1oluEK0Yd+91dlWK3wgZLrnu
yAUz761xC9Be43sR6/XtuwZsuuQgKr9HTYr7/67sMmYrooZvmj8Lww1NGTTBdq4J
u+dPncfgeAKRXBBt1pEXG9BvtgB/IeYN88zH1xKfx1w3MOPhCes2yFboyqAJyV4z
+JwD69QWaCFygexWG0KINM+H76jOA1BQRNTbd+f8XJ07KyaaEUvZLKs0ui1hGeIs
uDzZlg//mLVOqo1vqPcSJo7L0l3ajSnc3408RwCmp6uXlloD+lK+AP1PcuKvSVkT
/W4yhV9R76Ge+uKL1nDbZWzE6So4D5HsFBd23h1WTX9wvYu3SLlyZOp5iS5YSi2H
4T0Ig0BgKzad3MqAS4oOh25O3mgsZXAaPh/HrwwTNElJpIJ0upQ06bJ0x3S3tPJZ
vcRGq8Ky/UPfR2lZjfhYgXpSlF5zwLqnWnsLlcKHZHH+QErxj2LUoowpOMh09uFz
eBg//RRtNjnHlQg9OHzXYREYr7bPORIAtyEVI9zEmGawPjzdrFxn0oHR/TqQe5l7
KEVQKyucw7WAcWMxQUuNVLyhfp7avv6CcB8SBooCFHVAKm1dZK/8lxha7fRU6dw7
OnBNdlCEGOK/AqGtnRw5RTDzay5gB1fzUsv/CLW7G4cSx4zNytVcFz7n1hUGmD9M
9DQxovWFf0pWQRWY27MTkQRv0mUnSMMHErDCAJSfeJ3NTglKhkfnb+Q8ccSPwoZz
Q6WaWlmbi3+zw0EvMD6QXDmYTlbO8b6ks2c0CaLxbpKzlYINGAS4rshunNm4udr+
i/z8TbtFCo+92YCUWSnp/qVxmScehUbBTfsVho1soScO8Mx1kAafzqsMDKK99OdU
v7iQyLy+NAUW03sGhwwLCD/2KOJi0tYemmeoTQol3IB4LfddwMQkQ4y0IcGLDPei
goXfz4FHhJPlmiCfwg3PZ2G5PSs7CZTxW9WpUPBj1UTL/P3VAIeSA4ClTqWhcAct
C+oiQ65lQbwpcrOFPbUBHq8kxKzIVE49LnRtdZLibs+ZWtEpsPL29LmUUyKeUHVi
2AJ3/9ilXlhL4/yGSbDgdX2NgxQI5OLsbUZOpEAML7SzDqIjYpBD809iVL/O+EnN
NK2J4meIhuySVG5U7xJL2K4aO/EKu+O2uxrpcy2N6GPCFtt1Mu9Y8PzWUJG9fGL3
FkYKmQX2NUhDtZfLLWmQvDwRqIdGlmIIkTACrvwuCCXDAwL7QCWyhDimf02LJXdj
3EHcqveijSX9E+QM+91VEg6WHpogCbJU6KZdObuvXbONIq+o32ySXF5HLaNjnnNC
O0dA3QFcKDmpzA0blnVp+ZKTuLlRyXFyj6wxoCQEnWWiZ3B3ByrQYG0uDbeEqwy+
JcBj/m630uQitL657qKhQF4VwqStnvxZI7VkBQDSzzIxZSLfB0cwBf97LibcBjsf
behBLzwGKDGUgbUXC2zFd/ArOy9yACufnkBn8hFR+w4u6qIfiHewkFVsnpITCgqY
742rib9GwxxwvsIuSRyeA+T5MMsj0vsYtyWjjepcdu/RlOL0CazigxRp2zCa9IUr
GO7GQOOFZLeDXlXZQ4UFs/dEgDHrnZIjdrEnYub5u8KnGWYUNeRe/kxklHbSTSfr
oPnSyXoxvXr47K63unjZhKUjqFWUcacBUPwiXzV7bFd+pkg2qBGepfW11qgMir6L
Ln+vWCvTdpgIJeDIWMYsWsI16o7Jv7ozP9DxQqV0ov6zTg8GLosH8x0vNqeIFfZH
yAsc7+BqGp4fqogEsAOMrJKamAuZlx3sUo4oXxFKjOku/6c/utpGAWdLQSuuDUks
yqZovTAxhEEYPEd/54V/lIhrxt2l7m3TfKVnBcJxzWYT7fEVxVc0mo/wtkrxcImD
a7ibjJhqiX8qZEZmP0QUBnIvTgkGzjTqYMJuUE61Oxq9qkoDXEq8Qe1dkD9AesKw
rDDAoa+INnTNK/lm1B0cm6pTu47TXHa06FcH+vz6NeWMbM9WP3nBln+FStsw+QCd
2GsxE5cjxPTHV3llDa2k5gG/whyxbVjEqvlPiueqdheUPuDOlsvCtwatTFJVX7Yd
2ZPFNoCLWc7bVLaSbMk6avOe528cHkBv6L+NY6Kixa4AYsvIY96W/g8S1GYuPHLZ
VDYtS32sW6NbRe+Hkbk5nN72GHsaOvm7Jp+GKV/IYqV1Lamtmht70YQ2riPOkd0I
DJo2KHCj7X4P/fCaTFoYSPBiWRe2pZ30uk3wSmuNEGh0+zVGsGLIDlIpTNaaDd4T
wKcQziAzd/CtukdSFAOEJF+i/tSdYsKk0xqjkFcPMQzGJNOXvS3pOGuE54n/0wEZ
LnHg29ms3hsdm2PyiIa53DRkn8XqG7m+o/pAVkKbQDjknrBnhmNG2VMPI9j2Zfmk
JitmfV4LyA6orxX42viyvZ2Ap3eEDJyRK2B0St2cLsfl8YnxsZZQoxrnf0MFuJJO
MOddl1ezKlvDqJucUjSi5N8L8LltbBCmjtswHmKcEsi7ofQ0DfLv4Z4IblsPvpzL
mjKiZ6Uxs5QfYXbrVq3OP05YZkFJmQ1UEbbtndatKI4VOoylfh/qXRk7ZKrITDBL
nNZ+8fuvK+D8dywSHTGD2pquJx6e+gndvqr3LY9pe5G2EY9422jxiir6jzVR6bnd
8syRso2pVscH7sxRkjNQXVDYBQFaI8ToXmRFWsIWTyB1KhKV+Rq6Df7oUmW6fDMw
TfMbPeKGYxpEJ82mV1KwiZx3XEkN6QLZjpPq/+d9PzDQCTloquELe+KapBp8ssdx
Cpu4nALJCdyKsiKBQYBbcTNS1mLC7O/BiNjbEdPfgexNVPU1XuPVQauQmaR2d2Fa
oxpXD5Fb1LMnsUNg2feOVv9WZhiPAjednIPVDD0ATxTL4bfpeQAm860Gj4RGzfWx
RsC+nL7aNOPqauNa8kSmICcMEBAge7fl1Tk0/jkr9FtBRBhw8Jez1XQKs9Hc1PLy
VjLNinRVpvdnv+6/fzE2lRWSby6n+Qvf70alrCYPkR3EvnIz7daKPedQVEK07j+o
1JDbThOUb4l4Y4YeNc4dKAkJPDKMwWPBdV55c5dvgwIe2JRhgUsVn/m1OzgPk3mT
hGVllIvV6KvBIKSwTO8/IDNgt2u6RbO7Q8kT0pv8DA7R63EpIarg0SVf4iBQxYhv
SX0jProrc2n0m4P2agAxq+31rxbyTIdtFva38MszVGn1GoZsDOUJDvb1HYBH8n/I
t58/OY8h+GfDOzAzcWOkRcSXJLWXRy5lzkyEf3fBmLY+1M8ywPCQ9pWTeO8Gfp4x
2OhH+9vG9DRr7dhpNOOp6P3vtvAc8/L9woO+kGGvtYDDqhyoTf0DuIwzssawH4Hi
3hTsNzRN6kDodTPXGbf1QCCUurkeuOxKG+Ax60SVsqviBsfmqmwFfT0Gu2LE72ia
6E2cGUdYNrwv8uZAmAYXof+UOd9RMwwhoYEnTmoANiv2p+XInVZ6hb2CYwRWET0G
jQgJL71vuasz2rJQ31sCI9EpumeuBcaICJ8n8s1mYbzZs01F+DbeWLZNMgOICxmb
cLeK6c2QzVTd7Hz1RJgr3jSuD7EzJztgJw1QIHxbbRST7buaZ0xMQE75DEFEfVrI
74NAidAFwkCLaL92+mTKgXKR5x/EYV/hM7ykJRVkpZCQapWZI4Hz9Yrz4KODikOx
hy37QZlL8ARTV3P954oAtwkitrXuxIHOnQtXaaGYENTGvIZ/lp7hDQN0KIRdyDZy
Dqh93zA/NaxL31u3RWHPrVTVoftsLkcuB1UUYAOu+E4YfGn0+7Bcv/zbQdJWfrQd
a6He4b5wzm4cBx6R9zBKajp4m5nq7TaOj2X18dY1F7O3mHfxwtnEDf7sEX9RhpT9
CEw3dM+USYPG+O+jSKtmcb5xyrOZw8mMKTQEFYwj0xke7ORfnSdBNktmqPMl5Ixi
tMba0AFIdt1GeCreKa3wCs3DvzSBokisjCrf3lr98CSDJ4ibi9ujblG7l1qjqM/h
psSvCHphbbf1D2zQuPKKOYk08UA/HFUwwxiMwy6Q1pLcp9cND/yscSEnFS0UWRv4
rJ9e1ep6olqegGew+JSwV0uqJ2E5mTcAsvKDmk4ox8mRtSsEtLrJ/v678f5ZRbqY
2cUvAgigusQjsj7i3VWk7HatUZnIWv/N7tL1ibbr2ocu8EltPkaNjGpvhAovk5QU
/w2tvqWc3ts1SDgDXTcv7MstKeMJzb/ecTHcjWJliEwE7BLhpqfLUJNcK3NqoGDO
/sUk54tcQJUIHpWR+KWeOO1TsCYsSIPaQhZabszXPpnKW44ttQSz+zMW437W+EYf
aoYAS3zHjkElAr15ha9GBpx4MZxWOOhHIe9N16E4Nx/JEP4WvQFKoXjzgb+m1yf/
OaoqNR/wKdHk868CgMWaDirZtKDQPvI0gJONHnp3l97TsejUJledvDt0UQVa9Pk6
2VKmPICRAl7Y5MFuFnASN7O3uhogjxbVbgaWIcuylV1Ko2uEpBtYhW6fDaDNlyMb
NVjUbwJ5JXqKafk7crKSDCA4fBZhBo0K7VVJ715DOXrIU5110b+MQsij6fgkZYM7
S0kPywQo0AHRWbPdv7uSLgyY1ESNpXmCOlVPNaAkU75s6x2wr7Pts83E1wlHt/KZ
CdMde4guPrb4WB8aIMidB3JNS+qyVh9dlj8OfeXshIxMDGyELjXgpr3fNDkky6y9
ZTYwLlAAXSXxjnhQjQp3YRDOREo3BfOdvHKgzzGiUGsJOBLB+jLYKH3c/W9HQHDp
upjWfcvr8skEpUXcj/JsXvFLsOxhSRJpaMZ8CpLYdsQmgD49/zqMc5texus/jkHP
2BWPog7N8fcVhv2kKi8M/gNDgDsAWS8/4TnCoTmhZdUn9v0RiFedwlgRPvpE+k3t
SvFjrE38sisKlohMmtQ+B3MXpk5N6j2ptcJSLemW4gcr3aOPDXhM9X6xE1bmUwez
OwCFY0CXOMjY1o2RkXdF9eTUsjDEXzcRIei+JA75xPvDBosEaavkWMmX1H+L19ZD
N3jbotRksPRbH78s3z8051hXmbtcEYlyGR7qo5Q/Sl6SE9UBCKKYr8Yz1Je7hwHC
GugmpY44/gH4FFPLisBJAkmUZGNwg6KT7KLM1cA9qPXytjoFeuFC7/v33otLMxyG
uBvxEIUkGIKJulEeveZ5xedAUOKqW0uHdNGqfbfUuLvI41M/UAJkLATKceAOA6Mt
fYMPBymz4fMDSEyi+tzOy+8kkWmntOCtQw+tTyVqsEjinkuVnXZNOeADcpdFzcoB
7R7V8e+W9KLfrlijKbk3DznIztR+Wdx/IqzWo17tXIaoPK9Ycl48bfLn5f5CDZOC
Jc8M6Oc8tcRfUc5WAEthwdpOESpvq2tcOfacU02Hity4ZUB4P4dOZk7YpRzmYtg6
rszzXQO/5nlCKzc0Z28Qus1CHRj5BUx3QcZlf1hUv8MDBIa1JqwHMiO59U1TLlyl
Ef1a5Bt3WogQ9SGpBB8Tp2nKKiRPH0voE6G0tCB4BaoFi7uHnmLwqyXfSMTXUVf+
BjEqPO22P518ciDQdL+Aka8RqK4muLMNavClGRF4y/Szf+zfQcoNdSLEBUze6su2
amKJFjpaAjbx14RoTiNRchJKo0NiPDf6uYgwKEQplMdvnyZ0g9a7hhYvSIdTLq7Y
a/mbdiSpt/x0pbvSKC+nMC3zDONlTlR7VIawY04pwF7st3sVfB3ko7MHyA5nP6Mp
Eb7z02uTb09UoxFY/yeH+pCh4NhbDQwqNvWm1YiWW4kJxC4ooL8qON5AhHDTKhDs
8ZOxBf8uWTF9I8NZtY7X4O8XMl+a/mY7Dcg1Kk5+x5zA8CQ8uK28J3S26QH8Bkhn
shmfjZ4WN7k7IzvryAHFwZPzSHJZQ5w6KyAR90R7RoyPZgiU8oJi15CNG/J6Y0Iw
KN69tkGu67Oiz8RzqYGEVhyw1qPVirg0a4s/UlLQlyHzlf6EYQvQGB6idxjzviDv
pUJEQQKKMflLkm/ZBV2z7cE/Ak3oKTS0PUlQmTqr7SnxogSU9G7AiHeeTqkYBwPy
7W3UfpLM39GxKn8LCqzsnwbyHSVEkGpaSv+umeJDzwCmyVwC55ZZpQAGXS4XGmBK
RGEjUde90Mnx5ejnatKJeNRHmkl/ygLmxVwuSUAGNp134AN+UTG7WRZHQ8581HQa
erhI2noi8c1zYBVLz8i4xvSAkG9jRfAtg4c1LX6EYeM/tfbBqBX3zb6TNmNhMQH+
YPwzaWIso1if49IYweky/gWjk3LS2xy0actIygpfE7lrziGgB96fLo3cKajO/Aan
ofDaHyDB2xAPE0v6+/+WG1rI1dwCRFheo2Rv+hBBnTaLE8kKCWhiDCBL5hyTNc39
QU+UoPb2CmoFwu9BJomXLpnZqnCxiNQwcYqlba8Ed1HIF8kkprJbUZXva1zbtkJh
Wl7ioL1cgHJMe3gKKFMogswKGlb4vhGuzLfJi9qUk6EjyWaIJpRIJm7GRIMAhL7Z
W0p8l0+1s2o/loTeekcJ5wddm/wMjYY8vGZn/L5fBsuE9LOLyE1gCnvFL0WWojJA
oC7TmQMTZMbzlaQid42b6UYiscDar1Yu3XxvwbQx9yhFwRxjuzOetT0TfAKd5DRX
Y7i+lq3PEMd0LkwcMzm4OMPe6Qa5ooArWci/DdLS7X7wHb4Gq3+XWNNm+B1s4/9z
eOES0ZoMd2VzSmhzq8ZkFRROu115sYYjdguMB3K8anDVbJVGmYK6TIWo5OPK7TpZ
cf9bsv77mfSSgwrZy57pe7lhTFqOuY01W2z/f1KdF+fMLpmHVht72f9rJoqKCl8k
XwSNkMJZkMeBw0JzdeS5Av0Raa8eUU5fzpiIGCOmlk/lGu24d7JUmJEUuCjekHVW
NmcCFb1t7fSTkEw//RmuGZh1lLNI5RhcazhM9cM+yV4f1bI/kKbpr1Dr/k9C4Ss2
ntBoKtDqHS1z4obupBlc0m6DIqNDVGJhTFIHDpOWJS7UijMd3JjkgBiMelJ/L+RB
1zl0g3tljg1QfLsEvZNNF3XBmTnkgb3ST8MXxB/qDvHWLKLF46kao33no9w9QRGh
jS0L93DJduf//s2T4rLXD+PkluOytPFW+PGGSg3Obr6XUA2pSiIyXg20y2dHeEYJ
uvT28c1DMkRK4TdT9MLzNSmKh0c62VpnUFFRxtsaIFJoWKKSDict34wiTN66cv8k
A4C3vpnoQ7OhMDJgwS/49tw43iSdtTk/3vrdtp61KAltU9vOFYFWjTZ8mvmypRO7
Ih2963Sn5s6/xazYiNmq8Hg3O7D7CWZ/9Ue/dzd9mKl3JgvfivRovAdP1+HcMzQg
OEu6CWawTXS0ZBsOEwlxFuOHFIlMTJ6MEIzBWMCauTT96RCdxgj3/d+0pseKcZ+Q
PekZGe7UqTcw4FseivKrLUJWtB1FEd+6qU3iUuGT7dWvPVBjZaGQ7YD+fFi+DUMS
AdnBob2lD4JxG8/eDVceyJgPJPC6bsWi/+rKR5rvxhIcTpi97YEZCMIrUFpmg2Td
NX3L5tvThHeRRsSqJ5wYdZZUX0RZR+mjPK/5owbJ8WxEsAXnMzfgvNeRxOLlpgx9
JIxpd7Fr3L8lD/iWLmmf5mgYQZA//kvyV+cZX7KRDC1qZyr4E8Pd7jitv2IrWLJH
2cqERRmr3AeMXHAujMMkYNStWPWjc5Y7ehFBPJASmjXYxhsK12FjegbJAztYdJZv
yJZwR9/FRheJgpykDPWRQc+93upP2xL53LAuIxH/ZWnydNPoPxIFNDJtszPooONK
aDBuywa3h8gVqdxMJGrJYeR213Myvx0UbDWXwyZ/06toPXlOhYEW73p3qafCEr8m
WMdkZpklDRVK8/JAwARdOdSFJxuZy3K9oDZIdLhph4DXK7q16YUIF7s8jV5TY85A
VxuG38OrQ02GMvIuCihb7jniLh4QMgI97Vg9RcBQ+clRZmTCfbEIjo65PmLoaQ7C
Y67QypFKh/jhy5xWqCwGE18umiG6IQBCDdJuoyfRAQ59FdJ4qoKqSPY8NG5ZYh2U
ss8FH2YNjTx0/T11wcxQ4PSzxvwMRF7eLz2LTSbSDCSpNJ2tX7X9t8hbbGdjIQwR
3UdG8p05Cu+wuNIlc1qaf0m45rS1yG0XlmtvGm0cHqMVe7Rm6mTdy051vJ2/0MhO
se3zfPypExCtVUcwdezfKTBzu9lz/12j7JT0CWI1PqdjOdWwXNSdSCxzMLL6Diqj
GZgO2RJitVSocoM274GHnPY5XeZ03vgATBAfvj/cy8NHvMHUctdXJ3u+vX3ycpzG
MNe0mZXlNnlB8+LMsp6Bg8GwgFzklrZeau0h9nm8++P55CzIkteHYNaY9ZwhPt8Y
8JvWGB2JlsmAZawcV/xM9ubWFaYxRJINn2x0/29X4seHaWNGUn09/qnl/xs4RChy
aRiNnRVK3KaxgdZyOr9/TewPm0R9yUSzPZXvYfBOGoayhym5PvubeQEMEsVbP+yz
chsopVaw978/LwTWWGfQ/u8yijLsiwFodL3UzC3KytKv+H8JF4mzdM0yWNDbYXP+
tl0Q/PLHkXww2mgKy8wJHQu+nwNWdnz80RQGyyJPyeDaEY2JRk4G16HgR7WwOv0X
KyhZQes9sEe6WfQikzythXKVqe0wqyaol/lFtP9TgLR35aZW637eQCLnkj0YX2Bi
NylmqmRlSsh8G5OMQXaVlyyS7UtiAVXDGw1BS50Jsa7PxBDiyMzJSf4xxr8HZBYN
CSigYQFsd8FPcpo3Ebu9VTe4pQH9IhvLc+acNMmJVkY16pihbOPjpa074WxHgeL5
dbGuSQZi7HRaBpvrSbOhp1onmYdIHOy+lQXURCPCKdgICqm5OXkegO8dpqNy5ceB
vtyrmbwPC42QKE3JH29VPHVbbkOV1NsbfZYbnmMnM4fr5W6lGDQ/6nAoz+7HjoGk
/m805dJq22gJmKq60JYGsehEiQb3a8UCyG8xbRHi8eh3jKk1KY38MLKD9dNLJx+Z
yarmNZkU2QoftpGM/VUo4zKFHZ1UoYlLn3f3O6T7jmfbzz6hCYR4JagMvPb01W4F
t2H5G/FsWc8sbOfHpvruOfITF0IrcMzSXafMbVRA2r9bFJaK94dv4VdE/vzjADQx
467BFgHus9CHlgcf9Bknwr3cWROgnvDW6bNudCOheTngnwbBS7RZkogJq56t1GtI
q5+wg9gyBiCIWSNNb8fC/KE6RwsnROFEUqW6AXHbmbQZ0TdlFYg+jAkrdaPO4WR0
CQi3LdI8rXO0T3PbysVW8PhtgEcD7eqmkJmC8u5WNsQ4fGlHEUWrpHPpDIiDhzpP
UpHFz3mOs4X0aDzCebqfpifCczKVx+VtXSUPVwDt7FOlaF7W8w90NmaztHp9KvT3
f6C0Uv28aHgQrL5o9gsgbdrZUwMF+JG8wJ+dxg1aQ5LMJtajPIJCN3fI++CbfHjR
2MwzAJmipbmokTITwMSveoeAo/xTIu36p21SoU3fPx8QvTpCzxbUiWfhfFY9J+qN
/sbbvB9cqZPHBg7ZdmT8zEcFvTk9uc16MyPyZXNPKqfTwSnjaVXn3YHA/dwa/jwg
oNR2UuJ//Mf8BPDWWoR1dqjbthOFQKd0XbFIWzM1EdV85FIGiWqY7+QFK+MVkezw
IVtzhjeHSU3IJuZ7DHwEq7fAlSpszJ46MAi6tgLwhWzQpPKW3uhrysjNHm282ZTZ
jjgr2A7GV7TTuMBNCNyT948cWvX/EoR1reCbL4elGPGH0NENsXlKizDMgwI3aHwI
GxIKOfYsTLyI9qhoRDOXiPcjvZFhw/tYK7TOnQbRBwK25GDPAGu8F/9+AJRjftB8
I4QIvHtK8kKGEHf3ng04Zo3zOXnHFU7xbD1XEy1HDic2OdKA2kyL4aEyFHHjR72U
qYCCkbMdkFoTdhnVI0F+uaLDtffpdqQ/bwCY2Mfj+YGtE3TP+uJ5xbc2twMha9GL
sDTQoPbF3TvjtONAjT5PHSofHmy7FNZlBM+6S7m1vQb0ecdjM0e0Fv0VFb3w1lZ8
W4jrBHOvVX+4QyS2nFcWSGNaQZUXEWW2ftKOLO0ZO0rYiT7hlYlwL5tMZBY4mSRk
5W/GKd5of6a8SYQfVyVTymbuyxiccp5R0ZmN/uqpP450UL5UFKZJdaQrJ93UZ83A
IGqAqHkrdP/iv3eyodUOTIjyhCqD5WcJC0de8/r+D+6734MbktHC+EzbDKJC+bZF
/MRCMjyV99d4ec03ytB+oi6SU2brYft0I5CAEmomnz0fAkL00cyQbVplfdwxFWcp
0ZV8kcZlkjly8ygbSH6ADkA9KLDqAyxubi2boFj/lJCjWK+h1mfrjfOJ6McWZPE0
nfhNOjzkac2k6aWycZA1lYp5IB9+JMeOhKkYk29w8HKRWj0u+aryEyXwZ0u/Opf+
qqzDBPZtLgl5IzKEa2s85fzNQ63TLR0WKlAhW6gcZYmcs867u/ogy0BGKbzDYSFQ
6+V2mR5e4Slh5+7d0JiAv0emkYiN1Tn4SkiVcfbxH0ftPXqTHqa77Adn4y3n1I3+
lkjyEZTcJh6wqsv2NcVvhiiQ0G19/ON3uemIRAH0UYvuWo8xEM8dEXFJKye5Tdgg
mIVdax2Tf643YJIFammEsZWB0mY/tZkVdspdwpbEOk0MJUXw+mkt14My1sAprNgT
V9pimrMwIcvLpqLEWBIzW5ujU6Kb69cZbtEpK5tOA3caf/jxBdE4UinvMTXEIENv
4Mpf4qmyxuBU2WqbWVyYvQ5ps8QG2ZT0NF2zHtq+dUYl3NXBjkCkL3EjI2w05Ltz
VuYrLTDHZI8i4lAYYN7Y4elnZldXzZD6uLVgeJ7BafRxkYg89Knl5gxCUxGtCoC8
5LxjrsMc1EWGV/Ho2S3IBCFPH7+YxEtHf8/YJ/9GdhwVHuLEjmFei9P62HzT/uws
XAAIFBdzrtaRyoME+52L2hM6Rn8WwIc/+HFmaWkM446aweuXEsx63S2BBxrax8s1
g22L86g3D4l555Huj8kFHQoTfCfgogD3Uho7DiWGraKEN0pzj1+dtm51+UnwPb1z
TQ1grRrqGjeZByVwN2XKTWrD+rp1UsYXGm84PGQLKi3mnVKaO3rEyQpR+5yw6u4M
JLiZwm2q+QkOtXnTMpjxJMrS9xyyaf3QsG/bTmktparrIw2mu08XrHvz8rrJlKQj
55nnYUbseOGUS1Y9Z7WX8+lphB1xNIYyZ/paORdv/V6zwRelbDcXKgMazv+VllmJ
p/op+WdFH3NSPD9+lKoBM1qT5qs28RaWaLxz8oB1bNg3eo8vt34K6bTkQwCdH3Cj
FybkhOV7fUAWvH3OEbeS2gEO6wkjzqTIAn7zQ1ub8gyhMGp64DyghA2dG4wNzLzP
Pq5CNRbdGWFM2Anaubx9esSqWZH+M8c5igX3RktrIq2O9fPOcf4DYpP81aI67kdt
HvItyCkV0B04CkS0Q17vcImNOsvHqkDeSnt1ln6xGI1KzvrAUUcs5TevpEssva1Z
4Ke9LZTStSVx9SIMAFqcQ/doxT36dm3f5QmA4HsBCd7DpHKcoSl5LSsZZ4j4LQMF
58Ifvd+rTnnh+llEZg7Do+kF7V0ikWURQfTxaAlh69zpXz4SVqD/0ZI+gPIlQ5m6
ZA+sjciew5KwFcBhH1awbhshAwwrTCFFx6ODsJgvnC8A2XJ6L/+p+T4ve1nurVQK
2mVc8jiO/Oef2vXVqHWs+pkDYfn6zJT50FiJbJLU6jPOvr+jrpfBTvvOOzDjqLvF
rWzkJtXNvFeYqDfGuiuUIRh84lslwv2tMpfNlnTKmO+/sxS/yqxyDCkwU9V8/k1K
dYynPNmhrh7SqFyWg5OJm0twP1Qnvg4eyDiJqffW/idbd74uHHL80Alz2w6Ykoue
YM6ddKH0bSEyc6URh0qDqPaGYzCiQXsfoRMVr1Na32pxyagsjYWcK5WN6iBfNN0O
eL+TMtpNzQt13EArZyw/fPWMn5tHoHB0g7gXL12QFd7M5SI1nQUakVCNjj9ThXun
xYDP2dobQhiJ92TebilwT6N9E2sSOSqIAa15c3sRM7fURIZ3XEUgUAI/RjNBdGeA
CZJ+uYa+gqOkwimQgKt3tXwmCiNXeqZeRN4iaYRQF76aC1nMQHZd8b3gom+RdBaT
4qL2c52+7u/Mva4NRNkzVGq+hLCZRZWIiGMpn7tqGv2tcCOqDcC+zMcvwLqFZwxb
+YuuMqmaBvFv2k7+uVHBBrZxcylwJYKbMuo6QRkEo4BFTCmTveyrGDhRz0rznu6x
3JA9rDxndKbCKjceloCcMkhzDeyGsS1biFcpGC0yTID0Oe8PHbezXbO4/4AMZV0F
9kuPuisH3PjD2wGDEq3yqdMmHPpFA8fHTF7cYZMUYXKANhxPvkDqcX3bv1bJbO5C
vzcTmazBAe/VLQjquaK+HQxSC5jlsHc7kAHKYRNfuQl5Cbd6lolkhIcH/IENWH+f
F+2yY08LKVj37D53deOIMlkIAEDsSWi3QHmk73q3j6d2d31CGs9B6r6CMpRDMuDK
TmmBjN3fXOBxGVj9cm98FadfSWHiKBQO8HE+Wjqyi+ehfaD3eGfRdUFpJaNf0uZx
A/lxahpgYKGCa32skZ4T1yxu28qOALyr/QMS4mPjR9MjX8kN69196iSzel/H3a6I
a/mGdZlaH4rjT3Mbi4m3J/wbkDjWRaEDbAThPiDmIcKvUjvQqD7Mh4otrcoDZxWz
J5z6LxfAyqL+Cu7UhFk+zSD13qWLlqEb+CQn+FZJAVCas+mSq+wwrgS1OedkaKLu
tdQ4zFO26x4yDU1BY1q6hVy3DRS0mOPZ7z/tT/YyMuKPtoLK3X7lg8va36iKrIT0
v4lGn8c6JpSdDg66g0P7nk2m5iSJTlnV2ysWwgHqiLGO0fVSl/FHLEq+Af/m0l+l
xVRjwvvD5G23U76gJA7FOpwo1MGLV+i94VYCOFxMameKUNKqIdlwfRWvT9kWUoA3
SX7C8+hBxJHe3odTnKyYwPx+jvsNqYs/o05RPgldWrITsYleiZ/+xipyVshydbgR
kAc86PIRQ2IRTAaw7O52pTn0ak1kaNw2WZRD7Q63cLf2gDb+CuNAGWvyZcGQnDDg
C+r+p0lXPs0vsprfhB3xTK4rk5I3Z8d6LCovjiWPhStq5t+2ZJB3ApcWwbEybqTK
06ZBmHmE7RkgZNQupzEL3s1z7HmUx31S22zwo2vuUzZfC86v9PuqukoUsSGymzjN
PVYB++TSj4UqO91ZRfjSLrRW5M68kb3NzJNO76RdXe3Llq9MEvDAFEjZZ62BL8Qm
ku4tHDvmJsedF0tZqlf1VyMUPijLBSqmnTmWQdzJCej3AXDL8GtOBiGQe94lW+C2
sTGWTOCbqwzoHovMjm37Wdivj2g0mIC6HxMsmnZUrCsMkBWnSmoaAXJz5CNus/jB
iildTf1xZgsPehj7Gn4h5WBlfy7sCFCn68Uc+GWn3mg78BC/UO/YmsCOtdqbjJNP
cr91I1sxvddCZIUgKoiSIk3kQO9HkOIeFrgmuXnx33IGfDIsq8rsRsZhwgLdzOI3
7F4c2FEZ8DgOzwRf3UDbWw1GaCPb/CE59yhvyHasw6hOg7HQq3FdP3OVIXekMX+c
0HoK3lcUBqtySOBU3Zz+gv0FTmvxg/ziSeH/PTeZAsdHSr3bm7DkXsybw3cJfdya
QqbBVoyezILxArI7WrOC3sSTCa/K3ufDtVCOdbtmEVWZGkvTQc3lZ5K+cdv14oR5
CPnhAVaDVx6UBChBtAWcUfCgTkx3xU3Q5KB9SWCcjXngQPWlXWBI+J0n8eRSUX8/
UCeilKRUCOD2OwQRbONfxd6P61poAgnyFB30CduDMdQ95js8QddjsuowUoSPk92o
DEtFaLi/2Kxjw0bEpb9tdCRNtmDmxISIcj9LSclaHRg4olFhVeLcTdodMAYFnfol
0FpnM9XwGHn1uddc+l9ndGMnyp1v9VSt4wLbrplljCR1oDW24vHGqgYrhQ9GvEwc
Lgc2O80e0x+jLB1uxq/5pbLH66mGeZiH0VMB9jLZcL9BM8mDS/xiUvxCaxYAEsHm
q3tWoJmoOwZjHWt6SwDkrMLhZ/r2V6gFXhj0qGWDAJDnVLhl39OkgOGhvYGJa5C6
mu1NudOps0KTdrkNZjQP5IYg2QhT6/SpaLEKEHN8uX/3CSv/it47XaQMsFEKvce0
VUVP/IvdJbX5g7vpHGnS/WEj9uhR7ulN15Alh6XqwksXNeD96Jn08BCYgBDBhrik
li+d4PDo0JDH4xLqBMaFlPqxrp0J9HsTYHtJMnATej7c51iLXvMsb2CthY2vnjlV
nVP7Fmxu6ongpzSzsSTFxmfJSqTpdULcOXj4DQqnc7CCOIePsd3J399DHB8NTS06
tnNdN3lRV3kE2VhPFy79R+2A2tckFgqGF6fLnrUmEu2w7N0XMeKs4DzTPJ1v45XD
NOhPJGQyJcFpKRW4dxc4d6IUiukDlNUmGndiWyo2H/92+MqwyYPHY0wurQjfbqqx
T2dcAKz7Fvy42BWGUSSElJ0R+xu9oyxeTNlaKMJFnUewhISeaR/OxXlnGg2Nuhn8
GcyXa3E/PCpp2ZLRkeWhH4HfBfUdtbWH03HnoyaMV8jDepHbHmfbG6rG6VOGeGWX
+IJV8JOyzjSQPjU1keOHWCTq85w6AMp7q0Gxxr8EWr+9vcM5UmxBQphXOx6LRaO+
gb/GiFE4DRv6yf36Lh0SpPyzHPLRSbRo25IkToredRRR2GdAGIWxQBrXDoGgBm+7
CgOdrYzkSJStL65muTPhJG08OpvE8kOmZ1+VDZZ75Kpy7cxAia+SrEkRxrSw0Ghh
+A2m/JWDiF/MQXe6RBK3WZ3bpUmfVQsLV6ZCVZfTGOKku6uTh6fPbFU0Q1ctYw0f
gEcM/8xEOCXtd/mb+cdaU+Z3xEmfzwQs9SVe7Q5LlOjAh9E9FwlGde35bm6Azgqj
H+XkHltU3FMLnrvOMHnBf1Q4nrSBtTZrAaV96XevFXelG2A3aZ9epEpECJiks2I7
mQQop503DRNo1zoBqlwLEfRU2P6N9ST+SnXxOLi4Gler2ry9Za3nLZk1Bf1/05UE
t9WqyKRitG8crPi3AlnpKfmC0KOChbgQ8t0yHMaSlskJTefdF4yYkl325doB4REk
hwDx8d2yHhbQ3tntuHd67a+dSFfNisdcL1LMPc7IGLhTKqM+ljKfaX/SnGkSJnSw
NyqRpQNK9v4+nKi5dPE74xKHREILdF1zZ4mMn4eydwZp4yqYdqUtoZFehh3gwNys
zElDHPeDXeirBglNj8/MReD0V4gziGhSJqq/7v1I1GDaMW7pQfL/ecDvMFARJIeE
3QUiFLtG2+awILBbEdNBoCNm+E2WO1XNF9q1bvACPbLatZUtJFjAtq4YsRFrVnqe
xbwxjATQYfP6Q0UicEDrV/EH7zz0jhbAGSYhk74XzCHmFJZWVJKqJY1AZ5rGWqtZ
8drniaNGMYev+Q1yYiOjr5VyNm1yOOYflu/44BVPTZz7GH2oWNhrF/MR0dwt4XbE
Bc72TUo5SN933a4OSKVd7dA7xHpzgGtGZURTkHmld46BPJ7pAUM8QGcG7vuqtvOW
V8aGutyQAABdqSJKwz+r3rKrZDCLjss0+9vQJXJR2V1ZkGClY/KfnDXzhQxjnPEC
cf9CyHVueN5Ydu7KIdPsgaw+wRIf1Kw9TMmNNNVJiF6xszanuAw4b+/xpOR+91ws
oJAVtoadNfqkfS2pTRYF+9JzBnEreqdw9fNr7fMoMlVywohgCcK/D0qyeJq32qol
iUqr0ZUnRK/PiTn6emGHLH04GaAeBs341I0gvz3nUX7TJRs+UxK2Cg56aeWdS4aE
0rEniGNXxEw2bY9JH+xO7a1y5rGZ+7o8CMxgrq/kBh2v5beIDN4aPOg+8FM2p4gH
CRbm05zAfSLI18wI88gU6edKV9pfzR6yiMXmcB8V/P6+XHG63D89qJ8mMWq6nUOp
grZFh/3OSUXbPMMNhOublkxtmSA/2YzcVZMmCJCR8YdT4awDqk71JsfRbY9x+M11
lIMXuGkjzswr9fLGv1fXm6CoaXigJGs6FJ2DfNGyzRcnaWdm0DA5VJr+MeCQwCuM
seEYSAEi+NtRsE9JqF0U839NLs5Mea8uF80EG4136ZxzUBImmniTMF0G0SjAmdJm
kKxC+xBhWJFhu4ydf1/Na4bRozOfci4CDNTnvZiULvnrTZw3FdgkKGUxeBqqhQ+v
XQmeaQrCewycg7KV1N3dpqW15zUsH35GtqYHgwZwNpS5vAi0WNLmwmEnRpI9rJG8
Z/D2XPJJY6hlSzXK5n8d6QcJt+AnKjNlaOAhk1ntWSNCEcQ8DLHhNHrTVbMV/wqJ
v0fPDKK0g7r29TlpxfRogxiwJ7vb5lqd19iRriyR/DKk8Rd2bVAr3aLNPG34fZKC
ZBO7vUZPV3uodankPDwy02BCIzoiFZcDVdhxibKGYtMvnnwaC6UPTngbjyH6k1hJ
Xu2XSDD3E12EszXzYJ5B9Rca9oY5lCXGy6zbH5b3iG1Xee7Np/DKjC3ixn4yijxy
NPFpcWB10a5PqAEfDal/pA5MHJFzTl4iXocPeE40ySf+bSFhjO3RwD++Kr8HeT3B
slIQDqmAah7qMslamg9xbgdeZd9FSYp6yvX0nVqEQ5WKTd2JTRazRq/cQDN94CaM
BX4/VJ6+eqsh7irB1ZtPjingm8YNndMXxYZbYYFGouLnZmZZKbGVIp/2VRTA+/hm
cgRuedHvIBvVOc+XeJw8SXoA50ac4hYyUKghlIfoZWnxRsHZlw/UX1TPGPkk6o8C
IcHZV2IsaeVU/Oi1X7Szrl6L9kWA6XgBmKnmPGPs3ePcDzQqU8nyiGDmTlJ0eaND
xFOrqJoh3UQ/hMHYQJKjnqcUBsCCZUD67bCAXYf3QxdEZaHB5LklSiiQl1G9YE5p
4KpcxiasjseiJTYBdWaguRXG/vA6I6ewaxfrLB/YTq8WmRm0h4cqSM7pu9Sn2F0w
9kxQq6VjcXmta99AOAj5doy+y+6i83PfV16sZddcXM7dQAvqKLHdh927RABDNfkw
raoH2IRd3lkFua//QSfOm24Rk5FByFoyXw3XW/1T/3dn6Wz8ohNxJFutbb0V8cLZ
pwujFyDgYGEoDhtO/t1N9xTqePsN+/zlXRMcJHYpm/Zpfp5Y6EjxnIg1AukmqrTM
P0tdFYVPPeUtXoVkCMil7Kuq2yrvLgx0ox06YLkSKeicFH2RxSgHVwVhpjGqydwx
BXxpcixBcV2Q7+HHAVMPDGnRd8I/nkaFtz+Y6i03tRLu8bb6Q6sdv32//CObmTYa
tAjGxYuT8aQkUHbqeDUkDyTrxBHjcXHz5lGKOMl7acgoO8p9lcRiNWXlRAFvJkFm
v0zGS0ao/CBbMJ1erXekDFHqFAVOQWg0csVVFCCQqzYX308ILDGqXLU0eq+6w4Hb
AxGwaZMUIGQ1Bh835fp8c4SIat8GT1HCQvmTtZAjILwYrs+luPvmmuJxYUlhGWN3
U9Z67dGvqNit2OdDNIwSIW7NDp6aRK9p0EDPlRFhph2NbjqhF+QmKnC9hPkzd1hV
jqZLh5WcerIKtd+29y5+lQGqlhq0BPdUJQ3dUMn5ypK1WgmVA33bzbSKB0gTAidh
8GUEGmyKY/7qeH4OGpa7L/5MnVjRoz/V8qL+yULMn3+d3uIrjsLQEfQUYXI9aCLb
epNbF9f3RGsQsi46ndvP+6uOAVHJ83r72r/DmDcACvZOHVeqZkP7VPWy1piirsuE
s7pM3tbZOfa7uFNkqBvc1x0yCNDeacn2kiOdvV9DGMq8Lg6hTXmWcZxLpIVUyyGV
1Ti9ml2uiX/3fjcH8XnRQoKG0PhfRupgzW/v4TKVIb2CnapFbhLyAh+oCbefC9zG
7bfTYrriVVr0gO/T8tg+clKnR2zH6oh/D9y4KFlWpnpJ2GL3XI3mZl4sPC1eLCe7
uDBxVvs7T1IezVLzF4xObtWoPrwehMqxoRJZI9uiG+XyPtp9D1iaQxKWkh6QT4Fd
Go1c1z6jXAHDgR3SmSmw0rI6Lp+aFzqifOiw5NHM06avIoprvLHdLFJ50bq5Ic9h
WyqCRKU6XxUBAiT2hRR3HllqvFyRq2in6R7Hu4OOnfh9ye1Ndy3tZLWoNP1p5Ecr
ZGSIgQWO1XkyHDFglzz9I7KbxRa5M1HzY1eH4QQMQ/dtRCCCZXqpWKwxhI1k04zn
U4ZEDejGiW2Efh9svrQbtJzYDvGNUayYiVf+XnvO6f+7yJq6G8vo1NqoxGplHvKp
8TenjQtFF7i4Ksp4H2RttsppEuLz5DWGLJKpP0NGq2BqKt1i7MMBI9o7MGwBFgVC
wRLEAnCEjsskMBrxqRK/vAQYGbYbAj1Ba/M2LWxGSHTUCE8LlUKQUEmjxWlFkOQY
QqBrI1PYJU2OQori+Ki1IjNzI2HePpYI2Mh4sYLuf+EFeFL4tVVn8993cC/kl+8O
i4/MbbDPdwyKdPHRzrhc+qOBNMkfdLWwho3O72k0nnrkPQCRduMdZA74xVa58RdE
IuZay4McAhuY63xxBnMjjplNzcJSNemfywzBVbMOMdIhlczkg6CkUNHoEl2ovBS5
w3gjABrGKl6sp5rO/HddKDIOLc5ypXz7OBPd20SSaxMjQ1aS6LFSLNQ2NxNvO+qo
Yy6A5QZ821oh/lIaj7Jqn20Ia3FpP0MDDrIt/g5wo7lIetgT2O0QG+4EhsXvcpvu
zRU7tPCyRKsnurkYspT+kjoTStYMkM1hnk+nfykAm2j2oSjN9/xlZ8/D5deDmOzg
6K590QOU6DuFQrCwEEymCXk/5ALIZC9TmdT3fJftLQ6crrceeNY8/FCJFacVMniT
JxpIw52rAmTLD5qApIIi2hBeW8/sl8D+ktXiDj+mdZmRzq5iiCEBgDUaOs5OSw72
bG4v+DwKcYb6x5kqtakMeGcRtvORWGx4hBBVqM9pBHtmpkIfgeTzFJ+37xM+LShD
eRLsyFbCU5YhNM1y3VKNq/DgFroC8dmbuIBtf2Vlqtg0JGPVT2Cs5+GXA9BhKVes
PtF4G1wajolCNoKNZvQxoI7ZUB+FQw0LWcJJR/unpRbgd9b91qULP7mZaUZ6QyRY
2IKqPxGYTwqVPUQdVd16YAKGIPOSxKtSAgC3XC9RGF/XWibtt17r8YW86JWqdKIo
BaPZShyIIE6D+rHwz96URyC/lgYioXQbuwzXdFQvBKU2OIYomCdT96Ivzc3Eq393
AtNaU/Zl73K2Qen+n+tBRIpen2A3MFCt7CtdyZin1uKEPTcwHWCWhJlXGUmMAnuy
ZIp0uvDJwMMn2g5DSgGCaBcJSRKVk0wHCkVsxUPA4cKpNYHS3ePufvsL/1fTRYuz
zq/gl39B1NfGXoGi8Ns9Lu8jnDKH6wCltl9Ad4nL0lY0pkliUkzqwk16UxQcAJMb
LCZquvdbCHF9ZPoTc0y4s8N+mj0hvqbMix6J/IJNjJ1xSM7cdOKHmJE1fvYWqgQh
NDsptHdUmQkMgzobATf5FWFR0Bd2FHSLjQjEs77f24lAMrpe8V1CcU5r29YfkW/w
RdUX3uBKxLPK9OEDJ0s8SWALLyKcY3en3/X6M+B/A23NWOrVCOIChEG80k1MtCUX
1HNxs3rVtRqhoO1Gld0irfq7CI5JN9gJrL3r7QnmGvaGhlKf5IDAXHUVQXD4Aflj
vRXv39WsUpB8ampiYOHeuAfxrECLtf22Qri5BoUBecIXNiv4UtDje50Q/gv7ujST
TZXlkbIP1Q9ubz5iZcwOmdyjRFS7K1ddzXPYZRyzXD/amNCUw0ckAhGpyyl24ra6
6QSQct4uDUNWIMgucbF/dUlMJDAWhfV4iXqBcozd7NDLrUXQXbJ1CsccC2rIPeLz
C1p11NUJxeY0+GBZiDkpMHVIr+mCBUigel2+Bzha12V6UfHTppBm24Qazi3W4mb8
9Z1ivzWsdpWUnxe12tLaL2dbwj296WY2Mh8eCC1gKo/j0RG6NU++yXI4c7Ra32cm
Rcul3MS4E8N2GwhAwRq4D4hVwY3iArGE1qWX38j8a4ahpQY8qB4bUUGHDO09z6+n
B3lOoUEoi9Kg79Y7GvRXOnq6TocMd5buKM9kNqow9L7qM9Y6I/RedDqbqrF269i8
F3wLE3xaMLBWgFMsA48aiYBpm89k8s5+r9y/if1sDQtOT/cHTDqGrZ/Few78me+/
rqZlFCfxvwdJo6/qX+9bcX2j3VZaikb/kIbPArI7h+73541iDRy+uNNaBO2JPCVx
2eKz37rQ68MRxRH+M6iTpYofWYk3uEk+3bba03GRp8NLUS0ixd3smNDtr0jLS1H6
6QsrE6tIL7kg6FUhQSlH6D0JjlXbTZEQF3fTs6QTcZMrXuanCNzTJpgmx5nm9LDG
UvOuKrPTxGOQ7zUlpa2snfCXUs8q0TGVm/50HiOOxVpGQoUf0SnLBGBQuLd7X+lK
+eM7JtebJcjkW2nJxId4r7+spA7rJVTbit78vgsQ2ADSGeLEkvAVV1lREevHQ42a
UOBPgZV+/r/izzJqm90+0Ua7WWzcesg+Rdf1Dk9I/hax+8VoJkLfUJl5B3lms8it
bwP9vfrZq6mN8psZxlyI3+vcRii0rmKxHC7zjFFBd1lQep1jFi71Xq+TR01f6dxy
DcDuVHdkSabalVc/XP7N5lQoU+8156A4f7V2j5SSJ+1rvu0xT1KobvvLk4s9lOHh
pSJsGta52lK2qoTpvaDChbOxQ03FwlzkRWTIErkHWbnkvZkrIB9BcTzGiBS8QhDz
VvCtCpCanIgEwBeuyGMQxFI181gvnhAsI0Z+0Sr93ThImrH8h+S6JjE62Z4+TlPD
0MgaSpHztOfo3/8QCsdSPuE6pFlsQdcgYfV7h9S14Tbjebe3p1XmSsjnqSmyNMvK
5yg8TX2N/uhDUNmthA2v62+dglcZRBcTyKcstSCq6EfYFDE6B0mV9saw/DG9hYvU
i8gcTSYoG7RcwC0E1SpUsdV24r5MB0RJXIs9fRWgEZMmgGpFmTbbC3lkvPj0kG9Y
HUTjmo+jkhOSSbd902ua9vzwDgOTrBxFCfijUN9h+oTiINw9OXISrxB2eXUphWf/
T0YOQ+jAW8EaOtActUbXp2htjiMwrDee9moMon+wniI0sy5Tw7/aQ338bLdi2+nc
LqMy4p5jukLkTczoCQfdTEsCL+Tq0PqZr32GCtoPr1wSzPIu3XKhD2iveYjwn2OP
6KRGve8t0vOkvbPzhWdA8TBLR5QdQO3FVTZIKX1szmibKum7QXryWfj75YIkLrH1
3nrI+X2pGPlt3IpHHNkIrY84MlW8/sVfIfOi88u8DmMX2U8PFM0K2k2MDQUo6A6+
bUCPGmYQdZ6eaoVPFTG1L5S14SWhnzUjd/nMv8mwH5+P22BPBXwJnBxbdB9wRdaR
7FuXTIEVKKOovIa6uY+IXRFtE256wOVAXdrjQNuaC8kIfkOyVpyFUWxCV31gXsRN
S5/NyfMsUfG7ac4l25H7UHoSu831hxnG5fsXZFgRdCUeRUFF9T9jtkNw2mvm1Vd0
w3WmkzaY75v+hRexcGUXUstzH7HL0zIhaAIYvPqfd7yiNkO4ezsuTNK1Fyn3+mH3
yO9B2GSxJeSbVqLQvgIrBr3BgZlElCSCiiFl/2ehtxgp3a2HMfcgGmHP331fUIul
Ps4ZPaToOXMD0R+WVjaK0PW6BLnfmQaVwpZqk6roWe6UCwHtgDAXqhfQhGNxQ8QF
EpKHSRTi3H4SbgSUcwvfNac9/E1GljJ7xCMJYhUAyugocjqgyKK5hho0MKAah4SI
tEh92uAaP0CMQjN74bLo+7N/zy8sTN7dk1B1RSnBo1e+eJccQrZdwVqB3Jtiux+m
TyEc7Q0dbL8xr4KymnH8jVMwJyZIgTNpC4W53TeRBAXqFK4fq0kmG+H4isv+1+Ae
YyhkTCYS8qzuJpfZDMiyLv6DmhMVLF8ctpt+AipUSZTmvHh+ni5LhMPDqgZefFLj
hXvt3t1NBpS6TCatV6lQO7OrOtmnKVFa3vFXiFIcvrpv7L2/cTlfuddJcVc7qVu3
EinSHXRQTDS3QL4ug7yG+dEm6wjdKaDuBP8YX6OhcA3okhiY7r4GNdpv78fueDJx
78IWlKwNIPq9ojkQYLZ7fyJNWHfQMvkNCNOGlnCS9Q6MDTteZWBpj8oMlisJXGHk
rWDwhyQRq+dM738bgS2/1UX2ljDxbOzoxhKrSyyLmDBKmZhjHiWXHh0HHW8fYrEw
IHlvofJrf5IKuNLVOvbvhb3p7zHEEhkK85HO3SVNxaY+AX8FQ3FWQcv5jX9D4VLA
8X0Si8SxBmJRrvTApzuGun3yFoMR3zwDEaBnxkozzp+qINuJnMj6i66TAz2DrxpZ
NQBoZSnX8adjHC3ch+GbFal+AhGDTJ5F1+TakwQ2RhrEQp5JPcir3yx4brYMTBV8
ay3mLhK/3CyruKkENcuFn56Am3czmzGTwNJ/4jlkjJDHUTOaSRi1vHQLeRvd+DHT
zuL8YKAfSsNfU43SpB96EuhtDAc/Z6b/4R105spfcVE8ORq1K5rPFk637YIWDX64
Umnska1aqPxZTRvPqN0KZEgV6bDdBD3l3k73qOwdfiVrQwOcy6ZHXMPfDNTxgY6F
sglKZ2F89SO2Bt2Dtxcy/2A5RZXh+ACrs+shTBJXiL714zOkbnkAHztUpoS2AKHI
mjyVSXuZht5MEVNRig6pWNB7MS6YE7BySeEu8jZNatVtNLLDvehqCh5NVlRT8KoG
gpBZReyxLqPpRwomwAAAclX8WRaFTx7u82iVEUdeipl99uBDeek0ywLbQ42dh2Wo
rII0PDhzCf9hgCtJ+kfIuXHZVBg6C9VFm4QP0ACoDorzTdRQ98ra2wctL8ubd4If
Rbo8n1d1UT1sNBmu91/FNKjyGE9rgSoRk2MHvhVKoIW0yH5ppFvoHodQKYuJcDYL
bNy+81g46VloZ3u1rPG7EuSAngRRIDCCyH9hX6trTEHAWbJEvJgqnPTpdUUsbfxj
HIQLw1qlS3yeBfjhNONBPYDSjyCb3dp4aAwdtFKm9iI6jDEaxhopLMDDobrZMhUu
2p+ZWv2SVvk9sklm/ACcsTKAWVaxGsu0fxrtilB0i4QjolDnWZ7DRjPU4XpdBlqI
gclMqOFfxk/ZCzrPDQ9xm92sJrK9ew7J0d6kakmebyKFVILARDDVIyqkIuKFX52w
v9VlYrN9CdB6ZlY5zBv1unFiFHA9XJuylUyBlxHRlcaNPO0g2415P5wsHOYY7+US
ZpO/inITbhiBhz/oUBR5qBKdI4nBjQZYGpE4rDySHY2e1nE0/tUCpSbHh2mlIOsD
qz5iFxjZPz/T/LvirBAS707JFkTouSQs/8AZ4FxHmT/AAREe3Gbsrkyf15zNW8T4
6BNNGv0Xu5K4ljFMQr5TPIc5oYKTxwueYeKGH23qh3hyeeVMs4ZMaq9O5yClieG/
VvjpRwqowcm9QWh+zB7B/VBv2i77ZJmCLXKjRvIAQGUJ0CGwHTJCPC3PsjVZ71N9
7b4jPzq/04TMN7lH8NQvXFdaCJr8S7RWalGxiNz45H9llBld1lF3WwWUzIAw/QLT
itfAFPMMGuiaLs3nMHCUHcHHSBN1NOx8E+tPU6cLdEzF5Y8t88hMy6Fy13LIxix8
q5ZE/uM2sQI6IXC7ShKxwvLY8EcFqu5z0TpsseUN4wJw8sE2ZcnIJQ7GKJdk+oHQ
ICxt0UHBSla5hW2LWfZmN+FDsO/cW3w0WGVRqGPkMooLB9SLWp6R5hy51mCMv+kY
PlgbAcsx8g8+Bvs0xj1heZSRTv2QeojCP4i5t8A59u9lz8GdMQooV0jMJeaHA9wc
j/eUSCl7ou5vWgouu/dN4O/EAsdrtbN04hHSs6xt5jC2Zec1Zet+ZSUeipXjfYnr
NkjuLxfHKG4TiVBkWd3pX1hazFgVp2VZ1vigE6fyrIYhbEIy4jem7xhN6C3/AgHh
v2vhV8aaQzKpYdaPwZUPHOEZ+D/iEemPOlxy4PhwzV1Qt9cGvduVVtRZ+EjJhwLq
MzPRZxRjY9L2k+xutX/b+A6XsHXOXbQ9OwVi5d3as5PnoWuUHJ19lW1BSJM34hol
D2tQ7d15swpBl24bua6kVcyHLeDaO/2Pdf6ynMp+u+Gtc/1NlPHxWXZNzM1gq1hq
bTY4hTEfGggUXKzHGgloO3eBbr9P6d/8Z5c2GETEuEb8twitLuAvDZbBB7j7zWJ8
5kpUZt6W57FGVyvYUTIt0ihBv6VKajyo9BsaUmKkJf+5HAMPHTSheq31gH3lbBsh
MD3FevpRwFvnqQFDQyqPqJmRsPNchGvxjzPk0qhpIfHQnSH1g+PrL0HZXbHWx3aL
dOPPX5cq7iCrpt3G2SHMUDj2Qk68WnrQA0HmxYn/kz57nnq7k6ugdQgXeKDfEHNZ
tVdUs9+uPqVig4pTpW8QHYCMu6bnoUahMd7i4PxlQe56v8u62rkPCNxPfGEeRVX5
GIhPvVwe2TR9307zrqn554booe5rNbXTy5gn3IS6vwW7XWTuIpFQNPtRtpisSy+5
VfV5nIf9vvg+BeJjxUYi1va1OAGTmeMLtcEAv9jv3SdR0abH4HVcs2DqD2EqOqpk
ap6+TRAn4OPsFGkv45RsLj0q5MCsEzcjv0dukll61iDLi/TWrI34oS9SehPnFG5r
FJItrc172nf7cMbYk40TJxWQQ2tahOYOos2zdP4ZThx61N4QGnJ5IMPp7zgnwbLU
JMrjTJ9CdJN39/qTKtOtXXUzb6H5PW6Vz4wAp18nCA/O+jlWjeiNMgysXynyBBzD
hutH3JFekwRi+m/aIKN4+2vHDFkYLwqeCdmobaOH2P0Sdxs483X33bhMo1JH7ZzJ
wT9/Wy20n3ljruZoQqYUv7BbrPaSpF5hluZHbCysJrcn1XJf6JvgM1ycH+5giEto
Z3FWVERg0c0bHoke1JHGJmHjoOGGdvCYBvUVGQ6+ew4WAWUw39T/j5M4KBrJ/X1u
LLZgv0BgoD5+/Wk8pzg/kEFPIyq4DlvcUFM3vo3OlRuxICf1aeRT2CHxGSov0My+
qqnhiuyXGy45qIm9lDlZSLW+Ab1HwqCgVB753Ilc9lqoX/qMH7PzRoHZkgq/EkKf
n3/ezJ+1jDMn3yKUL2MWbQQIn+aPadGJfvqTOH3A5i31jrxdVYv2B1J7tYF8JVEQ
6n1qjPh0aky8J4VnkEOuY5CeeEMk0EdT7T7vPUSrLhzZeVptSHdpRtkxgc3QoVlL
LbgEmkhmYyVfVCcy32FGn6MwMysmuqPAS6IUEcV+f5yrS0raZdeaws2qmE3cl36/
AEm154jd2c/n+QtHZGf+UFFC9CymraaY1ZOhI4PQtpen96bUgqNDLNMd1b06A8VH
FV55fD+UBRg8dPS4aJOwAUUjJ6693pz/ZjYJf8af3uSS0eZgrYLC11H11XY79Zcb
DgnHYn5JM1X1KlplyEKSHs55ycDHMKiCyitPFtK4imAOjM6G/tDXfW3l3ST2h+aD
V++9pJ/pE4qXzn8sIlQwC34MNS8dmQCk/RIVVlMElFLuV0sNS+lKSv1cpJYtnc2N
NJUo7MJOg3JXAwijR3578v/OUHI1kbSzA9bbOgG173s3CjZnAsByadzpjjE6/ngv
phkSv8FywDfigaRl/s1+NpildFuuzx2kXowxJdAi0ZvaD7Gzpz8205CPbxxKmLIn
HV61Nb3V3swKRQy3M6UmWa7JhzN/8Pm5Tssjb5Fqg7frwGm+l0NX8E+O5MA23Omn
mtmMeszR3YgL0+ieDpB+9gm8kmXr1kgELXV1f9vOAKNVPuYX+uvCuDCuU3I+ifh0
yIJWDdlImyIr1DHmGGzYsitHXG4tW9m67S+YFSHtXXhZcypPqnrS+S8UPfGrJBBg
9PMxAzlswLIHp633vN1WnsCET28kfbD91hTcohZLye9QLDj3AX4smDpFEQvSYA2a
gOjLecJMPhL0V3WMQWgOfy8m7K3CLIyvYEtJ5BZzmd2K+mKAEJhZOvGXy3VpAZ7Z
Zh24J2Z+u+mer6UVpiTIKsg+KDUgVHKGyuszxxKQH7Y9frtfBPMtGW0mkkr28c8l
f4Mi62Tx7Z37n9jf2rpTRLAtrG76dghp+t7WEPDa4c09I5uLJdsmix604oUYqmXc
IKIx8rPZtqIR7ERdcIFAqnTMrCFGCyX/8drl9uvtyT+byHVyUamtlCf0kebG4a1V
ZKAZlKz++HtzdoACE9ZYBHARi9Wb533Su8WEdUe4FzPsrSMdY5NKyqE309g5L4CL
45OczRP9QNQ0BG94LvaySnN6i4lU5Sy19/7+Vouqe4bVG9QTHCqpI/kmqCpoO7oW
lRrEI7AF5JF9jeb8VagKxqknONBtYoDqq/FDURCGIwext1hukaFCWDA5ZJMboxPN
3R1NyuifYTPz1i2oG9x+mT5Jqv2OmssgeXUfF5TBNOSw3PWLBhkHkZOkX8yU31qs
j6zBTes4skQw3H3+u1/QaRBa515bNOOOBkiuudSqKfz87WB+L0iICfG0sq4Ny/Oa
ZLwq6JBochDUKBd3B0738/H1nWWnu1ruFYgMcBJkF5d8wa77KdjbAXh5+Im5dgmK
NzPslbEw/WAmiQslKc3bsIx1dljbtSUFsXLJWEBWeXt87kwlRS25iFhTQy8+nxjG
hqeiM7bEaKvfyOq8GMMX+gN+CQXmh0gQDIuvNk6ckFwiNDLDgsDvzu2ZBfGZi07g
PTZOiJAa85A6H6BFP1xprNKY3eNowlABtIM7kcViNDe4Y4FiFRmz5Ew4TGgeCAD9
xs2JCn2ptOGxLWcRvEXJBb7R4VcBHf70lbY0nQCx44IFcQpmvHm62f9tdWpClYSt
p5PhBfXz20Ha/J/Xi4wknigJNKftckJaYRGlkJQhFLhTgZc8ybUivYz9fIXq/++p
gvJNByDXn7Ktp8kyIoUwWH+7J+rS7MlQELqysfd0f+LKKtrtPdMcm2Bcy0bZoDOg
tJEgyb4dFbSphhJbYMB1hd5J2e6szdA89DTnrQ360a5EQzrKFlFMApDWg+B3dQUG
lGjjkB5mILmg9XvoYCKYuQfCIF6a3BSWK9n1Yr9SzrQ3WF2UoJ3RhbhTs5XPUyxB
5LPe/g0tVlBY8OPJdcabFVHERCFGiu2fRcG5NR81f/dnlum526p4jpisGecxzlVG
wWSVcKJHWZhmn+f2pxKVsLr10N+8FdZNJqsIYCie8yn0X9ZsQ7H/dvgydcuIUDV5
yPZ1rJKxmrW/5/+LS32TLFfR95jpbwsqfxX7UAg8Ezt18pl8TkkItSEUpB8ZZDLD
clPp/QcmyadQOUTnVErJ6/LVA1TAdVmyT0kPUC7gbrfpFq5bhJQNXT9++25d5+r3
vkep5FvTy4CYa9RhpulWV55wfSOIhz2XgE8WfDi8FwXeqIy3IAGe7aHiblHCaNcQ
dOsa9XFR9hlQqTXk+teUcoJ7hpslo5+4tlON0kxoiyGgK+7guCy7X+87gXb9H9h4
r8mz65+wZMakfEBm+mD5LgniWPYOMi249X325BEuJ4Sf2qSi6Dv8Ik1tjFfKWynM
80E/AlQgCI3r/kuv2hE/qeG/LOeIrzV4h9Oqn4Xg7/REiAgZqhW47KBNpbSwPfpI
ZgSWP3AgA1VJTu6/lfO3IpSJMF/rCYfQ8JysGSdypzU/9vLQK3N0NfJ9C87/US3r
CZoxXXFxKMBA7fspXuowQfcS8QKQs2zx/XC00DGDy9duVbKwdfXrnFyZjybx3Hbf
AdvwcZbGGQ7DNZrpmNDCt3WYHNMtVxXXrpGDdQaPFlV5IPvpMUslRV+2GurKZxLc
uGHI8D+KqpzMc3f7L981YDISzrPN22p3qBQEjRpQPPOEafc4NDj+MxBGdt2c0IcD
f4o69/DuBSBCONFJ1rGqtQn75ayk305mUdTvqRBo2TLiV3xdC7KEo/4+S+BSbUbq
eB1+V0J/lWRFCjprXrj/9TAxu8mVTXA2yMGCZ8GwP+V3bt8ctTcn0ugyrorr1yJd
wHeii5eHDmNTi1GSgXG6bPEwcSknMAVt/lLegj63SQs0+loICcexi004GPSp0JR9
IEIj1Sd4LUhu3yAdE5AwYJLh+cnBoY8Gd1pU27bCU/ufZ7YfSCv6Thjl/ddUz3EC
KFI92ZVUj05UA7INM6GJI9HJMRfTH6MItH47JynCyKjZO3Dmv/PVhmiH89WwB2af
XBEeASwpG9xg3enNq+xbWazfk8tq0+CZENVklrykL8oZSkhBrFUcqYWugw2gpLBy
zMk0KxuGcLuwxlB3MRYUYqOPK57vKWDJAK35oDRrFA8jWqD12jUaWBBGXJ7C3+5d
F7kuDZDWsCFLqb87IA8dVvAs4b6V7hKyQH1mlZSdMNJM/nt+BvRCbZAKtflOStJq
NHHKB1CluTwoAiQNuxd26QdtiTBgmuuhne0QQaE1NHXXAIOJ81BU1pUFa1O8nkkN
U/VkgSwPtBd2Wmb85oediwgdrzNhDwo2ta24U0eOEjClupwGaLsLicIsuZXBQmyF
NUv2U1hpxWa325boOIGMijq0FiSQJce8tZrFaUVL2GdHnFGfPSLeQOkaFkB6W9vb
t6MTx1EHxYdx4ojmxl4ONrL/56lMQGW6q8SD+dx6u2H88HpXHhI8L7O5P2ufESHB
mlWNrmHe6Ujj+W4GyC9twVXqL5xsbuHF2PNZ2UH35uKUqmzNzmilXmZlj2Mp92z2
0VPLqF1IE8o5VLPFWh8Rr614/gnEcBb71q5OxlTMAxDbE4Fb+soyhYgV/VISAi7V
YcNJ9j51CfAUsLVusT6ef9ONYI5exLMvOHyNrHXmTL6eaL54/uPdd5oPoDH6J8eD
TN6F3SEZFqXwMbv/7QsQgdMwgmjtLRO2+xpzvlpIpmBcpMx2EG7Y2ufY3NiNWiW+
iFezkLHJ6ZSRohLgWeY52h5dUFLNWQogatYm39naoFlZm2IuDMlupzfvdvnhzgw/
tSB5pPBCO49q+CavTb5+wTcajAES2mSCU2sKWwScEJKNAhx9Dqy/fY7azchkZR9T
dd//6u1mX1EQo+uytwtFKSGctshMWdgmkDLXscM2jYR8nLxl9ODcMWuVDt1RjCjt
tFYB0PZgTU27im7cBJ2fyPBPdWYYs6N5rgo0RTJeh1ljS36RE4nFDI30P9Z18Cey
51TSVwws7rZVr5ySYK+IQTnpy2Qne5MCjFmwEGzemxN2beTKhB+UOu87iKh7VVQx
imUyWFSjLwXIg0Nv89v5KDeOh97/69mY2hsGCXlNBCCIt2Q5YecjqX42Sa1u9YCg
jZSvm5JvcuDjpV3OtfXOrfjQdck/6x+wLUrm8PEPfcR2fOvEJBVt43m5yQ9bFHKW
lgZ+VH6uBztCaENpozfRJ8+dASiPWDur4I+MxpMb1O0o3wYVuNGVvenVosxsnyud
f9bNZXIgq0VMaZfpcPf9BGH2PfFMrEto3OCCd59Glh511PX0AzuSnQMhjiQyvX6k
+sFoxFBLtgaJbAruGs5AuCQvSVpMYfm8/1crDQ/CNIy+Hbt9eNdhKqbZgq86O0tn
iPCAWOxOtJOMccXLYYuHGhH8VPYcBfC2tdtZwcBgCpdu9lbNnyb5qh677oT9HScA
FvYoZgbegFG/rF7yxQM9Xz0uTPjUHPGsepS2Darby3BZhqGhoZWP40sE8C3LBPuI
VwfccZf/FXrz2FrZdI5pRpSqddAovpviCnCwgcVMTNn82JcmNTBwCe/pMDOxeyBE
XDInDHv8v29CFlfyoVFMnYSnL5kvfzSY13P5U0K8ezYb5NJjiDnR15gLr5Jeaubj
Z2B18OOa7BpJ96j7UoklfYC4PzQ3MdcTFDB/pzg/BiV4mLJt+RqBbGGURSDA4F48
EhgoKBSiafgw0/+4z9KDLuW6OC6EETI4Jfz/EVJX3xVawO8RmCv2ipIMY3TashJK
K8fr3n+3RK6s64I/tVS51/m6YyqQdcSV3iXlwpfKHHeESSYPRW4KrOW2KNElETRY
gQhbdc4WbVAOn5fQlalOLE19KHMqX/ZRA4g5skFI7HeuKGVsIWp+Tw03cKkIOEma
3GfH+gRKPuMi1vWEqRtJf+p6CycAgl4EXDIktt5fKPfWvFY54NubNuJbQq5V46oi
U9GlJndvN7iDj8lb2Qx5U5UmxqQJBA3Xorb9o5Xt5A/K7vwtjEq7nRwqA8ZhP5NJ
DOQU6k9qOgLlZECfW3W7Ic2L+wLIitS2luQ7cHyv73CsGRImkYgPNZN49XrFnqwL
VWxbK5EMEdo7JYtuC82X0Un8Dfy7PpBDBlvO21ltkWV08yhsRKjJ0XHXaHfk5H9g
JESWuyBawYNWh8t0Dts1AapKNh6rMXGLA7Tcytf/eyyIf/9b2YyAPsNd8mrOPsdc
pwoySpAqHxkuf4gZ+v8ySPKccIB1KltK8NerWk9Uk9TBrNYkKAHAzd8zaxnyitgJ
M53q12lznc4bBYO+t0lhjmMqktDsY2iRYU20TnAwNqhhpHF4KdHe1ua6Y1oJBj/b
nh3Opn446mlVHTNU8l+9OB8bB5X7ILvqWBhTu9XNEsMGad4tspIsoDT2Su9xraRq
dcjdD2IjqQ3e+Z32iC186scl1TZk751LvKRWgWvXn+9vze3eC3pGC0CeNapZ5J3l
Id518KewP1SkxBR3ARqiSgy49ltGURoRXui797vt++mn7Xw+NzPiWUK1yP6jyjXh
ee3v5sfSBqeSII+P7fGyH4XjRpuMdoRE0q+D2rcWF1ZIg4ZcI6aEg+LVaeZ/V2a8
BYPlQsdPZCGi8xkg4m0Rm9lUMsNX1oPDT8Gyh5eCwzeWnIntFtcwkQ09AmHRnIir
iteXejfeNK2imFiJfZZFPRhp7jXmIXizH+lWAFjq6+fgK5LD6jYE7SAEJO6hMrsF
8O2fSot0RNK6P4DdyfIbUodYrXKcRhL4mKSQA2JV9zKYAZL8ka5QeEKkYODl1F74
iaJiOVwAOni8bmYnqDW0BgItDhPkE99QS6biFFO778w4asOY56PPQ5FiJh4KdsY/
Xko4cK6G34bOts1Ah1eqfBT1C4tSXr/zphI1dm30HsoQcovD5vGX/lC2rS0Xrhdy
siRF97dhpp0nDpcyGhWyYMReNtmRceop6fZrKy2Z8h3g+4zoDf6lBm5jan2g928B
ZzSCFaNHO054/cNJEnwPadpOnYRnGtyMa6cJNOJWdhrwjsCeJocfVVtzNDFGv/Pf
boePcIgM1Sz4zU1SPZxymVF4Skps+tze/7FC56yqX76CzDCLe7UIYIGeTEvuf6Ys
RFYkmkbB6HywTgRWP6jhSoK6D+IaMFk93x+IrOg43+hMxO3tLNZKcPnd/xu0oBhZ
DdZgj55w0X0ELI1OhKNcL8YmitBs4LOpAZw+JqLhPSEkaqavVh28SnCog6LyxIVd
OMWHXbRiv0xlBq25gZ3Mf2dIGaO/2Km9a0M5fm6CD0uIyMAsYBrKc0xSfSFLFF3N
EIH1dp+LECIhid3wet3R3cDwwIs+IpY/aTgNmUCJSc7JB1UX6foC7Hf3u1QqD/8O
yagRNOsPVfsBVEPpmY+JFsS5wv58kUgUkCB1cK+4cGN2hXPnqwUg09HlsJfDbnXe
FMib+CDrIFM8H++BDJZd0EmCO4dvc56oCAOWWwaDXvIqDufYMT/nixTtYRXydsZQ
8iOGu3CYXkAvF8KIre8EFhyAP88vJjWuWF5VWzdCPDhpy3Ip61WZMNCKPEg9RN31
m1EkyKDNAfcfsQxwOY4jLTr5JpDu069WR4ZPjxLogAiQ0mDqXow1kr1GYflBXXKC
t+MBiIAzOxRcren2dKB2bIZxcTyOsvNtDKyQYJlpHLyrlI+X6+Fm3RIaMtwqo5FJ
0N67pK6scliMopcMNDkXRrmMUhvstr+v8iP9iFfXcASQnYRkfP+vPcHCr5bRebbm
b945DcaJwmZk9WKGmeHNVOhiYlpDsD7AIJ27qJNLOuXPG05i58notZJKORhzniN2
ccdknXgVcQXruA5pXtbadzC/PAp+YtuLkpQbl6q7hxtV7A9XMCFsfXtbcw5XqhaX
WtJOITMawC8s+OA60ZZxf5H9UdJWfJEDiL3cB3LS9VEt+zEcseM8oX2J5O5qQqRY
OTMltNQzUVNoTDmIQCSd4+E9AKHKFsvY5iPRZyRoC6CDp6oIZf7+M3FmdYrbx5yb
MbambHtZc6LAvtpsXIznm3GwOT07bY5ZYsPMXulZ4dPtnWji9oSz6co39wiS/Tvc
faDFSaETyRMH52ICVXQvL10MSZ6MLu75pzVs0l/0/hfqQ13nvvwMikBhOSc48rWq
hJFzlpyTYGMfyjFBw8cW3I7BZwUXdQFdaikYmqWa2QVOC8pXqLtUFg2CFKEvql29
Scrr9P+9P8c+PNa9tEF6n07BQdxsTQCuxqL1/lrbjamSaimq4+l3Tr5SRb9kp2RK
V2V3UZmhfmLOLxaTmpQDBnwAWZW3ZBoUQQ415AqbgmIfOkusSORbsbT2ak8joNgY
zNXR8qT4DZkgj+DApLEjOz9M+RdrvB2fQNRZX4DJ9bE08IcEpE34akQqxpTept7j
R7ADakoApQZLxFpow3WWjFQjZCpCl+gbm1T9xp8WnwwezVLXnMhP/EpcMRJn6soy
CEDjSUg57ZwRDQ2EeiUmD2uR2U852ekW+vdDrwvOrZkLAXF8eai+V1sSjmwDd4Qh
sZlgj6FnRVuYT9dA+E77kMhwIYkvp86dkt2HQtxiGEIiO8dJMAZIdh1rFHxcz43I
bXbn6jutt6pDIQDo6/66BcUWasuukDHOQaFOb/Xas/4Wx85NIouz72bY0vzD22i0
CBz4GdZrnpZqb9ZDoxdL0WpMflPfokXhDli0T7L6lsBjI/02UjOXZfeP93Pn3nTf
T2/o6o1gxV5GR8jl3jTjbU/y17KC582hABCHXRN6IgX+u6oz4qoZOFoJ5MeyzHk+
Mn42HxwrN/brAepx4WuuBP7MeLD1cT0+pcVe9h8tXJpuHDrUjgwChlGW3WvcKcvP
J05Bd1Fzo6W7PmfmFsHp/gpbLCk4UpAhmDzGUN9uAi2iKjgY8HIR4voh+4JuiCRy
KHtEcg2dw7HkH/7Wt6ZdIilVPc/nXMRXZjUeKRkCZRnfrhcOhQXFmaqYgF/MPBmD
4pMVkBegk7HV3oKlO0ydN4hN8y2TeTqSoNIgYKs8JP3r/I0N0e/Fro+0AfGkxA3R
NrGXCWoWHPl3QHNmzbYyWUMNX5agp15WT4SB2hkvyuqof07Pj9r7iPF36R1xdUai
VIoKZoFcEd0/gaLY4cxf9Ha8ZQupaM/QL8rJsFxM7/rzXtvorUc4tgnYacF4AzlW
WFzRYphsdlXz8+gBw9VARlbEiEwlkuDDa53xRfEmM3otQfFptyRQuWaGTd3Bc0Om
fVu7RbhXM85JXWimstQddmKSz/j/sW/UQKBI6IPDVykSRNsTbs9HXsMlwtc5pj09
X99WYMxgbUHGgA4UR3Iopn3okWLyW/51I+0I1+j5FdpRt4i2wuRnJwHdNjlHX5vv
rDhHFXshG7kM16E7C0feVKsYkrDwudubjZpxJ6KJ9ZfDSH7+EC2OukkzVDAdZRMW
qH3To47/NAZtEyOOhgFuEk1/dRrQGj7/LVqAW+0penjNE1I0o82fRGl+Vz21ZYw+
Cz6ZTezcBUEKc7eTAbZ2jZfHePrX93dEw2fcHnjeoy/tVKRl1B7whEjwEP/xYFKB
Hm0U58pG5KetedcoTxSpnjodp17XS5rporcgXLjc8Rgf8NrkA//V+TeWtp1os8UI
iThfTEJfz8Kbl34jzGwDqV4vlozf6LuF5wVl1kHBRZwwSqf/Ie8r8X9xkv8wgOog
Lc0biWykT6w1Twdk19bzkkHwVU81qlNmXZEHsjec2yngM0PYDCHOC21YN9yjEh57
MVWSdKt4oRe/QwF9mxVfBxlQcVdldkJE/jiWUncIYuwtxJbznCCAHv7pcsguYmIi
fAHSJpPMPNYNeKuY0mOKOB3DRc8RMJhDXqMzkOia/8RbbUfg1ASkY4HWmjctyOLO
nlvvVuR23vj4d8RHWiEOk7SNBAsb8rrOFuyon3yNfrmdGjyfbpz6V66nKg9pWN4H
yD3F61SQNIYPnTwcq5NvYdVyGEzWOk+c9+PVVKphpqHvuGdK8gOz2O1OGSkADZYb
FF0upoSmZE7z1l8saaBcPJc288orekMJhbXzkAgWnGo1AEGvHlQaYxfWmMuCIgU8
wKj61D+xqUpqA1aXO0SJexS2V1ScpXkOg31DqNvvzxrbxam/fIssY+8yqnDzEdWx
Nd/uMZQSowaW2VJRKbO90pZfj+vkON+qxAeVbWvtnfdgD7YajHH2Zdm8S6hsyp78
yi8FGIGMB/ozhMaAHRrBiA5Pqjn8QxM70B8W4iw3dVF3JmSci7M0WQhoapTq1VM0
3NGBNFnCQPzBFFgaAaqK3iI3ebdDarBu8tcezycVkFZdsMCVAYh10P53WOfyU8XI
Hc9sxyojg6hUDWAgfc6YUhZj51eay1G47UztwjZmBWXl0XuBfkmxBazyPcGeuxwU
eNVOGe+zOCqBoNnNw85NheVcsC0DuuXVjkzIWSROC4LFREYLVSPe7MOM8k6sJqTM
nnvmO5D3yTAGmzylnxgBB5uELmsNgS9kFLiwRy1urUXOFGJ7kvKV7KEXx+sPoRRp
AfQxB4Gmr5VrjhYiCZtXCKBecVJSSYxi6XUzcMYMqE/gNqRLTN9+1rym416j02un
VxGmDx8K1TXlKvGRd0EX+pkL8Lbs5wR+BFybYpIF6zSNOVX1880bjQSh9Yz4Gn5V
6cU53OsMrG6EU9DsVelNp7zTakRrmT1PfJCBx9HcQ2XqGsUgu42YB3HyNfZB/UVN
4pQmn+NMxZqjnE2iIl5bZ5kYn3C1wgnjE24YOffSNgSauIL92/F635aMSIgtaurb
WrnH2eJjxVksfEExyV91m0rRlRIMUg1dthBvmFV7Ov2D71ZF3C82wyqJOWXfSJHI
NCDKGhdJj84iHTQznRfSyFUCTbz5fNuDRcyhHTXANpxMzjBT9A27+7QctpgKIOnT
mAM/ZXcHxTmABKZpd33HzA5t4u7xZ0gwG6u1Y3DwzZ5P9WonKg2vEvhN7SSCOgYM
dTiuSNZRGgtc3rN3B2vPRrxlMy3Ja4MNOSPynIlKW2HQRggnJU3MgelSoIvTn+Gq
FcQ5EyxzL9ohwojRqVWR676glmQo0mtmFfYH+MVk12ifshq8Q9cmYk4ed1qCneni
WsWyKfh8lV/4+9yZJHB7e8evMJIOhxYCbMyzRpXlVQx7QH5LRy9zgJo8WO101IF0
Vh+k6QWskxWLWFQoaajg4fiiMZuleQgt+kNsqgnSHxZPnpXRvO5zUNtFw1k2U0Fs
FeSCPtpgYyUCHZUie+SpouCwjwgr6GmF2MJWl7qM9FZknyS+uS3876JKC+30silo
5lyUmHQrrGUOB0Hb1i/oPeZBDR8Dlu1DvzWPTpDOK2my8WybAVYPCwpDjwV1S5PC
4/NQv8rbOjn2kLsu9L7uIOg/Ois4BE7sxbzx70n+v5vmSgE/MQEhg8l3JVYa3tSL
t2cDgBqzIfaV2JbhNdtJDiaYnmNxIoAUqVTJRQiFXk1FKI7AMOHhL/m1149+ZmDG
AT+PrRxyKqG4ENa4E9WOowIPxSWTA5OilesxuXa0SLTxUDkVM5szlDey0WpaVz7K
feMWrFfCUa8RGKqggH7m+rQqFEogEomYYiv4i1GCBICLqWWGK6y7RZHJU2bTtEe6
x/Cc1kghrxf0aNCFLwZvWbD2BKlH+bX914ap//oh2USlDTCwy32xzX9HHCo6DiSB
UN4ybAY9thHc95EASmKbwPmvEKW3HyVq0Z5lIEzZk0i3KwQG8ZrfO0zw3gjAXygo
JVnc2p3vRjRiA+RYRKClmZpr++/vKh50VqgdFKch64nYIJk8ImYQMsrv2fMH7/ax
VbG1Emerr2Ico5mt9fRgn/Yiqtc3NZiRuebyYFmDIK2RFcqAym+yc6t1Vp4hS/ut
T2TdwwsK6D1nPrKt12Q8wC4pGxemZpEhpGqdLpPBKOGNfbiD6v4ilbyPcJ+2QOVx
c77FI408Y81VPnDJ2CdcP23vRg6mGCBSN/n2mlhgz8ivXHL/LVrTq+LJlSWRxtGs
RsFOV0CPBBVBItNsTstIwtWMcJZJBbLYZo6dgkRlbUDRbvPzX3ZT2SfgDfveYa4o
qBJU9ICrIhVYbjpsODawv/pjc2FqhPNk7TwB6n/t1SCImDG0/fl2Bm7M9FXJeM5I
eLyo+4c0uvRffQlAtFF+jlJXPa253cU3F/VWETlGnJypfsAJAb7F2QpwpUMJhIK5
MCErz7WVTbrE2zyZsyQyGTLgQzJmlYPWUaVJOoXGKxfgHv0ALJ+iLDFbrLuqFXYC
d5ZedsLXrq9lPaBQ3NQR8tMHaHcMwYBDLdA3dPW/6dUzD2WzFdlfshh7rMOfecYG
AO4aIT110YmkIm8edOkuprT7ev3otCM5Wb+m4j+dt076Y2YpK/dVqcm8tBaX3U/L
DAzblnIdmoudfdmXMr/g0DKovOoHNKtcaLqvro7/INfTRLYr+pjze/TLPpAULUiR
I6bVFtPdcGe4oVx38nxpgWCFJQXVtIjcoli8RDqDnLSdN94WTm2RuG0ihRd446b2
K6oXYDTLMfGSElSUi6p9yqP1v5Ac/+G+HMlsyclagvhPNLZk2ukPMJpHtp98CtVZ
9ShS8bpNj7pQPFM8PPPnRagRfWggLvKKELc+cGsQ7kvPCe7XFe45sf18+c4u2yjf
wOSR73k+yEvuUn/xspcUMAnx10ZC9lgHaPizy61JsRVXw9Oo9ZxwBty86z568ApD
orC5tlYXSIR7BfuKeG52tpZrWGYujY2jL1t28b0Pqm9+GapkpgfMx6Csd/NpB744
wWFn0GxuYIkJVCxJomgO95pJL0o2fB7cR7bDHwu9gloArjk95vdzZcsoz7/V2OBH
V8TO/UZ+GE+W1/0g8CIbpGC0TnBAXM7fOzyU7ReyBAe6L8IkPbKGNfv5JbkXJ4JF
bRtvfbbZ2dqSWNYasf4jHyUth7uvyxbH0l7n9licSheWkb65bsgZazxL3sYJ9b87
UYU36sGoFCajV8eaLHLV7IKVpmOsdeGA9LXF8f6jguze9Eiqo2rxroTr8XQAghsV
1VorKmDbSHvQwJCDa5u3gkgP2k4r8a234cWJrnivBq3LqyA6zO6zEQcxbXgnWmtj
Egz4oX4fmV+pLj6zVnO+qhLmvwRwoje2oF1R+1hC2Z08uFcrLlzBF7sco/VYcaxS
Nk3ljz1DXBYuYEyEAGGMpcInQyif0VRQHVmKpxZ3ZwyegTOH3lzx3yzW2KxY4k+s
InkNfefURSgWyDfzqYZhlQfU0MyOWUhI7g4ozogPkEyEieQsq7CP93C6UB20M2oX
Opvr2R/xH4896DwcuDUaSShGjMcrZQ0NnwfCnCtjzG8IfqAY5CC9xqCqNp23Mh6V
JQ91hPQA0+N0mtnPOHMyEgmCwgNYx1SEsbvxVUte4OKsAY4/N0jFtKWm8RWOkSt0
RrxsynsjYVDKwHxyizHLQAAeIi7WjwYFrNXy0qBNzmDqv+iZuCrbv1GbCk0BGyH0
OK474LRtcP9FYbgKrs1tubTOClQH+Du1xVWcl4ggVj3/1GV1mvp2AAp7moD2yUnb
MPwlZKT2vJ0VsqyTJEXrZybn1xzxYbpXvAta7nhBBSSyuwBvzzJz5bQicBqj3wxx
UnNduH3bA+ESGFv8TQYZPXSICwW6XrkOoZs8Si07qIy6xYgPR+gBAzOcTp8QxATY
DXRW7aJPohn/OZSp2lpqABAVSj+iDJksYPXze0cYCsXuItwWFF4Xv2E8CpQo/SlC
Yv/KOVRNqA4NgatJJdiU1Rmf9y9WeQzqEL+T77SFdiLWjHYVZzhzOrthem7R0xyL
Acuq0nkITTsF60BdcI/p1aRcgMja0OgXg0WIq/bhCO4kZXJEa5m8WdHgZFsjdbLt
qMS4SI8F2+kouLEQ8hhnVwbRytGnuP40X4wB2gzTwE5G4Ms5TFr4nK5ymu/abEOa
kzH92Q2Vaghbw+iRtT2AzF5w+SIl4L+Aoz2/JxL5+42ZUrYBGBz6i6PWQvb6HF1o
yQPIfq7mvKfhowkkfNjvzY+/CpmT8T09ylbk60pM9mprBeDty6HA2XmaNo2r/32/
IC6JFwMqc1a083OFArk6rS7vkkfC7eGQ7LsnIXGi3nXuNw2ROkxBKGPuIQnrDpE8
RRh4rVcxijhVsZ0+5RofKP91FZanFUW2xa9JADE5/BY3GbdQy8D51SFzoDanMXKn
491qxXaTFCraLqebxYi0vv9P3ySo+C2NDFHsQCFNxLC5o7AUHWEBUTfqHQ132qki
2BTOs9MQf8qhu/y2m1g8Kdox34q77U4ZJLL8rEPOInQKznLwrcxvqnxzFPpjsK33
Ymr3beKKdeDKwcUF6bZXij3iZt7fbR8VQyEz0PO/js+uyPHBN2QxzsP9gwyAzkf3
v7JpVT/DrIuReSYLgymJFC0YRsZSukqfhQPMIuXPY/5/p9D8xAwYrEEn3/h5EU9+
y9CxMNJHk1WDnQhdIswvagspVtkTLdJCseWiv2l96LMEXQIosfZmv5b220eYwILV
M4zv3aWHKA5M5vJuQcRWzeNf8NTvqZXOboYWgKbzi5ysBgA8VxoYMQBHVgEAqk9l
KS9mc+fEXwgEemg2Tr+oGfOH+C5fgKbeoCAI6lcbrPLjqWyO/H8mmzwz1n8Sa0wP
E5G12zFgipuWvW0jTNiHVJXEeFLgKhSXRaaNtZapWz1Dre5/mWbYpXQ/plb5Y9Yq
pj/wEQhR0P1uOtG/qXKMK2KOdclROlCFfLNLsfkzh7ioI8UrbQNu+uY4Bz9L/FB+
RbPM3eyIE4Tu96xvrPEwovAINiw9eAAfE5TlUcRU37bdAbNwpfBMIL1lnJT/UD9S
4WiF1aASI8HJF/1d2Pl94f8HNbZCt6GNRdGm+iSKZiZriU/WfxZt73FL2NRUDsFv
/rjrB0IZeJWjp7KjN02YTUjlq4HIbbGbeqATxDlpvBTTmYtiK5nOrmFEdBlhY2TK
LpJUBFKa1VXFp6fmzM+tDoHc1lI1YhIcoT9W4k/ikg+3LczaYSWXeZdAtmTx7vSf
9vnO9BCT/fNIYyhoKADD3JDq9T/fF5KP9P3NeqJ5TPHOjsrPKaJsqCaWV1/3aW0C
pI79/7cl4Tl6gSXcgEsQo5joYmI4WCG8TBbN+eQoYiIly17Yoxo4cV06quRaW03U
A4R9ARPRF7ZFCLitpYu6PPpwOY6Qk1amFi2jMaP/YgRwO7m9jU1bWC/aZCHE+/w9
8b00de0i418bg8CEFV9SbZNvnO/Su0zA5feDdMUcZg0V0CfGT4zdEoLMc44+d2lg
K5VxGTbNvf49LcyCgjxhytnUmlXAIeY0hM9lnCAIgNDlrBBe4wlIsSFpNb+midpO
FACV0Kz3EKHa72otSlyaE0PkEfBh/g2nrwG+Fhq8wYi+T+By/XPRFTqpZQyf51VU
rv1dKQ3lvyew+Jd3h0kPj9s4CtKxp2GwYYGP8qDLWoZJccyHC94GVtX6IPs+mWiw
WXdLdkami800jhk9glLDW4q/dvuXLb+9Qoo3Ei+OUnAZSVhm2guOCd4YXNFDw0No
YoRv7jLKKTyfsauw8LVwONVxludO11GxHU4b6BJb+xE91/+XuDxh/cjsybr0rs0j
wMVMurqUh366Epp542re8j/otYSpvTkUDU1sW2dv5InnWoXmx94RccfaEKBhGpqI
p/7Ry9CAH/kFcEPFRqDXMq5fxCS/YnjHh4QLTW7i7IUf5KxlPQrfYInWPP34u4F5
GVL40GqKP1Dw/X4Oxm6Qv73ub94Ic4kVw171Drr5lWv0ed4GmvribLVbWK17gMr0
Nil8txyK4hBHmFeTMDUHkgLP20I9FMHWCoCmw4aGekt2Mn2GLnGvWY16o2OhmuF4
uxyhFDyOsfp/bn6qsQMgb+jfp0/is0bjhIsPxh6wqGL/Jo10sESw5nPCLyCfCi9u
8hx+fDR04rK17b52SewPPD/ohccB4CL2lw6C2VnckpKDycsWDzJgxxmQIDwqmZUr
lqUZst0mpezlLMg744ZPDnqcMyVQUoPSaSzgUyV6yp0PBQv9C0Ooj033ioJe1/b8
6il5NGev4KfiOk7/xpfCsZjdWtdMu7XtuE/cTox4tDu97ReiNwwSwJg7I/gxFZ7v
cwr1xRMjAa6lhJKU1Fpul2XJKl0RwuqtX4cvCgKQaJyA5P8uaEkxc0T6aix8Bg7+
7BdjgVo+9vN49+mF5TvmKpZI1Dyo4zNRYmVC0pO4HUsDfFrWG3BsCT47Zxb20FHK
IjRE+7M7IdU3D7ycAvm3/TOCyH8vgmsBQ3hhrE2/A/gVBJkDVRXWvwojHJRlturF
ofNCVtVYFps49Bz8Kv0K5ChD79ByOt55LTW1O+1hAToOa2arQQ4Yj6EeYgGknN8X
gWVFSVbENBMfXGX6PaIBJVxPWoxDx9M9NJJRlWyk3jW0jV3krWRgzo9700Kftxi8
pc0o1Ta4Szj2a2FUH4UX5BugBMonmHyj3CeLkRI+XJcWRScoxZh57eIwl0/QleMn
x0HaSBJLAVRc1aWXcUkQBwg/Qyf6KX70AKCnfNPuf257wGP6SItgqmJG1c3vT5eD
gAfdZzgC/qhUwi0W/SKjik2GwWQyGvd+bI+HyvVFfHJ3U6QBvRdOHAxe2SC/zFsp
Hg9ioKcWhx1DsmZ50aOV7twh5Hz1D4EMkyFgHwLOKypQZcdS4lnyLqYXCk9cUBDt
yzhUc/jj7aAu188i48vPCzipXb86y20eZplJmMzkunXUfw6dByTFRwKIOJbS+ZVr
gm/BXGhMrdgUSSICmFqiEijE00QR0nQ3SiliPeeN9NLIIOni+vK4lySYeUKSFsCE
mmdKr87I+6I3kYqe++OpM+0b+RdovYBAS8qhhVqS5fPrKB2fyd9LlBC5+6WGoVWn
IO6Fi5GfIlnLLeFJKZDcdP1Hk70O8Dl0L2H66vI5uLIbIldPdkku9C/3rNo6AaRo
Wd0Z4cD2i6oyFusof+5aE53i+xYqnYTp02iDmysxiDpTH6MPWBBptyua9m7q1Zzp
1MjpqH8tc560EdcJJCCHMvYVpYmAU76usIwW8Sg0jjLN1kWJRYRw2FsoH05IZTqL
3mYaetfbjACFiWpf1pZvxAqJheWSEa3NC2+yKq1+bGVsaakED35njW4N6VP7mMBQ
pegC4xqUu5+OftMoiU/ydfVqV4TBxWkSJ20k6zOLVVGCsEYTuBNjiyXtEyBINEtC
2XkhPax4ztmC2n2oMhk1nJ6XFoD+hIZopvJvW6K7WsE1m419Tcql8bLPEZF1gNsX
At0Vyjd17NXRzW9s+7X94QU4QHRD1NqSVW0yZaPoXGfnwqQtGhXASsKkR1cbQiiD
L7sYDF0nYykizJIoJvC73/rdCWOERAqcmTKwfflaWax/eWkaQz3zx5el2TllsCBW
SLW1Iey8mmtaUPPAFJUioPZIbbk6vvlvaVZl08VhXjOyCO8R4mALPPZpsX38CZ12
HbyP5r6GisSIzE+17e43GTtNdR+KZyEClQOOcPsMYx+kMvN0vEf/tTU8MdEPqVE7
ac3lcpf/WqJ7kYkyGCnNK2dPCTS/14RbtFTn9ex0jLPbeArzNbVLFlG5FXTDHbhI
5u26up3ezKj2QFsUSt6rEwH7ozZQaGJSeg5hbELmw5TQ2vUQHA/qauVWXtY3XkpV
Pb22IXa/GIsB1VGrnXMT0Sg2LxqxB8Wbg057HPccoYhThso2PmiFp45ymcfJWoQG
OOLQa2C07OPk3W4ZkvCKoB9yFGkdnDPH8hBA2eV30oZvUkhGXer4acb0WvSxw6Q7
O+DyI1D6k1SQWFMswkQPM6cEkT0rI9vHyZxZ9PeCv/Fgv3bkzdNeic8kEJF0O8GU
FDzsmsmDhMbKG7wK5wlNlsq0ejmSdXZ1U5K33KoVrgQrA1G1joQFe72T+uyZteMQ
SRiGO4v3rz6kUBfsBzAAg0w6wGQDaSIrn3GEC7N6DhOupqPZk3IUcYd4i+eDhANC
aJnhG7jjTJe2i8jJU7hgSyf87SPIdHaZW68O0PErXIrLG8AQhfmvRqc/55YMkeXA
F063dbPFGgmGqa/nLJNl3fyVrUX0or128VOPKb1ApOM1lGImCw7FCX/Mmyhjk1Af
vLu4bjNw84NSnU5aVuS8SdlLR7JSGO2KmwxJEuwo4IP8kj47Eqs+NuOkc0wawj0X
4uiIuXv5F9rjp2wZWJl+Ch68y2/uSgEQPJAtyiDQ8tZkWWuFnAAae1ea2rKVRr26
1/hk0jVB8GPLsWOIOSrxMXu9f1RQIF9fLwbna1BiSe4X330GwkePxZtgbJbB8MNH
o4TmtZ6xD7aINo5RZRq1vxSXYfgLC18u5D3NLHpP18iD/MUafbZWaGG5N7ug6AXy
MAcLisupXefezHWIbfnZYuTZhgIzui0+G5peDMIQK2aeyUtSzWImJWv0gSSbAVZH
xbBKiGNhwNxz/l/yl1eer0juF5vpS74O+JY9FfND8TxYDtcZ93qdvja8sFdKZ1Lo
xiujyUu6RBRHhFiyPIa5HAgcUQYy941TVExtEbE00/08iTO4xbAzLxZWH2OX4mPm
rCoeVbPvynGba4lu5sM6/gO/wQ0WqBhfAC/BsmvSjGDoM4uoZW0tAqHdC8ejrXlp
u0uGgPwXPzA7B1LYsJnn5ynvbbNx4akyFktlA3HtiC4B356KSar+DYJTwFJK4Hyf
Nmdp4e/zxGitzcdIiDWqmeHFzVSlsmAq4zrkUjr5L6vm6lHJ7sTzy6OXRrfIULlz
ykmDb8mugyvdgqRrx+fle8k3etHFVzOKWDeXuQga+nE3utOTWYH6m2jPPDSFbJ2c
iXlIGMnxdAdzDrOQf5F2gYc3hELsnROxpzy+s6igoACtnkAcqwfihzzYlGx44+Gp
DE9M9rrnNHDQab2M9hNzKKfSC8HRuw+3K9T0cb6kxJKeBiz9W7EqkRqGjUutYAa1
ulupWELVV8uUB13lHOdTkuMCbl2XUf2NSDQGmRg1l1AQktTmzMvic8YXtQg8oNAL
7Wrt1YVKie/alE0aA1kLwY2Ifg6X6+alrDj++dCvTfQtWx2Ri1XH7Ogm24rMe9ZD
ky4ihSA2eYV6y4e4c36WbPAcnyWaLMAmP4d3/+hhup7xV6ABZFsL8aGy9utCzyc1
ZzqOSJfI6EOxSiqkrypTMd7iUjMY8A9iSYkvK0V70eKEHDjaZBUEzK0mwxVeotvT
TEwiyoFJkm9qP3YEAsdWcUqwkKsP/Xev6A9x9+yjQijgyCKA1cAJC6XbGeCDXG3D
UeWFs2Vz+1ympgelVMadIpMI7jGkqseof7XWOv7lOF3fDfBja8P66PHrnK09cVkK
NttnJhN5F7ZBRIh7v/EENaVbYA83Hz9H26761U5/IKtDAbmkJZyQgb01juQYddLs
xtdi/BT6SfJex7tCBGg6D1qLMVZT8MpLmoE3ATtXndcaZRUy52cyqvVDlLTM7cIk
ZOaTWRexHSNza/SZEsWzxwN30xijHd01ihe157mW601iKkHGpDLeSSDuu0GIFd6k
UEFhS0ZgyvSYvOQE5WJG7gjW911FAYKVwfi1xhq7dCNk4p6j6w5A+yWNgt6jGh1b
EEhPw7OUxwdCEAzUyzwt2XdzUYGKmbYmCVfXWgG3+M+DxlCfCmZqVsxD+uAGxar2
ZW8zUGQjTFteWjoFZD6EVyc1VYhS+bdHDxdkNomOH8YRQDB+pvaXhzU77QEM2/Fy
VAh4Q/434HG5FkSVIGMcVQ6s+OP+rqtQPtu+w9vjIaX3ILiHouRhgIRuKjFt+xoB
baaeUmTTWvi7Iw/d2YQJ3ElyV+qgO8L/IrV6sraKW8z2dnDmskaRCxFzbFqRMc75
+8a8RGLFG3m3WMfOyIS6S4wecQkWsH4duT10UOwLe8mbWS0ttHt6T4onunWZFzCf
2WJy96K11Hx8KAkAd7O3o4XHZKInHst8dYRw8J3dKqfdQQqT3+FA2/ROumJoWzgA
mSBcr6gKpso/9QnZ5cHNyJueaEAeWF0tV4ICgJcxhvjLBiJAQU3zCYe0pk+MFM7J
t277GosfaoRYzMGk3GLxq9u5EDcLtfSfMCm8UHmG2efixLASgfZ8Gt03hvFUIP3Z
koO7Y3M9zagXiA8kYa5wmKOKIsltY6NCzG+pv5LlcXPhbyffZF1btcCMhUG6d7C3
3prCVPSTxhbDurWymwMj3l0TeKJyZhtNuXM0GBI5VAzLfIWJr8PV5WOA7pdVnh9G
b9g0QZ7cPFjUth6m/e5xksQ1CZfAQMHJYwftbyRLhgvrt+ENpACgTjohp5fnDSL7
HSLx4Sn5uZBFXim5b4Jgm+fwN9pG29DPLPmXPHlQBJz6kQ28+6k/UqyjXGDw67Xw
U7sW/w5uyE+BkmspVxMroN+AgOiUsp+e2W0Ib6sliRK2UHiHs05farq817e1XVTx
45x5HPIGhD/zShCBC7Q7nToE3+FMNar9ZOwJsqVnW/lyBNnuCRynrnSvd1p1xiKA
Etc2jQij4fnvz6w/Pe/UIi6XmXeCmVt73T7CotkXu2Hx2lOyWPTd/qg04C6Rb+Gg
TaB8xzlJKhijl+qjk/IwSGntPiGoCeqR+eRn4GsBMhKV8MGa2e6RCczYzK7qbbxY
SmAzWdk6un8YK9MMhpW3SE/K2OOFmXhkaREyKYrIaawanP8TlGgMqUQVSz2EWjve
CzsWCtuNFqOItXcPraJUEsRu7Aj5Oy7xf04yKd5KEbfbD2J0fVrFLq1Oqp0koyms
LaKAk5AmOvmmWTFidylZswO5/QUfDP2Pw7Ohx85uJYy4hyN4zK993kamV4hr77hB
etkgifTab4tg0+U2HJK6kTIt8brcPPucbohu+I9s2QQumX0G1huueEqoDGam8Cpv
CQjaU+YxPFZHxMaemuqZ5llxYQg5yh+tG681XOuOZ0w4r6KAytNkCtkO/rJpghdp
QGN+MlxB0jLWXMIV1YJUGfXe4Sn5UmbCDT/IhdIZVVWwKaiVYNMCXLyuKVoe2t/L
kCNz2wTqtXmw52n3YMa1ba8PB1j6la6K86xXm7H8T6wjtTuiz+WdFhaJUaBu2j5Q
7VXJ7jiGgjxCTu9HJJl3q4q7dJiXE/xeqKcGE69lcFz9t4M6rNscLe2cnJqkMBSG
z+QouTOlTmMBydGLHmG13jsoehtuwlgYtV0XYcLfhoHCKl8864bQ7OtmWhFsXm2t
IHS5wakz0AqCjvw5STd0ON4DCyFlDibx3+4LSncRQk9IM+CdvsrtCqd6nzKLvv+G
2nwUGSEK8vJrZ3OVtvduabtE6PGYd2WozmN6LsVBbFN0dmDyMQBkKxTeVr6mEqh6
tFuFXdd4Z24navDuklSg+nuzcaKK4+Dt8t5ovBLjklXH9I8SBKInIv1VURGoRQjx
P9tm8IFGv+oC1Rq1az/+w4HkcCg1KlWPmhclVrh/sTJm/hml+cY++lJsSyqrbhK7
FGv+V0AVua8zTt4xm/9X1bKADI/Uwxs1FzBEqhrJuvAZ/i/R2OgdkSOcEBI5n02q
NmVz8+fecqTNmcKOYE1Wcxp12RteYURet9Dmk78jg8fjPlNS+4NmHJdYcBL3ykzN
iCjD79Kv4hPQnGghQj+ZZdswGDvHseZhf60cJ48anGpcvWfoQc0kScQydLJnRL/5
LYLEZdzWfi3oky430xnruKLNPgZhGr8Ne+HCSm5hlp4qy3fwtz1Iuy59kOv4Ex/S
hu0782Pqz22v9se0uGXDLDVH4ZYdPiNmHUYrh2beVjMJyunLc3JwY+Txrw0PTSO4
gHDLvjqBHZR8XnDb1ImaO+isgqMkBt+DiQh+kpRU0+fSPhAGWRECfWBaZQvCh6sd
moKA44L7YIhH37JdGuMv7YJj9yuCm8W4EnWMbBnYEKXpA6HXc7Ak1pspLA+J7b9A
kP7gEIjZHNPRY6tGIF9SgB6xFSv00xfzTzGjOjRgJGonoFECJisGD17Y0RCdqFxl
K67E+rNT/Uqda8Na+zfE0sVOXBTQ+KJ61lRVxS0ZCVYLBvZxZTNTZ86CrsCRChfR
jNUku/4sXgfOo16+8htdjwhEPyENRBqy6Deg8C6zU8U4z5rEbaE31lenGWgJ6H+B
C9hqHkrwos6j33VimO+FSX5F4/g8FjtbfTh8xt5FGPtrXcET899sJZb19zR57ZVm
ikkK/FuGmsY5/PF/pfIUwtJAKCKc05CoUDwjSaT+t/cUus7+2A/cBCsdtSus+vNv
k6YCtQt2xfzYo9ozLHBICtsfsag41jw/1gl3L0Rz6L1cYQQrbJi7Grf6obHphjus
+PcUE0Y8YXXKbLdDT746IelgVMGO4cS8nAAHgz5Q4IXI+sD2hZRBOstjBlebjfCi
xQMSSHNZTxus1uSPbGLiFWJ3NFlCdzxO3zxGdlXFr5O5jRoAFlWKyxKvXuprRZjZ
yvGbItR0xfTX0Q1lREYANcqikwykAIihYIvgmXMACzq4rCb4P0FwBPKmpKHWNCLI
dCUlFlkH79cct83MuR/6izLmpMOJnRcoyf3Zi4Dbf77bMyYdwd5lHeda2zXZuazu
y8/cITcvZJ4M1dd4rpn7GVGiZzu7xhZrTMWdvMGfoSI7Cg0pr5BIhoww3fOyW8bP
6yC+lvkCPJ1M+NVSmmuo+AqXK/Sqf7nVQqXQARQQlstE3E4GkaHHMBO/lKyO8dkw
n07gD154lZNfrfKXlkoo8zvp6xALF4N/wt/uW1GK5FbTphn2zhFKSuTFLTvMuCft
HDwXgR4dA70P+unjsfk6Q2LoOQMLWVm/IT3D5V0xXA3rXzM7xti1ziiR0VppFjeQ
vc33sGdN0h5Cnz9IndomxOipcqirtLEPX8C+8oYt/BAMJjd4A0fLoG2UAjWurg4m
AGq/rDD622YsPFaWrMPU06iyodE0H/wjQNC0e+lvfVOoHlknXbStmzOqIwlorWAz
EogYT9b4zqi1JYaVW5e4+OojW6eQZDAd4/FV7Su4FJoZuJSaVTumq9dPFqkwWIDB
EOcZxndAXVCgM5FuH5ULbZDOXDSOrxZqPXbHTipNlSOjyinqAXGu7lDySe/1HV75
n7v/MNY4A5cST2culpgTuEvK8/30VPRle9XFKzxhka2/ELlwH9zZIbcxnCgZUR9s
0knk3l1EXKHX1C3iPvrEOMTEKsZu5vc9k9YxxB0TEp0TD8YGKuHnJDZFwr6KgDPb
oaGsgdgm6kxz+bzwyOtEpuksIlO0sN+tCaEGn9nT3y9Eo6VjWKA3glU19nxYGfD+
KFtd3wmekZDbSgu+7V/5mnoLAXLWfyBDphohLU761kULfRh419A3hZ/DL1Y7T57p
/hiITbY6mCIZWeZqj/X0zrI+xoqcHkNtn6t/LLhZLCSn3yb1QOSB3z/rUn2C7344
9ffiybXjnaDAjzNl+IoTiWZmLXQQ8SfBo+nLJ47zC49Wmtn3RUlijVmT++ds4Nhh
NbzO3lCOo72wGrmBgONgr2MU8Qj/6460UUOq+3Pv0F/KgYWPFejvJ2fOu+J6suZ+
/6ONKPp4P0amkzlOh14r9yfMS6bWEV6P6etTQiBdHVSasHLSg7ipoApG6Wn38gh+
XgJlcOL3tgsOlqFxkOzGTWwZFH0S6WHHsf9SU2LNC0vCEUijmzMz4V/5Fp+68/ju
1jD6oC91JRPTTnPOR57cZwKhrJBbrVbfTrb8lPU6TABAq81yVahY7hoBLCzsoLXy
/fOQ0dSG+MdRlUzBBehrJkSMk2ONlVm7aNIckSOxIUsdKsynFFV+AZ6ZxKC+NaA/
g9YMO4I31+V4FK30yIpOPNbCATkEx+hf44wYU82Y53/wObI8GteeZbn9oAv/1ibN
DX8n5ubFmvabvmFg62Fyv5nOns0hW+kbwviOiTtCcz3PE4eHdTqPU7FwzfRIdAWp
GV6eun/NBXMufpdgvUvBpsYertPaoU7yiOH8dQIcD1pGaUW6ZOK71+xOigIuAXVp
uCqKVUZKpmJ//6aqAA7wApJTW8hUvM5FUHryRxJlr1M6zDoovh/w88K693P0ebKP
vO/s/tfaw7cUAIs7hO6Uu4PN7FE5Okp3NRw0WxPvJ0JtT8T3DlovkhRQcZSEANTE
3tMeT9NrN86wjapN5c8GSbj3+JnkcUWITL9xJKCB3H30Fm+d7+wGdrTMPppyYzf2
zxl9spvbFClszD4a/lHxuy649wb86OAK2dpcSpKpC4X79kEaNsJENHShYQ2mMJsS
RiZTOGxBhN2rs5mgR3kLRCIbaqLqCv1wgTwjyvzFaEGy+Apo6A4ZUIUVEuxAi1EA
A+eEqUkbnpsWnpC4q+8ltlI+/DIOLZ18E+XuG2P96RSqaRUKqOj5ClzyufwBHSix
qSND1DMYcaBNSwAJ0ig6R9neAb5aWjlKAvzxUeSiBb1JTEdqTcI5scHqdP3frhe0
24q9kddzUqvdrSP0u338s8m7M+nBCMcfTSmZOK8sfd5I8+N7mKKb0lXdqzplTFmF
saSgx1mjNnwBhTz1nYspXOFwctYO7meVLhz6SKxANeSN3BAbsbkbEqneWjMpVcu+
BeAQsBAlIMJ9bH0p9ZOFEdEHuzBQb6ERIdcCjDGYiC0fMU9Qd3OuGmq+KzK4tseX
chT0tIUNrgIMn/0VBt1Z5O2asSOO3tCok53xHUTkfT9x/No27ReMFx92C5u8hv2c
9Xa0KaRJBCERJqbD/sehQc5Fc/TKycOGXWsEUJ2oGUmANn3Ouklgse1t/sG1kZHc
tLNOf6nnn175C1NaHG9ZMwZ7v8khMTrafD7DqNmskStHlcrIMIV3lhbEqMylVk7f
Xc0V7w4LvtrkgGMrdSmYel3Uw8HhmkI7wSAdxSzruVsyCqpFYAFxO+OTerJ1/zpe
PPlu8rapVvsmxqc+RiVysC8mevA4g+mYSkckxv8k1qGQfTYJBylPmNeTVxcFJ4Hj
EBa/VxHFzVDUBANxFsAZEF6Mk8zCTMEuRUV7rBYVENcMv91YYlLLaTGcj+STTZvq
JD+hesflNBJBnlhlKepFPgUTa9Ind6uZ9Odru6pVUPhfoPPb7LKk3v3YEvIlJmxi
euzb9DuJv3aNVp1zYRthvQhJpT8UTtKFto7bTw480wHpwea/3il1J+HxrBA277Yk
WOtTtpmVB9iR1ahUSv1q9YnJigRkPNjrjyALaRD0qXdIpZVb1OE4M6gzYvcK7mQJ
JJsEPYxcBUHtefhw/YPe+Bn97e086RvYmmbJwVh/LwUTdaxheJaBNUxMKlz0tUPL
rqgRnP+hfPRy3Qu4DQI75C4b+RZ3PhAoZ9PittdBg7yk+UYWzTeqNhNviVXe2L7r
0VduFMQvCzRfzoywE6HcFRX0ae8jiz6VJ1BfhLTMrzCrZmFe+wn0mSEmmvWN5WjB
Iyct5rxiXv6YE22Su207Uw1aMMUhM2RNPxWFoxbFIOqHF2emhY0wWtQRj/U7MSUo
35vtIIf5AssrAcG/0Sb7dSPfXepxrD5JzSOB8VHpBSyyFVt567VDPfCd61tu1c/U
kIukmP3xfEHC/sH60eDFQkQO96z9RDuDlnDZV4T2OTbc6RF6K4/F3NWURHAHAo4K
weceIAsOGTYTZ9BFq+3Hc0tkVb1168K498lUhbJ/bTcq/x5rxNcvvPfUqPlp9EC+
V0+9ryLA49IUi2FtUhGr8HrMMsGXG6k+9wS2LW7V5tYa9EwYRv4izBLaOs4KJFh0
bZdOdE7eB3Pz+ZwECEjOF5pnw8ELYsnu/5FbJexgjssIPUR9FVjQYNBuZz2PTjP9
DD4PyTdqrPC8pC/s0Tz58l2y4ymwpeGbfeZkNbpWGnGQM7uB1S7oLghmLEC+YNkd
CED/WIjgVFo4Qs8mQS2+MyjjsjI5/032IvzsjtFVzl7Ja2vQqCdtyd5XR4SV5v9d
3TMvENy1VwD77r1R5rDl6zrFEp0uSxNko7/X5H7r7iy1EZxGD5YMZx8obEP9Q11h
QpFO6g+V8n48bo02a4ur3YgaAVIht0XB8LWXXXkcDnAHGdP5sPEG/uDhjH2hnT7O
NtZkfffICIRoVSoH0YBLEGuc3Xi8JIDiz5yp9fHpBunJ/FHMcFn4pgRiXV2Zm1TT
Ndt8tqoQy1vkX7E9/LDkse2r9drWU/IsZWKCGxxTsVbjpNMtD9aJkBedxH87ss1L
zwmsCIA1P4S6yezysK//5kr8FkNLS9MoldheGoOUiwcPriZBINJevx5uHpIbT96v
LguGcak3+RZ2TRwilFEUa0O+cE96zOxh92AcC1Pdwo51aUlGnJaK8Uq4Fob5XMbS
fJLpWp+uDybk8Oqzfz4euCptezrVuwOBfuV5RIt1/6nUvR8/6I4svUv4MhoskeWs
vTjxWa3y9ASRMIHO8kRrlN20cMiUJu0hgXIxwJQGZwtqapLQNkxNUF1yl2yU0uUi
ogjvrW5KUVB0bcBa9z9VXE/NsuE4+0W77uLlYraSGVUR0YdHVvZJVQhgm0F/r8ll
gZ/n7QbkYkouoCS3+W/fvT1jvES9Lc+20frPD3DdIYY9c0S52G38RFl8u2bSNdD7
QORtNDHp3oELswzGKSiIzoEf531t8Henyg3GdmWfBL0bQ9AgGH5oiyGNt5yaAIxN
taoiJAYppXrn6H2JWtoTzhdJVr8LtXIGw+xMD4WsrxEpGALWDYREpcNmTY74n/xz
PtYVlEFUwQSd7pSv9y2pmwTer32TD0/bN1A4MqP4eIf2LwrLrJxU/2NAxj1e2RGe
pWiDBcPPUTAfHTh0P/Iizr9L23/RjjwlZo3Nhd3yI562CjcqriP+WT+LnBVetaaz
ZFH5PN+gtKQf+l9ym4b58/53KzKiV+XPgXL8Cf5Mu+R82e9igAaGuWcw3T8OqHoi
wbEw9QfFPyWlHWTYhj3Uyyph2zUhtUEdzdGek3xp9/N2FbUXO0LGStD5/GZHcv3j
R+TWrH5kYFNYL9XxBXfYAQ34iebUGHtJo1VuTkVzVSHgh4lbBV8r9gNWuH7npwOk
F9geGw9RGYGqGgCsK03f5PkctyV+Km0YvFqHaBF3Dhvv9VbnIxNsYmmM7MiGOUma
za+MYCG2xPl8DSydmJFHBFujlFrRU8m9qjd1RZfOGT0P8VbDa2hg9kPV05N6B/B6
bs0d8jKcoTO9FlB7jJw6DdbgbYu05d5gjK/hh7vs+DKTAjoVjDoMs7H2GZI7C5X7
L0ugDm9ASjIkEk517fGnHY8nZ4HKb80sDViTlCiOy2gHlVz0Kx+Vq9lhokS3ZXMI
JvbPQ7X6elvJFd8ZSW/zGszT8RIbaiHyDQalJ/TRojVqKd3PpdbieiYxw+DzeBYX
se1RVfDcaKyFWGTAFXe/q1+O0+PtxAJ2NWpCIgPaoonpRVpZvNMbKnBuNmlx9o6z
buZnY92TjJe8amr0tHgV4osCgpeFIqLDmyxFTKN6wo2mj+or6lOS+IAIvQHuHdLK
IS1Jgm8CrMh5OhB+mof661C9oAQQFhA4K8+3naplUVI/W9M47qD4Hq7ZKIwfUOKT
UJ7PN5rexoEA2jD7d1oxQ0AqGjopmCXuvEmKvqW3SUouQjSXinisVoA1vW8o+fLn
gdpQj85EQhkJIXW0Vxt/85Aao3hKHPxyYQ1yNgPw98aUeV4LK+0MoHhutLury+LO
gO72QJteaMhNtLWaVHIbk6CMiy+r+ikZbU+DL9E/OUZ/2QR4+loRDUXogbGlgE6S
Zj1g08VZznV3/SjIpgMhuqlYYH7djdJi+UDi+ZBW8XVvl+ZOlZ81CHmWqV+EikTv
gq2bpO6yZLj57g/Zg2ngVG5Ve863/CKNkYkOxtcVbqNt+8KypQt0UAKmm+fH/FVu
DP+H4OLmTFep9mDVf28qURUuCVjLOC+588PxsoTJSqiqULnL+nFvJHgY6geOciTS
iN2lIHInrngqegbOlihg1HK2hXWhiaizy+2Z0VlB6r/bcovcP5KxMN2hVmDtDL/Y
C4N+gTqYoPj6Nrg5BOLLAgLzijcu5UyVAAix4dU2sxeeG6iNSqU1NVYjfsMK9ieY
fPjpndWUxHzLbEMICqgecBA6XdZm+b2eu/nq9ADXYTzcYCTYDTTR49jmmD6N5ATn
1J8J6aRE48oDWvuS9t9Z2ubG6OKRtu+24/pnhfL7rFSQMaDnBCCAwf7L0r+xG5K9
HYsf1mDovWT2jds8YNuiRbIEYDj6Oo6cB1oxRfw7FBmVwq0r/JLlFs6qAeAAQ+JJ
erd3/xbtYeLCeC2qJRRdz5qA182hvdwR0vSmnU+S3DuZI6MakQutNmhm1qGNRfd8
rIcOuro1jvjX1i342kVk0c54h/qtuEbqL2wxEt09Rn8wVol8lPq6xHUe7PXx7bxX
Z+DE7wrlXJ2t0aYJVI5pNZL5zTQs+Bi89yvarK7Tabp8664tTx/dEQ2L1WuOxnZW
60vRsTc1rr9gyse+dQ6IgKS2+McI7tVSEW9kS0RrLE6UTDBeQDzujX988ASNvSPu
1P1sLpxWgWvW9icVszyCV9W1zuj5xdA4Ch5eHcOKrlRRF9F22z4on6lsqi6BFdvG
MOTsvX5AxGNpp6RbqAi9sT17MOkK+CqkmN4v03CF1f7/eCxcFti618ZjmtjAVwie
Gt7sIP9uK/llHKgCpK68VXx55gQFqlBrkzGUqBDlMsF5Cm1/kB6N6G/qQuLLi1GJ
9QRgX8vubj9HYnpZOLxTcQsJjOSTYfQc0Idnn2U3Rq5frQ9zIRfGWzLQlaB4DdNd
mTm1Nf2M4dbdNqIbO77fk+r6m9q5CV9brPLgFBljHSFnxYnoqWZJ3OTMmIkNnMzm
JO6Ak1oA99Zt9u6+b2U8aoHvJdTGAlxVzyQCF6A3dVVA6o/HVogs6xVWVd4fUZb5
Oh9Lw+SVU5a5cVHbqLQM0Qcq4eWELPKX+k96qzqTErRtj1/MWR2zBqQ5Kzw3haXa
4pc9zpi1/pc0lyAA/5eB+3NJB1V7CkeIwR2ZTOEYS6NVosGjrVhdT677z1Tj5LdD
5NfdK6UGKUgzLoCvpqSLjZZt5lZnePjjyvqSkFYsq7EF8Fs+mi9hHwos4o2Bigb9
h9tpfaxvGKiP14RKxArZgmBtfCWWBJfX2PDMOnTvi5XPVu6I0KEZFbDDmAJTqHBF
99ZUn3iPCmOp4e9udZuyIramAZE08iaxyRSsVbxlaIrWHozPKJY3sryHfIoxLzea
F5qlVcv9sqn5rNj5zdY99cg/NCrWTiDTzoKXdPsRSAoMwAF1wfTHRpDJJuGHJ7eM
OpbXKg6Krp0A6kAp0wbnhiK+2xl6AwqKx/m1Cki2sz9I53LAXomujItUTfgZPGDN
x/VE6vYZceW7VzqKvdJdjvgCq4M1T8uwq+KjUdocdnl5vzKf8CrsEY/zqg2N9+Vn
M5/wNmP5d+kVG6eJb0SmSi6BF7e2qTQNa/CRracQiBK21SIUvGC8n+rLOHho+k1W
CArBiyEbQErAHOQo/ABVfsaKwMc/ibtA2fIEChrRX6Slqp5PnCmLAzlC0xgzhF8T
a2lKrCxGCP5IOartHurS3hrh0H01pK9zsujBKk24crDCVBgAcjfhK91KfNn0g5ZA
oxb6GtZQmTyPwwYEsfyX/XssOCyoTnFoS1lufcTpQ16TR8q7SIQVsoCcdoNouMpH
wKqYYFEPnnAPjmYwX1VNVcgKcBVhpAarSeJFRrXwpmn7kHrp/x5YRrQJijIp9o+E
PM9Qww56UtpaiKVHuPJ1qCN1iT00282EoJYEPvfiUtxwZDURJ9R4L21l1hKdERvA
fZx/LH5tEqv5c/VFf9avva0A/fvEO2ye7KYfkG7e9FBi3SD+FOfm28O6Qq3tweR7
xvFeo0FsOUwDbI+isLE/RYjPx7jOSXXQWVKbylqE1aPSGvaZ4BHriXrJN8PFJXw9
Z/JjAuN4etv5VnN4b2FGbeL/jZdCQtVnRgviJ4F3cUNgm0uwtRiUQU2gU79sO+Yc
l09+P01wx0scWcyp4cBXSqHVu0nWTfW1/WSGhbGbB1Z7mNM/sqzSIAODEVYDPMMz
y4BWlTYgd09pCPY3eepJVi6hudpkeyvwwwwhSfXEsKr6/er2Lir29msPremoEKW4
3ud+wFQttBvwZmWOIc+o6QfMPmHqjOkc99TPz+BnyFHEjmcp50sFh+vHDMzD63vO
UYCEcXeixiDfHGPgDkddV2RXyqM1MH5IvlC79RzqRLjOsQhGdNJhKAosqOmc67oO
Kb5DFAqJsJxRdteYQgkUoW1sq/rBz/4CcSP0q48Q3cl0XNUBpu5InXZc0JfQXdKg
DZ3udI2pLevKc/CxmW85iqhZJRhYioRm1FhTEMq5E0DC+z18saISjCMfr8PdTxst
VrWnVbJXNBRO8DQmf7ZEzANNs8WaRNs794VfCHgMpj+3AS8ZIIRzXC8DzPApQaM1
5t6iMsaqzIGb1i+c1j+V6F5GtleqYrHadUqsvRcfz5HSD40X4BFHgov827bRxi22
0nPN/cfayqPXBWZ7NzuUM86fLTOYMGA2B3P64yH46eG72XhwsDPAasTq5Dg0k6Dm
SoKN86TfUBCEZ4IEkEPZjZSb5sp3C3OJRJpVQLihb4xwMt3j03PBkZZhCcDWWKbK
7Yosv1QTKnUmUb0n1s8bypfveRJUgv0GbWpaWH4fPoqrojU9y2rL3g60uO4Gx0Im
PbJFGagIcvym+ZVqY+kjvFZ5bwVXecxpqJm0ICo/JJKo3C99Jbyg9f5g68hSc1EB
hCSCn2xY/k9e3NEgB4rfsUHn6Ss8ufmiWtNaJJgK9OpJRkf0BAUgfuPJCbv6cG0a
SrYxCX8mlVmnZyjQDMYGXSYpi3MEWElD0bkIJ5nAQkijjJ+nBD8m+z/BGAxjeV53
aPuGVW5M95GGhhjWMkPvXIMIQO+o1PwevXxb/eaRlSB2v+K3H0/BiHg9kWVGJOga
vMAjEBBvIXxA0Zu+TsTD2emkRUqBPA1vDA4vtP3q8v9Q4GlSj2flNClPaCxS+rbm
T9qmV0cvdwi7stWeZ1FWKNkk/eiuKtA4l9r88Szr2b0ozIVRQY8my70DQXSMKapC
saMnmD5uYwL1m/iYks4DoOwSUkESaMSfEXA0+fnS8tynzksGyeTkrSPBBaQhUimG
8oH1KY5WnaKSfkf6LUabyahk2+sc7ggqGvrHsEBUohDxOsbuVj0eYcKViwbhxFxT
GTKTSK4SO/erQ0gfITF29M9I3Q9kniup7OOaib5BScDxKd4KJsf3QtexDoSTpxkC
SrG54KknC4h2nUXlnpHSEu0UjBywCNUcgOAWQ+ye8z0NklujDeoeajvMdYo/c4d1
/gUNDytmjBbKN2nSwyUq3jRHx+++upzOolu0QDaTLCPQnll15rAoCy+wnm1Luvwm
16RsuAbMELIi/kD9rDZizYcuF5Q1SA5A0arbLsaLQP9rw4xda2Vajii/pmLz5Ngg
/Alb/BUKX0+3MTgxU0Qx9HbtrScAouhmI4mWo8Xtln4Eg8J8OAyViDzLaLTl01wJ
Tv7U9K9nVFEplCMRj+2nHLpb1Xqfy2B7GqSaEjjXI855K+cECe7QXSAZ9Df4+w7L
F4f5ZhBAz5YNuQaS41C9ozeEp66WdracQdMe6STV+9KWTSv2baBiiYjtxAAgPTNY
A4OWKnVSN6nb1ruEyw+xzt38EcJDwgsAcj/TL87be2MXPH7oMekxhVSRIHI/Izq6
GomT0ZaVq9h4E36T4yHOBMRJMLpbTvhZ8H5sKJpbKzcTdKfY+akwlMOjkfqIRTbg
NiQPCu1JXEpiat1njhHqxCs5QnnCic/1WEwy+cIYEceJ7nWhKTjrY3xUByO+tGch
yyPVSbGHbvoam201B7EPM6MI3UeqCYPetrXnp8pspZ4H99OaEExtSVzLckNTlfm8
8Ka6D5Q8LnRF7Te6edpR8E9Nk45WPkGY8LQnqIlrNTJcfeYxU0EQ0OLJGRnQAZzz
W/ybnkyhRmuBzssim3uGxfJnn2Vqt1kDrLi7xGnFI/wbgMosyrbOArwKnBjlsL24
YUEup1LVqMgK5IG673EIvCOY8LlYafkqbzo+JBR2FHZ/keeHsujrfSTTAvJXLSwG
K2Z7bc48ItBGtvebmZQuh5QgYgwzS2WMNbxVX37YwLy7177EXb/1M1CLpXWR1AWJ
xEZzKDS8RpUxDvDwvvjO4qSzbKHhtpLi4nrtxk3x+414vbA0GMe2C/8imQsgB264
MCgeaZPwCd51riuQPpWkRcgNNCUfngkIc9HsZikiG/4MT1mvjWShEE+yiit9wQqs
By1tBq3fewzndvtFjf2gy4Vq09URBXNdfgzK3qZq15ZH8xRE8V76JXzqhB0FGfYz
p4GH4d3AMReYK8MxCdgikT+hQeTXQyl73F9Y8nWnLpwxr0mOLSYILElOQrnNkTFz
JziCvoP24/o9Gnuljx6yarcXxseqlBltdVE1xL2J4/7twEeSlr+0noimHrxFNdjB
VIXWiD63evVCqTXJCqv7GivqYDqBTh07KBVUIaT6xqdFfcYscfLV1u/PoK9fUPUi
ihcSsE5I/ChvDCFhW1E4aZSwzfVNxGD+2MMjZ3/xgrEm+twSiWDvTgt361UG4qyl
UVSZBJ9mH7uzgVqHu6U4Ttbylb4xsVaSDRyaFMNPiUC3eBXAAGR0KMuxi94dmHap
fcsfEjkwpMSJme5bLuoB3ecmPpDaiSzKvGAdIKfMxUa60qsjG6jExs0oiLdGXkkG
nDyZTYLykGp55vLUVMlK7Ng0TGv/NgyHeTPA4DV5ZsnbKJ8V408hJoy9OQ7eyVR+
I0zYT0tzNHYb3nRn4YoLKBs55H7xzsQjCYC0C1KEvaHK4mNc0G/WPA8wj+CE7/fX
hLMje8q0dpAjUC9HgLwmtCWwyJhiRfUxY3t1su2g9URBSd2BY/bjdv2jY8sgA5Yp
MTw+zXqM1RbY6YLNvEFlnduGNWRjzzmpF5rdI6Auf7vwDb5jvUeZAcOpgIGbaxj9
odJ/gQ3UB7ALU/iv7ClzmvZwbMbIq0+SkSuJDyGzqvjds3zwNLKUxiDVxTe4cSfN
/9d+Ci49Y70E0X9GdpO/ZhMXBv+1DmdqepQZE4u4wb3GH0U4SnRFuNrTMsy6g9fU
KSF8p/QfaL2WRJpcO1gOHbx+9ePmjqpJOl3jCkuSpu+cylzOzZf0AFEDuReb2psV
Rca4++QdbC+X3x2ko3YfrQ9sLa1xppxuKNSVdY7uABYdIYITzEUlF+2VH1uvGW+S
q9vKH8Hm761nY9fRFojZmztR22s4FKfE0lshVnyhw5qXRCg6KDZVpdCzeh2c2dAU
tsNQVsVWyQh6bBXFXBhLT9F+VKjNW5bgIHs8oTstZu2La5pFn/0quD8OL7jLwjEB
cJ1BB1AiQE/iVxs/ZDkttuXNYOQah6KBmbDDuUCM7vhuyTVs8qGTFPjMazk4THJB
eUlleEMFL8tQ3id/iZvn+gXDMuARQ3F2AXbXJjMvXAcc5ch0gASgh/QU0fPf2AlB
cCqUrMf+dvEioMcMJKCkUeCGQDqS3IkAtgeVMkD0yVBjBM6nCBXogOnlLC0wEHPA
981/bfXr03ISQ7esbZ9ON+2c/NKQlxbMX097G7OyU8GxGkELKQjZdOzeZrGPeOwP
3P1H7WuW0q9AS08MD/ywX77rzIrLka0WX/VGAj/v42BmjyQ8GsURSCsQQ6JLlSVn
yUo5k9fDn7ExhSV1FY99CLODZ0b7x8N0qaH6ILLr9Q9pZf4s+c3r0UxzqE2Ebfgk
xTxixw/3Gkxk/6ltqxrrT6whaB2GlTmcwwozUSkhW342YThROhwi9mNJqVEYbBju
tz2LcBFd7XSgymiIWpypokL1fXcqToeUBCn8KcxrfoEB29KfTu+iTvK2F1Zk8xG1
20CecjEZTKMyuLIo2NK9YqP1JKkt2eGzjBTrTueJaIZ8QayHasgjg1H0Oca9BTMj
uWcXh/y3SwttuNTPbZQzuSCHdjSNZ4u/EyPT4XOGFw6bI94wUz1GlFF8JC8ydg9T
GN8fephZx+iJLhRI0iRNZNLhI1i1V7HuEaP1Z1xWYDc21dPcKJSIVWLJXQbuDElH
PVwG3Zzwc3D19T762ceh8VsIcUXWze2DaV0SPsSShX8gSqh7q2J8xzl4gLvTvVYT
8C51FpDAmgTGx7nrWpMkW8Np1sQ0gaVNm0C+7/tQvUTjJHcKCYYlu55cfyI9W2yk
SVav3DKvK85JKz4XFC2mLjpZCG1kc2lffWD3ckeJgXCjaNoTQ/ycT0QOA3A/eRKp
y0Rox1SuTldcmLdv4Hx/xooYQBTfOiy4PEEaHs03K9531zFiz3RqNfoz/Kxk9C4K
GQvY7+8CPfssKxbp/Sbk/C7LgaZHmcPJ3dL5UCYhZg5qiHZYyrC+Aud42HDQU8JC
RVsZeWpEIpQ9UQZfUq8g0BT6ao3sGpN461QqoHeMKW3h4Hz/GeiqTwMWzaR0K7UL
PwkszDwMIdmxtPX5ieS19cClQN9siM+XIIgwIsC9gmcGmydv9ds93dfb7z4JMvW8
zfcmgA5uvq1xj+PPMaX9mrCxHGhNdcHfrmCuPibHEF95S3E8RZOnJ/kmXNnUVQzf
cUDRu/Vod+uhETzeakAv22oKYlFhXUd4p500+Al+iZO2Ia3eRaUGU1ObnS4uO9Xe
TIab5l6sC1QXR3W6KN2yo+vynAdqzzjW6O7Hc1gnpJMcg9A+B2D2GZLbRmi84X1t
jbKNeaBODOdRMW+KI69A/O2ZhNVQ0V3epflzNNYho+VaaofMlV0OlrjgZARdmmmV
6MKRjUTM2xKBoR1LsbgpW9oQjMxOULukI+XxKlmZ5kXEbOl8gXzLle4VpBzoQN3X
f+aopf4xhMRh8VeYZFrFyTQhapdhgDP8CJHQTLxoMa+VHnPsBJPPl1f1OJm4610O
XP1kKOdJD9Z2u2m25QnRAUU5OuE02ImQog1bPD65Y8H5YG3tzmxpSM4v9wgm8aiU
z9eWCxN6PAkcpBzydZn278uI130XzfftbV39Esh2j9HjaUgOuMDH6hysk4l55+gy
fNqhXHXwXcMCKx/g9zsxN5E0TA71YD14nB/++omGuG0sLwnjMVvDQX9ymd35wgts
Sr57IdHXjgXXNCOuqOjR3beA6n7ACxRXn8+aeYbsO5nn9wuhb72pqX9IE/2PxDy7
xODuxw2FBdJ4oJWGDw0Tp0EMA8Zh7EixelQ2DgtVCUbld5qhGw4XPRIvIkWDVHsD
/nkPIZdAwfv9Hhc5k6UF6KTcASJIOlpl1oJAyy+KFg1HLM35MdMrKnkIwUIPnl7A
ybMZo3x67x+E84stq3DuwP+r/xQsxqG4QtaaRzOlmTVN1VLi593R7p0eRnS3Cd/G
j5DyQGl4VYI8QvQ3EO7mBEKqLVzMzxrLegsqGB1FY/20F3CCEVY9vi1rqOPFyIMe
YIj25kgHLog0omSkzYToePYliKhVbS4fMp+nSyLe6Mbl2uBTfAfAXhRs0ysKnbih
vvUvW89iTMMZyd16lWQZUCNyWQNDunETqb8O1KxSBMYI46rJKAKMv16/oKfO5kaS
dmanue1G/a7/ehHWT4GhOl946xwlluAu2JqAyqQ+9mHhaWKuviCqCXifXLJUeLJr
kXIPMf0m0X0z0u+n7zsAo4yn1MjCSfmE63O50pjBIoJyWqkiVB28MORGfIMGCxUt
YsxCo38zJL2Z1G7EQ4RBBSdPJnHDQhSkFK3+hT/XZoCU/ZRFp7CBI+/4kGYXpHZx
POb9PZmprb2hmrpyH8NGJLU6ChDAfyZGyiazp7ybdC8F3QczTaYEt/A528sI0kMt
fVcgPc1BkVWKhBr0QgAp9255V0axmrfzxzfU9Hk0gYPfF0YIhW5DN1j27T2yKBkM
CV+TZkD8cq/Bjws4RiR7LX0Liutiaid08I4sFWb4RTrNCrxBblyHXYcp4J8G6mXU
+28Z1b3qGw5ji+0kAYmMI+VYNggKKghGbEOnFdr3Em8R+54b/HFVuvrazKH+urP9
BVLrDfuqo9bkcjC3ZCN+fkm81DMLo8a6T353ohjkAfeoumIEqRAwnRzeYjZ0Ft3U
J7J05hElPOxDsMyRl3pCx0CZk2o3JgMdx5sHwh+mrqy9Ce4BcvSb1ShwjB7QbUfe
i6+YK3Uc5qXK1OTvPGLeUZ5eAPnUtmO/ZTOz8RDENzrbV6wsrjw7xyItnTWLn6zp
NwovEdMrbzJBrfi3uCbgDRsG5RRVXW2/EGHmpeXkeepcUifaCAPiPRdj5ZyKoUlm
Ql9P0GzrQWgEHsSUePXTB5HnC4QDYQ+gWBxb2lVBP8Ce4bIO4vbU8ACVERon4K0/
Z/+/uH4PP5JYfWRen5wGSrb7ADciaXOYssBfKovK7e+Dz3lqsukTw27FdsiWUZqZ
1xL4mhBZPcN4u5c+QJ/VK5yEQ+EsUKwpbVnWpH6vOIWguYCfVmZq2dOgreAOvstz
PK7JabdZeuGqJb4wz2cv88ebdXqO3rAmh7b8ZsMgOYS7Gl8zaBUBRbrMDk6IL/m/
CoIt1WK0SYaJ2Ch6gDtaaHwAgRUCVa7fCeLExc9wTPg3MkI6XBHOrhXrMcVySAiE
G4ciz/JgPx318VHvOX2ZpvYextO1OyC7Q3L6jHl/3doZtA3ohzMZyk5HoCPPUWeH
Y3lpLNXWAl9uEPU/X+aDKJkebOmZsXEVdnACunWgokNlzjLYK6d1yafvFr7KtY+f
gYPUXowSf+Pc3eiVrD91OIL/iMQkJdmvlfnqgK/PgxTIekWlNgAGvTldxTAIEL5k
PvtwBGogazjpgm0fExkzhmutIhggVjMoYriZSFZKvTeYEP11OwvWZ+nb63vk9eQf
q7Z1JIpRvlD0eH0FCvaDeEat7fw9Qp/FaDqQ6tf6P9URtWTeglsXEQhr7ID6l40w
JmHOKRZgYpCOC6thDecCQCIEFVb/kSdMUEjJiluVgUCzpefkK0XcVGxENPf8CyeT
g6UY7wSxr/n60fvo7yP9bCHfEOH5y0gm1pEQVUJMd/EF8Az37plZh+SwvnjKRdp6
3MK+WHMm5q8bGEJYjUcATnd7/z7zIcmDsoyDLldvIggGh9eC+/E2KR7x/swj25xs
JkhA/16kl8qneG2B+dKVoObVK0grk096JIIcMD/vOEjDIBlrUjI+A6biaJA9QFld
c1I6JwaT8p4ZgpSR7Sq37+XpB6wEUbMzMZD+heiovufQr3ACU/y6bYhmNQ5XFKS6
xdxe2Z1dv7dhklGHrRo5mliYQiBQzKYspSiIh8F5QzfDw2jrBRWjVzjaUrlv85Gu
+SgjJruJ2LYpoWRzwIK5bhOnM9SppPGpZhElCufpT0wvST2tCh4zX9N86c/hR+DD
P7ZB5M0XLXpjlTiF8SUUhmisyjijHq09mthRGhQoUKeAVXccNVcoPAbtVTsi2Qqw
CF4ozbczT68c/bcDXAdQIQSE2YORwAIXc55fZfHpf57vvXEMe2G4jv9kolUknSPr
CTmidWQhMSN2Z5GgA9WmjukFfePVzbYCrcXQdPqHTRB03Iz/8VwOKyKm9ZcG99H8
etlFsfBeiyOtOQLGSlPJQyJFDToyN9uHyKzQBZKX6snonldr764Ylh3EMqn5w8tT
bHLmICzxgcSAEyl7pgcP9eHvvZt2ESPFxX86BK9VHl/kOyQKGuo+nEKqQSKwVQvP
uBCLwklb5MzrAZebvoeClstOgtfRkFur1Dn/iHWhKaNpVg+69yAY22KKuav3KHyo
/xVfMuzJJYzdWcBCPIq6S90z+SRalVkZqNbreGyFx1JIckGL/vTcJw+3rs7CSm2z
yxTWl+3LNEZSbX1N9uh+AFpi1niPotlzqzlZS9FI0HyD3iWq2CKeKCdu5qUuwzRS
5ZKGHESKkx7GrUQeoXYNI9hhzVV3YjAC+JbyQBwjmo1XOQ8Czk49P3QCwc5VGSA3
Gxdk1UQXULv3soDJhczAn+1OG0SACUBwnEXINlO7Js/UJa3K7n4TcyN3kJvb4ntY
SvTZ6f7CzlxKE2Q0JlTh/WAuL0eQvThF/nV99If7CioUAG9XnUawZY5joqzbiWvP
j2nhrfBDIZkeWLK9R4o+DZgiILikpa2YMqjI55NpiDr8xsebPqxF4dug4FnT4E3h
bSg4oNNUfYurUmQNgfuh+yK8FM3LpLhJK9pxLDEivG6nkwm6aJTVVA6wy60MED7u
xSfOshMHbvM/PHSeOGBwpBF3YE1K52kJPQ6FVDClsLaLM0hNNhhAUyPX7WfRHrbt
DB4yoowjAe7yhWkkQgWgmp9OjLiX9bA+XEA//bgsxG/pVXj/jzflI0wBp3arqIaO
SB9bRQM1zD/jbCq6JzQfoxm88o6hGmhRDbNwWLDMyyWmZQx6p7RQKCFDVwSusvEA
3ZamGJWop1fNhDAzSUipNqeo7kv3Fe0CUlliNtdHSHzrRnbCyKNmCuyD3MBJ327C
CVX9yhtiuKNxgNcaRZjxQJOR0/DUm8TTQAks1V0uf838JsQES13KGEFR6SF5TQnx
14EzFDJSjDJAhbtWUFT8ioNQNz2V4BWYJPouBfvE4DCh0i4fOBdlALEQRhPa8tuG
VGgNFpBOnZRl3syohVQ+LKUDAaC+DQjJvkLO7/yNHs7iREJj5Cmty1GhgUnCUAXK
SZrNgYvxzBBaiVlhY3WTRsjUstE9Gz/XW31BTcWY/gn0KHyM75nblZFjQEWbFERt
RGGuJxg/xpC6wlW5LWf3cDacR5Pk/GWVJyOAL5yU+QTVsCS4tOFERKC8thUMQY2s
ZUotqdHz3L+OLdoB/pYRrKEw3CjjhaIM352fnf8SVE0z4oMeWO7OG4F4h8FMaM0D
lRzwqKL3G+hmhYR3XoxxyK+fsKR92Q9liSdC/2DXDX+sa+2AnkuC8+xVE8/Q5EuE
Ymelr3gzz5NXmPmQiqTkeynPAx4bzYbpyxslcdlMIMzw7ZinZLKPYZa/irdEMcWf
Q8vtgLsURVe43UjGvNfatbDTjaVFeugzFDo2QIc5RDo9aT8cIRnupCyB6HnM+FWk
qAbd1/izEvWcVwRYH5UKwG/dUaCSonPwmgiPZQ6nGdI5V/OrEIYrFfqxl3r6RCIa
ZNVwkHNrbh4tDo8oqEFrfcFx52PrL9UtXJ8KZ2JpJFr4Bj5jYua7S5M2z16O86lB
7606Dx+A3QicrSD0IkM03LnfLeWiXZDC/kX/AYGnFUzUf0nuHwTnxU17ilghUKFy
CUTQDwr2fYKS9jAtpfrDvhQQVYhMDd4yJz0FEZVA31Z8hDaSJPLkyjutjdftIs/P
tRd7Mp1q07JUFBaC+2+PUrKUnHh9pD70c+oKRU9wFIiJ4kEaW3e0wbrfcsYBceHH
Tr0Ls21NeQQBNzrj4Z5cCUBqBr2KfDuJ/vzWazRKzAOj47NbeUmL8enbIsLFtcAr
32YtO0WIpnYBWFWFfh8qeiZu8jHXI4D+ayQRMgBreOkzL1QuDQI8ooWjeuNqsy6a
WUslysi4TAlG0Vr8lHBswt1/qd0WEvsYYEdKeamQCxvyt6GnxlA6VtY6EJGuHMFJ
oHgMZuZ+Cp39jugMLjlaErdgz7oL6+4XuQmcfbZKxsQywhi7gYDl+HzWgE/PziHf
cuEzyJwUtvLGx5OAzjWn2O6k7A+eupsCGkSRKbMlU48EvQd+pC1Da9swshv1rdIA
AenuSjLUgAyfQAa6OjY439ZiNiTcHuKKCER6ZMa7h6KeV1uR0IAoUBOVry13M07i
IQWjuEPchtz4qdtoTq/cP69Nc6fgA5f6HYU8n1BGL3mkJwiUmm4RdRo02CG+0SU1
hguMuh54xVrA3DxCKAVg0/JUqoIFn2P2LtAtaNyKSuLjokXoS53Ptrlh9vRCiGRJ
jSddW6xoCLeex4mxNozdLEKMCYwF1Z2H6OzU1NyHqMfGj+VNB5yRZg++LOaFhLXr
aYhOqVued8T/i34BUAVhzV+pziHk27v9/sh0aTjjoth+If8kxHX7s1DAQOGK4J9a
XtTz3ykRYnYF2Zn6bXEq42Tm8T5YWua7RGRcUJWXKsxLlL+bOZxH+roHtDmp/r/0
f9STTV7q6MFtCcG5L8lOcI2kH8fEyTQmTqr8EGhXMbt2MDsv/7rM80uuNx7t6Lq3
Tk2QK87r/80iOai2MfWmySmBOsDLNgBbYgtW8GEtsBca/PBMud1kvqHiuKjtE0+S
X/w/ACxVtPsxj6p8lcCRDQIX1PBRkgCzkHHywIT+OK7NaITMI377d9dtIz1u++nI
oV3dYeuKXeWetcQqP42EU+thVyGLg+YFlee6CdGIVC+ROJNoHf+QcJtI+VXpy2Gx
WDCl2SutQV6z/WziOuRUtNogTG5njXh+1pb8OMvcm/cmN1lOROgV5JA5gYRmQFVo
iccfJ7IEhk4lT2d/cj3BUuWt1CyDvYSs0oZaWZL7UsOKF6spR56oEaLlZZRrwhw7
idmGeJ1pzSIEuqfGl6navgx0kgcsAJXVQsdnWpRgo3xf1IiBBFVSt+bOF4MXQd9K
7Hifjr/WJDOOPnyns/j2pbybit9RwxMuO7ANtT/01cNFrtXN+q1HUDeZCtEnYJhR
ssOJkWEf7Gg4WMMw4Eu5yxJkVV5FI9z25URm5KbFhejTsiPEvcmfo31bV9frNCmF
+ZQN6YJJpuA+qWeuyXatr9UJBRLucbKkXM9ditl8PKvO96NIKDZokPC4O3EMR/Q8
H+NKS6RZ2EWeUlTRl8eEAFkqsYL296c7tHOkgVfZ5tyJMwfg9y0OY6RqIY0CRKVt
pUJRb+9pTmRsHawT9EuRioI10ucmMOl0krIcujMFD+vFRxSZW/Uwsp14sHBrPLga
Zs+TvXC705UDlrrO4V0JAIwSC778FTPr2Fd+Po/EpqKirE8FHcJsRtuED4g9VicK
sjMPb/WKm5zxSY02YKLr5EeWaYy39hgcv/7UQfcijdYl5wF+q9VtMpbTKH4taGkb
9SP+VH7g2C3dzLvUljGTdCsw5g3g7wn0dc5Z3JtZ2S0HwB50Bu+p/JivnOMmdTdk
sXLNmFqTzcDAwo/A5Y6bTY7oQg0FHl1hLQdqRUnoGxW3zd5er4DSmnyRpH6DClGj
CHiu/7TbCuSHKWLRD94uAPOfn4379HKWqJGs+s6e91kTpe6Vo/yU2yNa4alCHRW0
ucT4O6+hKw0eZLV9gCTk331xI7wpQhx/MMIK7S62lpbCrOTBuUskdva9mXMoV/at
QJOk0kUDPWL87pgjXLPjGnD5ERE9PYYLSk21bGxkzybPDipc+pKQ266wpDNWPvez
NYaqsz20kLDxvTdkHHMbJ0E/zCICWAWDqGx/CxDEwlyY10crUpPrXhA5huBT84lU
NJUMqXUIQ13IeVQ7I08HnMDhSTMoBi3f9aklpi8heT87vOkbW2Lj+uaBrQi+nSYR
7U8jEXRM7JcePCDW20gDzczn/IgBGBQqiCdXlfHLqVOlW0ZLyOFapKtNm4EeZNfT
hms8vd4qnq1x+kpTS4omb1rEM/Ir2YDu3QZ5RTa+R56QfVU/MlTXmZ+iyeJGpAgX
9t59vR6LgD9epMZNUq8XRKsF5LIP+4Xnh1vTXjIYb2BKybNzjozP4WzS4XMF7R7h
N9MHDiWOvgMUD3jU4l+32SCGTdjeGkiO4JAYgbe7tBPXfM5BLIp5sCETAGE79+Zq
3VTanpvPCeOnCGpFr05XXUihr+2Drdsn5+8M9alCIOm0QG9ntOfDCk4g/hvvk3G0
QYFpHsoxzlJU+E/5kT4YzTyeVQXFZxJuADgfH4Jmi+4pyQPXPZGOcQDoAsOuZn4n
OT2020p0Q5SnlH5kuUlS4QYRRgmdsCxSrEJDYsUPhxMgsWJs4BT/f+KxvDXbRAHi
jS/RyA2SbPE1c9eZmkzAIcsl8FBe7T0bbOwQu5OVep7YAVjEy3MmooTaHtM8zBqA
41DtmYA21Yh7pDGvEU/+oM1JTNbmN29WVaEqWjujKWExAgt7Zx6TLI+VOs2fkYqM
u5hoclscQ/6+rh1j29xR8ptbeAnUC3xnC04BaH0nJBkIQ9XMbSVISbpFLgA7QdpY
Q7gVP1SytPS+rtdIkWW9+K59OMvrWqyvqRkinwQr68ghIw4m2M3L9iEStk2hf/qJ
nWlnnCQ0Gfs/XJ1CeXrM1NWtp9WFCMaEmjA5dWYvk/edRSxqAEVpgrYYCJw//z5F
Cvk6OebeXklvQWtHh8fc3a6HtsBQwLuzut0fyeqg9RCcken6jTAxe8SLn2r+vWSv
Y7wRjVHdU5GuzsNrqHg5KUmsMC4b7lPR3BfMxLbYyurU2/fieCk1lQDHqwMbp0jy
Hn3VkqcGChch4OLggyRvF1y0MDUV7l8LzFdis5UdKEDOzdpYbPAimWnAe6R3DRWd
uT816rsEVvKQm1LjfJW0kCf5Ao4v4C88w6xzvlfGTWjh02cFm6bJgVlgiOYUsTnH
HoXRKeRTUmZTurgCeyX7XnyNDF8snbXDH0Ll/QznyQMTmu2daqCsiu6i8FMKhZz5
31bvvU0p6jZScxUkjHCt1KGmYQvbyu0FvudOYhaMGkiExiu5h2KFJanEH+hvMqVg
cxjRiAuh0xLJua5lhjO+NLvC9f95k/3/M0cdsB/DnK4ml4iTXylhmAEBKn2rO8/R
1HudFOrbTv8wetcUQ9MZVg0iZHCXxInrd6tDP4ptSreXbOc8ll+hYeSrg145TycT
qE4VwR2eeox6pb5dJCoXaksDG7oexYtODKtQEkvflH4fa6caO64UmUWFSWrxnz1w
XxNIPZANtV5P0pPO1cN1eAiwkj5gapVV0ENzKsHzSd23jHvTe2zfDTk1qkXoig5Z
M1PHg50rDO2a5JyAMO97Jzy7hreNoomwi8wF3LQ/Te5QULwMuuEDbEwqhEJMpNiN
rCqiUn9CwHon1zkD9UH3Mdr8ERM98IAA225a7hql+QmCW7xAiHnLGebPSt/vhR+3
mtYtXbWw11k+PlPBNYqKbLvBGqeVp8m72H8C/PeqYsuZVFMeM1oPKje1uqC1rwnX
uJDUYY/nyS+OGEz8JVZwx8xjrzjpMjA0V9hXjB6+x2PX0+WkQ1p1KuUQo2toz5PA
JhrWYMIshVRJUVTuM7swKmqmvGfPt4tHBfAJBUAKL6GgTHaac9xQSuQCw2kW+l1F
ZDVQOBDmIRG8ptxaEdc2pmfdOmvito525pLKFk6nMb4qNGlrtvjurDsRZa9wOv2i
fWIzKnFw4EnclWA8aN1hLIA4ri29PU8/8Qe/f/33KVsUjzTtZsPro5bV/JJMRJIv
l8k9MEdDsUuuVEWLNzH2XQx0hQrqoWl+gFFltqVmd/bRiyOovAUFL1+RS4yQuw7I
H6F+dP475C6PGG0d+9a+7mMATpAtCVJHSO+3h4ovF/m+yiSYzC6msXUYTJAcMjDB
+rOYYdeXzoahjwAoE1BaDW42bTlpZdlZJSQRRgE6zdjD8FXwDKbUF5kHdCNkkHnq
kOzhnWpePyO345gseodDh6hwHiWqAcgAP83o2ntMk3n04CaXCkVIy8NGF3KeXOk3
YRGCDPLQgReHhsIaG8pF5E3o8tcCfE+C4l/6Zk/qfFxXLpcNdyX45VfcmAbvu7w4
7ahDF5BCunc+xxSu/82F/uum/DRFapvAyf9Tz7dn0E5MSxnPhOGPFd+VMZjaA+A8
OWsudmU8UfHJ79Lo4MqS5ZUMxWD3ZhNJ0H5BLxqQ56YKP6asAjaHB/qj5Be8xney
IxYqYrDyH9FQveH4ge7fBIL3y8VTPYTs4gKq6S8QP0VHyIxcweBi6wkGfPQmh5A6
VTPcVaCL76FK5MVZY+L4I13s+W1WTJ9i7Zk34c01DywGL9yF0mmfn6lOWxIupXTZ
lucnIHrCCuPurTVOQMXWpke3lLr5oJLJkAmqpsGFi2UIwBJ2d9mVfmfrZR//0N8m
Ruq+oWwCgA30dqyHHVO+9AoVisIVRi5tzs/C27lD3L7P0xqGsD/HaUF0FDWeVLpK
Mqg4YjL1iDo8dyXi0NJib8XMzcfRhOyLAa/bo+m0qDL+UhRZJtYPHMHyi+534Tv5
VJVR2yCU6SNpXJz1xnElm1OlzaS6rna6cEmVXH8/xblxn7CRSB1Le+0V2cmjvymp
epGst2ZeinEyUOS+IcMpEW72gHSqvT2SNdO5ZvENe17uLSnkQKhLZgCX3wN3JDYk
UG6+Ee+6En2AbwOGr1Qzmsxwc2C4JIfmYucT68/D9dEvDKBTgfJwvcLp1OiCtki5
q+BYbXsyorRyiefDCp5g0bj0B1QcoJcFVR3Vvb9+b40cIetOuYk1Eu4z1HIoTXJd
hItF6MQoXSyrIYxMLTbiRL1Txt67D/e5cVG8PtHJt7nSMCVSwJvgMXjT0VcZ5bUo
ZMCPFeNzDe4JQC7zI4KaoplXrkdx0IxJGSzOenzL60B1yfG+Gmr1ZDbGmnHOfioO
oCvRTTG2EJ7IQ01ee8D2TGvq1C6Qmi+/63uj+2LuJB+hm+DBAu+7p+TNYgq84gUP
Kk+6KpGye4p/+IoC/CZgeei1poWi93FBCe0vF6PSQIuKfBWbrGon1kzm1FVKBeQa
/sAOf6qnCysdDNWY4i3GxZcWQy+dEmcQvqx/3iX4Gr4G6Z84aUER0FeAqvM4mUHI
UAM1/oxujPuzaB8H9Qo38M9W9baaOQ+6MbDb+GYv3A3Prt1hZPAG70YWfWpBFvQv
vIkpO5lZoT+vNbd6ykNOwSNmfsVSFo8cPfAEyupzW0sHyFzMoJ2qT3X4V8DIHS7U
NuFw8kOjPQG/SSdKBpJ3BUw0P62sqaCUnHFKME6aiX7mBG5KygLENoyIqASnrzFw
w3NuKLA4uU42xoj4XN3iSU+OpwmzKunEvt68BMt80LdEUB0m9ckpMKTTRyb7xvCP
qFFCU+1caItikVEkak14o0VMPQ6+6X/eSd5Dh4IppJUStm+/s+4DRpasGQiZ3Miw
9KNSMxdq0SijSLQa5yMu/cxDqBufsuEEFYZi0JfDW/WundEcTzIBCqzbLVznGspE
MO3nsdReVsMmfNyNkuVwWIEUa9re8+cuXMSMkBuzuE9oTMuQWCpQxeo3Sy1/NAqD
zBAgR2SeVknl6QopW4k+1RGDetGocYPO+XS0nxUJEvwhChohcH6lRBVn12Up/aQe
1h8IJ7RYHzXpJgTzCt7eUJKJ5KxM9bgGJi35o9Yn/8IjvJyHVHiA/yH+nFXzTHq6
X2AiebsEWQ5diyr9PhegkWeOUbubQJM8IAuAzUsZH3Z6cLhOLl2vU9owr2vF6537
F0Svu3MBFVPQFwZbxaC4pZ594JiKlglKR+7dexD7BKzpZuGjPvRwF77/gPa4NEzh
LR3NpQC5qPca91vGs0I+UBLmypSjt/tfvwC7zdcD/34vOFDktDJRPx/0MgBagGdC
3rznpRo7TIaYzxsn17zgW6fNhU+iekY0YHRlk4Y572UJMcllaoRdubfNIzXXUqUz
CLdZNQhSYuNxFIJT5lLnRO6OD51JHYFQR/q4t0PE64vvLEr/aJ/Th+C2RF2E6uCQ
0qxR6eklWobwOr6vMXTJp6GSz3tPNOGdGUn69ZcVan0/xFjExLVYLLY58oFEmGS0
jRcyPn4oE9kKtP1eCs3C2+ILttPDWjbe8E9VWzZVr5tAROenLxQ4Tt5FWde/F2Yr
LGMQIlq/ywxoWA9WV66I5ShPcg9DL7U1cAVNvUaxccHt8hTufTlIS9FJpLpt5Mtk
k7byM8Yf/aYpRK0B4Faf6okdXt2IL/kciIavPdFcpw2r594KjxYdW9GWlnQyYbZh
jhxyTWx4lYW7wsbNEKAKXnDQw+w3yrCsvhWwKW+rvNV7OJkQ2HXWg84n5CicvcOW
US7HVdbVOV/qROjwe3z+yp5NFtRk1rX7XQivsfuR7gUjiTt7ZuQ1uuT4gQ+meijd
2yOJoXVck7L72ZY8FOTxnE3dNz7w9O2kcyT/jxJBx6XerM1rm50l9BpJ1fMMGZAA
AZL/ALw9peZwUQ1Q9J0yuNUGrxOK8vpgRTxb51y5KcCP8ntUrftmkv5c6efpybNJ
CVIMU0YDbX6RlWTYQsywj24YcV+mjM5ZlDzql3005eBux+JEUYyaR/Ad9Q7477Go
4SYEJ5QzuVH6iYcI4lea+CfWTbXyPV41+1ajyRNVKtfC/FWeNe9viAUBJd93h4XZ
xMqGw1IcG4NPIG0mAFKdZCZ5lbK98B/fox1BtyZxvkUXc0U9opiyWkSLNZQ0qPp/
WwDmMwG47fHFs19pZbJ9mB2WIAcPRTLwe6ttf1ZdeSpsK14e9YxS1FiU0OvJonkL
wCa/Inhimm4KnToJh2Zadvs3SWUQr2Qg4Zq7xpfClWoGLFijes+qQSlG5rfTKRW1
i40+IQDFCyyfuwz7VRz32PA+uNE6G/l+92SVz638b5D+yR7TLK+WFipjWh8mSD7g
UdQyRQboIYnsyeKtPk7WTIAOpJ0mINgUtluxpUSzQ5ghJBv0/ZduJohhJjeg23W6
zGd2Xv1oxYXGgd39XxoF+5rxDoc6iTMxnRDZv9wuDd/OPawsH2FURzVW2xfCWwM6
Xi4TSfgHz/UUZNIynMDAPaCLTrXXwQWWCesa/mY6vIX/9eXMEeIx3Aa3HOT9Ilt0
9tVcsKg57MGpv4MENSXVwUwMHphi2mrF4UCTt/zTEQ0yEEmCIwMw2hr37lY4QPiX
74RXZcqbO7N0BzvqYdW/Dse6balemMmLJGq9029ZBhdMmbJDN6Vs8lTqxideIn3j
wBhShmTSTafBH9DW4mKTlV8txv0LBojWC5fLAzfOYEuGOzayPUGKcIHPDmhwZ37w
XUnszbagwMiboDKwKalcv2eSwuoxX+tlqwu/TX4eAUEpd+EeddilD9plm5RTlWRX
m+UzLxTbLu8QBgw8ZqD0vL9z1nA1YaG4b/v2gLR1VhzUBUXRtTxXidw7SGOBlDyZ
vTzmhP7K+cxxJgNS40y8XoQ6p209qMtJroiI/QQIAatDQlhZqe0QeOfona1Hf3FN
gprfUOHyxiuHg+LpR28+DpbcZDXOHDVGipl1Yix0SafswQFJLlMGPgOSge0xt0TB
BmN+gujcD/Jv3OPkS73cYawdLmzl5Cfpp/iqT/cs9dE2SQPy8U5o/jdaAb99HzIh
NjkwJXRABkutXzlM72SIx68sHwAjS2QkXLjZ4D1KHbv6Vo9bCkKiaHsofrSZUQb+
vJKjiv1nQCuZr8tl3jV1VxECA6ktB8KQhm87EUjfGSOPlbvd/StoVLF65TiVAQPd
6kwbJ6ppwqFaH7Y6KYEzeOoxr57yvp1agE38/ZYMM279lX/dkN/YRNwdGrxOS6a/
OugedtInw47m+saKzYppJRYrgggjg3p12gih4ryMGE2L57dK4wOndO+Fjs+Y9G+S
yvlQiL2/tMJO7D94lu2eaiTgahrarux7CoUsgBD656FEkPMKdHM2VsQ5bo2b/lHq
l8Ziwb1cfSY0Aqyvow0/+MmARJ8R6cH0R3q2yMhdZaIVbz99nGrqxPo895V8V4wX
yEMeVOcaZ4c45wJN+OatB1cem2Pjg8k7tqPd7xi+Mq+vwcvevRQHL3kmHDdcI3Qy
iLHbujYPnfSWqYEJZT65024Pdw9FunrI1E9o4F2InTybEQN5NHB59EhDn9wPFlRw
pUvzbQPrXhBI78yPRXm3vySuKyvILrIVJYfvoLecKsKYnbJaNO6ehbOW6457Le0h
P+SVeOk3aGfWlV+jqJfpeuS5I1FTeJqXdpH4WevliML51dz56u2S7zkCUcdG/CpM
AWfSuzcKfwxUkXBwH+A2MYt7YLbXObQGw3RYS+pCKo1jsMeTINMHRgdUaaZa/nUx
+Arp5E1ruiKqGLW/14xHRWlHT/ptX/D4fpS49r74xFW+K73jhGLNfVxtdCXcAZwr
sc9p3TXsdxNcmk3sCfWvqSYgPHGP1qk74nVn3QPrhcyrk6o2DnomoY8/a66yzhtM
Lxwjiur3YOXu4U76DDOIOZxMlGhbPVFECzSfLKgp/6XLPEvXkcRmA9p/wP5gDmSt
LCPL1HPDmHKDr6YhOaXM/uBZeu9p4Nsz1Sp72BjC+44QuD3z3dStizwVE/1x26HH
N7sG0zrBFMu2ZdckBDHpp87aggYBNtl9Nsurf+Q18L718pPNzqIQuWas4nXonKGi
0YeL+ZwadUOqOAst9BZK8Q+hrhtITunXJiEsDZ6GrVUvhOaF9BGeBebwGwfY7DRi
eecfX54zTpldJCDDzN7Zazq++aOZnwdM1ilrfVbYCRCiP4Lq2d4iBy4ODRDDahez
cc6CS8fx42VlIeHjTRv4f1fUPprM2oMpqTqEOocbwDFpp8Lm3NmvDOQ/UJtYjN39
hKay9Nv4vwA6+4R8zyXYXfNZVtoccE9YqVjd45GjmNqPt0K0aokzYCE8Ltkz6eCv
yDe96sHlFZ0ayhEuJ0LTZGVtBNbPNkr4CE6eQEdHCezo/a4dK76TEOLKMvlEgfiS
7TcIqyyAnuEb0/B40z8xhhoUTEGjCRB1G9yZhDH6ammvHi6jtnl7CnoNWYVUXOp/
nK6WEpDh/UIPHIDcy1iXQCeKHQSuCJRTABcvgc+uwNsSiMTlbFMy3ynPL8o04qdl
0HTCqY5hp3HD8YQrluYABvFQO7KILTzCFn1GUqpbrgjkZWLo+EPDpiOI4Rpr2Lk5
JVyr95A3wjhC0A5YdqNKDhPGLWNoS7/UkUc6yDhQH1ESh9HGT5AFybMuMr/We9ey
1UvOX/bAWASF03sS5JLO6r3P1fi2jqfyUCSOHeyQilmbzyxHHgcjH01rwvMmpB0+
mIOw3AKm2KjYztYG0qvzqki1oKO+hs5e2q1ZYDAod5cU/aYZoC87dMzWOGVjrX/b
NAdTdueCFZ69FaKXQVNMZCSpsuSifDtKaGp1lBRfuz9/8/Z5ZAwPr5BFbUrluGtt
4JQpzM4oTJpYRdJZ+gsRq4y6cWhmcxMOH56MLPwsOd54tJ4Tg05FGD+cP70icc9/
bFEFbUliaonK2Ip+4tVTEMceycMpE5Q2QhNcdaXXx46AscfzkuN9P6Ic5TMiJkEx
1Jyts9ielXF9bjntFmc9KnD3MBf2v5ihuIqYY56QGGL8BQXNrJ7wOLT98ENNUtay
IjqLbKM35YMClonm/nhHw6F7BsZvOpSLaRsn8MocrrgCPwN7DKnkYmUbzoPwRYqL
mYUkneDRXoOaoiVy1LKsbLpjO9f6TsPxf/CL+p5NWHe5JmSJFCwzMGbD07v86GSo
y/cTcxOYNCqqSBi/4XQx7HZi4Gb7hK8j9+p0SH5bh+FmT2kveT1FO1x3honVOxZm
nOVXAKhLvJi8nMYRLOU8Tr2zNMY1BpjxUhyUZuC242SaOINXYj02e2djfObSxguq
V0dcDjMpkJPiHbuCx2dNIZvnw+2vZvrLWPca8/nTUGEF0cMd0bLL6Zp80S8PlSXl
f+4yq/ABbkuKKcvvLapxR+PWVesf/aFz9pZ2QaGUZ+V4ohAzoDbyVuIgHscn48ag
mhAkob/cgO3O5wKmxX+d20RUKOEhr/O0gJT2fdLAe4VMUN9FrEduj03enyMBfvaE
+WxivpBWYUdhqVriaeH1KcLtsS6muAymsDj/IQZE4nSTxAHjEi/j5Ohq/1fD/xju
Q4xegNsexQ4wApvFmQPMmRmNbHVru8O0yjRGZE+cheokI/zPkwuXB4j4Pj/2Uifx
ZEs3xE2EA11gaAASoO1EC9cRiT4suKTj238uVnph7gKFhY8YGjDZtuU3Cj3ewikO
TjyPBXF65ipoPYfP4U8MT5maNUIfrl770JkzGP3ialz1So7YV4Hj4JePrfJhUwVX
9nByC0fNJ4K4SrSjq+dhOmBcwW1I41TnnjBlR/th27nfF87B2SS7wphsEoshMVZT
oxFkMNtLR25+4RcfQ+ekQdmuszHV0F2ZJk0Qh1p+gXItjcd95ZBjJwLzN6WkB6vH
iHr9KC9HMn8YynJW+p23AArSCvDin8p6ETSnUBUhj+Mbpa0Uq74Icss2q4HVmz1S
UL3ZHiYnARgZ8cU2ensefsB8iezjbIGDfNwAdTooQX+KY1DRgcghSX07DlIcCaeG
3vxQXbyyqdHWsEduDM2QvORJ8H+uctheqaqCYJyGCsYCj7FjYcX3WUuJLG3oj4qh
solrSTrs6W790nK9+ai5mn/vMOx/oKZq7raPNw2j08lLB+ovlVD/67DlE8VZ/PBo
EsIFOtiwDDdMuh4SbWwazrwvVIXMwgwXtPfGNAd9ehhWYjpk/TGgHdA/ZPiJFued
LmNtj54wd3eCDAajJd+CcgyFae9tH+DJwZeZTQMdFMexNzlaEpzFc/j/VcCelSiZ
KeoTuOzMqM0eTf+ISMxVCI7qLfPhL0WRSJjcJqINbsntLTDUO8wn7ZLm1T1qd6y1
3iXP+tq1q/QwVrT+fWn33yqqXyLs36NzFwsutJ1vjqhyx1o+FPV2CcCNHio5GPY+
Y+xqZTeDcI0cha0qIBXjVm8YazF7O9csy3daNrAaUbFZBw1xMMau2ApJghS1H/ld
TKWLC+tkCeNP6Q1w2tmBbOYH7vs19CTkWKHsQV6kOI3/ysTmspzgpVxGTcX/N9BC
DVclikOC69Cb3BJJCWfGEvBrNOAIeLuMngvZun7O3dXXZkyQeAWQNW2w+WBUhdEp
DxXgH+ubJB0AtWEf0EEO94EzKEvtjisYtkuzUjobQEk9F65/7G5CtE+79QhNigP5
mqH0aPx8aKdPXluQIx5AVCINifwftz22v8FPTjxDyy1vUdbdvWuiZzVMxAe3AITR
Cq1BkckXagAmVbqujRzkusezrrP7TDyMxUjtFFbm7YbrEsUaGnBM1B8U7Ic1z8nr
E/EV1wULz3muZzRl75NjP8hmRZrz59yD60C8gKz0XQ55PVw7AGRaRfDYFo61GDkm
wJhpupOafmYz02qQUB03pv7Bzu61WIWsffX+EhIsBV6Wh/LAk8ueOGh6s/1eaFUx
oHhGSr4WI97WI4LO5AfCJ6DRDvkNWsIT60TXvG6CNCYtDfOnSQhBv5JfglCQHISq
6Uh0YZkM2fxyL+aiAbZxJQQ4AbBqa/fCD43SKfq1EofppbRRD1Dzni4UyIwKX3TM
NbAQS85gbm2XAzUsT567qGohUU3EYV8ygWVtE202yN/XrSMXfp3q5EZGJNzR62YX
EHqHMKCVGKHzYqoT0QRYaVTRSWga5+TNinodi+OtAy4LEq0QWFfkYCOIOREab/ce
xv8e8YiTpmNz9JHywE4p2RttUlEXurnkaRCevT6j32yk3QlJxG9Vd4elQBN/Nt75
8t2Wuw8RgNAMcg1cxMQ0+7xWfkaYxwMlA2H8FPYBpozG69xQu287oa32wvfKmqXg
oN9M1lJCrt6RuvBbet+nV5yiu4tPnKr3krQqCUvpcLh6aH6DoXirX2770kHLR+fj
94HJ00H+gWCbNXY4m9g5s++KAgCCnx8v03BSbgnwX80cSUt6UQ/7rBtOrBtoY0Y4
LIGmCqeYssvUpME1COkf8MhBMok0XNg2vx7fXxSXgaIcbpqB0jWf2R402vK6tSun
4RqUttJGxi0kPePIZbZU4DSiwkrU5wzHR1DOfiu1Y6wBcSN3KSpUZ/RnEx7OyHvu
CFQBe4tp27wbnfUhnaIEjSXcAxyiFrxCjwHUQgnPMBjt0Y1nFuQhwflaBRYKwpjl
qsvjqOsYovh0WZPvIc4DsE5vbf09y2iSPFHSGMwfLGRHzE3RVVxXy5KrjaMHHYiK
NvymoumrB9eX5a5zh6mJi3kIsLL15dtg78Xgwrd0oezhs06Y1bcmAeF6K75qW+DT
199oHfcl9awqLQ3757jLM9CNkvJqMBmMXCeu/pYDsWGhrWC4BhJhPm17N3SOeSHs
QDRvo2J4r/GRoiCBjzQLr3b3sTtYYKQhSAaN1a+86ICp+zIDl5x9D65DMaZHm8sW
AbEZDBKjRBrMK5cHYPVvV58jf4p3T52MS3L16Y5M3wZw8kSivPVtHjuzhfIa61R+
FUQkkMYrD1XfhPljURyGQcgsb0GnaeHT1mm3uTWFc6qHeuDwICr2ekfeatI9LyT+
JWpdSMjR9/44Akq3pLELG8EzX07aJlDGHqbeMwTXyEmj1n66rB7S/V9sYT5Vep6T
p9vW12t3t/kMy9W+BIvSnlFWiV6xy8XXoCL5GpoQ94d6iaXKfLDoSG3iiqeGpUNU
IlkQuOtUTnO6QQh1WC1Y/ERxPtQyC57m9OmW9Rq6jB+WJCFgL30wjue5KqzwaCtx
RZTGTVBls4QRecea1yUJ2VAl3OFjz1jDO8+JKlakLKWNtSTazA9OtXKJSElcF7FK
RkE5HFK+YI6HlanCiBdckQT92pib+//xDuZeQhgDZiDQp/I+r7HKUFOeqXLsYGYz
DBcBVXrFB5VL+F5TwvojumEn02ougO2A9QqzyZ6AnJowyGTTqFHczuGikmo2fPXE
eN45Y/Hle5px0vrax+kdhhhNVS2dDtgxXarJsHNpYKXjRr2wLQkpKhGYkhShY/ft
09YELJov2IDZzWHBT03RkfLbA3HoOas6wGOLUk/lfNbuqYWBifu69U8d0M1v/s3B
GL81ocsgEeF8q0pnGQLUAzozFvVEENsSD+mZ2SHR4RoRltmoaE7j8yowsAuWJc1d
gJCMbOM/uA6OqRbL2IA1zkFH45OTfOQ9LaUTzrTesCqNsnIr4qjjgwZQESjjxQfI
dSE/14vx5u963y6ODyqbn3/w9osyMDkXp/K+XZtxJ3gq70WUE0eBu0n2Uy5Ne9BE
fYPvYn2QXnlwg2qcV58xIgV47VwKfCHPwM7HlJe3YWBnoIXe45vLXqV5ubLF0Sik
wUshMjmP3hl9NlwBqrhTLEVNytf03h5XgyhPwA4x2OXtvdX0DCN1aDHL+LERKcrh
1uzRSI2TRTJ5ATeMAw4GYWNG6j3WvQ0sGD2FyEm9JSQU5eN3zRjID8IquROIGU62
WQlenUusKqNLQFXP2Tn5v1yt/3AyhqMoREJKuFQDJX36IwewHl6Bw9ysX80jTJ0W
lOH2vLzZlyI0kCIMDtihkhjb4OOlJsnKvXn/kh7y1u36TmMiMH7XE6OvQYe8igg0
8fnqsMD+G0UeXEZZ6y1m5BJyVP/LhobPi+8CP8pHHh6Dawtv47dz1ufOUHA6PpdR
vMQKr+g+AP2gQyKxhQ6bcIz8obUni1PFUs4rhhHGKuhozFv/JBD8MMHLCvkNVtJ8
BSBti0VvG3IwFjRCoC8l282x11Kn64tVWFr6QtJ3G2vhPSlprWrwJ5cp/U4ipq3b
gnPMDMb8r2BVUIr9LMYvCFDAZYMGRKijAertkUz9IKsL6XhRAHWH5jeHUtjmT9lB
yUB4qQ/JK4p+45ZSkeKvhCEiSNbsMKDjQg34dovFx3zACDne5E1jLqPf7DWL5uKT
7KHY6oOk4txRQFXRYDVKKsAzTqUmR3xdiKI2eIBv+6E9WfxMTn6OSIe8devGhimR
y57E5tEDfEqi2HfyUfvWH0TqpmvV0TmCqktxv6mFGeuvbFvrYWoO4vQchGkggSO3
dSbreQE+/r/xZovei+qSXkocvDCEzvqbuobDLawNNS4aIfia3Cd8SxdCXNarf4U/
MpwVRGep3LDQhJTCnaTFXP257yZfQn4Z9ny2lzh3w+3r5DZ+pPO4TLriYlqjWLvn
/5QdxSFyN/V553vS7m7863n0bnyMyZsQty4tVIpvW4EC8HFT0ERxS3XwfTnAZ5Pf
4Bx1IoYngeiZ2pew8hzVQtx2LWgn+sAljZh0t7yJrmUA9cIfo44G0S00P9mACuRP
3+wYGnVjMbUGY+tHfMiNFJDwKGPWvfUvNzIiCgqISp/tcW2PZ2wCmzn6GvZyeF6L
85M7vQinLFhBSYpZtLAwgXmsgVzwYuQWVq60hXQzIYeX9T++o/lhywIrHjcY+zZJ
y3eL9dxaMEfF+Dkr2weYQhCMaPTZHYnNCA7ww1UzS3yoI1UrCz2Sg5tf741XgpHq
MfpnGkZD3s386wIfrl5BK4bJie4JGQDnLy0zZfcC6DUnMJ9TZeE+GkNJBWzt1UIv
ANBgX0iZs+P7r/XwFrcihU3C+RS140jl4VTYwNxPkgrppRSSh6v7qcVzqgHjumFU
MYRJVjARVMX/PB/uq2MFGoz//SkJaQCazgDDd9mz9afzNBd3yIcDKHPipgmhPq+P
8nLDIRqStwbRNX4d+6XalYzPLlyLxIUXxR5+8Lz6oSNc8ntvPVG0tB4u1XjRM1HQ
Vj6j8rIJEMKN3C+4f6BN+HAYYhRJz0yrF6vS9ZJD0LENa3cjRcL7QQHSENp9Etht
w2OkkVbO/ENKT3RT4RQgRFJi0zN2fUqAJdR2PmVaNOirikWf6RWvp0QQTn3ELgIz
WcZ1g0F33ModrRDWkzfCSBqPhm6bcz2xcbLjmCRmkfEoHIMuX+BvMzM01h2bwqoC
5mFCUsJRoMVBJhhzp5N6hDmKFzHSv3HQ+/L8X5uUsaYsb3e+RA0Lubw4H3SrRi4h
Lc0giqqF5PcZgnpBPD/LZ8SDI76YbEeQTEFlQ9t+99aGpknycaOspvhQni9RDhtS
SAPV6bDkMaG7k6Fo88mJA4wI7wWZOsxvXeYDYIeOiq8vPaqArOXOX6w2NZxEmXBi
DpoGXIXH/beeZ4cTwu/VyWRjyEg0LCWYS0reXpK775B3bKQRi68JcMtpGxBjstOG
LSogIsF4Ddlq4+Hx46eoMYCn44lgg3+50g1l8Zs4xS9n0IJNHGFuBVZimlxZb9US
FEZFGN58w7EGL4fKqIZysY87DXwGhF+ShZwdZklWFQYEG/0kxvoMWdzyEZBFkyPc
JnaCKH9wpRjZcnvpgKJmEy+yG2MVWvGnYbJ8BL9/q0S1Giir00xa9Q5AYoYHEVTG
lnmy6+mKBzvp4yzJMLEI04WmzHknun1P4SAaK/sxObOZHiSx5THfyj3v5Pnia5Wp
o9MmyFQR8erC9Smv0QzUH4qw7pzugq5TkyNjaHvXO9HAM74Temnu503sAFc5xj6u
G3wFf6gClQy6b0Aot0lqD8Ve7U6HyHvTOzBbB2Rqdzll0KfdOxGWmWaEzvo+fyxb
Cr468DgA4ZpEOsxSDioUAAbdTEsVVilO9vRXGR2mCa6cycWUXspgXk/RUGftDs1e
ukPVso++HGrVY2m5ErE2oH04XJ4DJhLtq+9IvRBvDeSStda3D1RWkFVh68c2xayz
B635ETd7MLlL6KFIWtvE5HxX6hPhCawnZnNAGPmVkotYGfF8+PL5KJEwyn/MkRRZ
y3h4TtQOKQ83YUGaFoMTy33OPRnfbPu0oDw6j1CLF6IWb8rLXjL835iXpMua61+v
ksPcwOVgPkICsszV49N/r8ETYmfDOmKTQukcjHz0oVxDoa3GGCnk5VPrnJmE2XAk
vQmm3GqEO4cOWV4U+OJLNL5Rv7tdWWk/ygjU5NlOKUGQEiR8vLxAvvkg97OE2q7x
9723Hy0ZvTupGG2ao78/yJM4DVbvj9nfM0V8ooylxXhMgv7FOrRfbOR2yvZPVw47
yC4DdiJU4+dDGW+3N+I9kdgC3JIXHnLDqo57T4x/yX+Q/bVsSBh0HnxGAWkA9nTi
QuIgTB8hAMwq9KOYqeJcTS87BuEYmG8hdrohMhx2Hb2OHKkNMnR95UBhyQbJLl0m
Y4vZ4Lv4EEqmBEnH6L6V/mMWboMTRBa+WsqyCwKVEpECDTYnj95dg0dEQ2NdhW4c
IjC5EtjglxLlc+5LxvkIDbYEtNp1jEAoPmsYKUANjK6KH+sQY6Xz53bGuqzsCSDX
Z3RKazIN31sYJKmMq++u66qGlly+I6lpdds3cJNzbLmFI9DNxWrf//WYSfsnEqD6
k8NzXFdnVEt2Nerruv1xEO962az/oVrA6kaHRITDZ0+4rE7bHocDDFZiFtn5moQ9
2oRtLRcyOyZm74jOL+8/y1Xjc2UPrvRtIWL+pmqpIZH6UETuHuWqRmV9hElX6E4Y
W9NQRUez/yI7u1xHrnghniB+zElKWvnGZqnudD8M6w4X3340Sop6KOzf7FSHRetv
IcZytWFq7sVX2z8NPzVf5XV/WrEeVb2dmaEzJ8dj5yPXvfVczznl9PRh7baGM0Zh
/OYwZiyj4AUGk5yE+ZyohGdFVRL8uWzlRYHOdQGfknwEkZNFkAzXnvTwe70iqEEV
nM3hdscuuvbyMtkO5xg5gGi55TBg2Knnzq/EfJ/fdSM0/QeZsov+ry6e/JXBXm3S
oJ6igC/elaGHwtZZdxqYSRrbaQvOK5GJxhQDsyOKdeqXTTNGol8JaqqXFGK0qSPW
kbY28nho5nuBug/Dk5ifnv/i3XLl/FJ5fv7JpZKu9GvRCJ82tPnPexIgUtc9e0bv
Cva3bR7JDNjcc1jBMvARrF+azkbSm2UNmusMigzTX3TjqDOI/7DMjL1s01xXY0Dw
p/ToWAEjX76hLatmu012TO+eJxFeleDj0OhUTfKyWuqwNRCO/3jJfW6PTDOrCUJ3
viV/a4IJ0t59nYd+8azznREbMPs0GCme6mxDpsr/bmxec5MIUUNggnk+fLgdf9Nl
rQMPCLZoIRlRAAVq0sxawWRnEgqvMfedqgWben5+Vzq37G+Bu5x/pemVFx6JXrlJ
QyVmQgpkrV+ys1B4JutDtCqUgO/1xoD7sLdbT3nfFk5q4HcXhY8Gsh6pDGjPUadG
7cSBxl0su4pEA1FMHROl1Q+hLuE9wGrXICK/J1+gF3DRl9t+4Cj8X7+w97fPeDv6
Lk0uItiLT4infgGeWqwKLoFk20lk96gGJSUNO7J4q1UnSp1CvjxJo64nOrD3hh8X
/h6te9622NuUIqXEf3/KWUG+NzYj6ijDH7x0QG5kZVZcWQ6TtgZ9VJ25ZNtz4K81
U4eB0lkTt959pOYQOFp/QG71FbKavOmX0ws0fYYXaRtHpGGfcCxWs4mc8ErK8eU6
215NpTDg5iilFkkFOnjazX/ndYfhwcMoK5qKosckii2CtdRX7rM77W21BJF8FAXX
rTHG25zKF4b/3VW5mXHK7mj9MmGiBey9RoEAKLlLu04rDQ/4oUQ5459C4m+aNm9S
UkEZRasoC7YEBTZhNBNH9N4P2ZAYAVN1HARmxBrKSZT4Xf3GBTgzt9XFNNxM/b0w
0lnPqXeM5NsWXT8UMdmJ3g9FM9DcbZcIuawSjI90IQg6k0F8hpPOjyNtTlUvTI4A
nIIKesENJIJyhHbfcOxtNvRqc06HQJ7Fz78ktRCegtEkpXlu5eMSwPZHCtHOiId4
noUDjz2LqJNw6UkUwwjly5W6Mf73pCFRgSN+ZsYTsQBxAckesA+z00qGlBjhiQ9A
bi7OD+zsUFA7GUT63swKS0GRHrbLLRBbbaTyNE29XwBl9R924z5O06PBKh8TUlMc
yOTcBaf7lRz4qr9aPcZFtPg7/8wYF8IKJPC0csKVddisPXMhzlMoHSnjCdU2EJhK
O/pus4cCANwVwxa/UdDpBp1qfse8cZiLALobL7nMn3cgwn65V1G0qjtcmvTzx221
NCSdCZxqBmQmhXoomrtq/7/p4/rRZJQ2YOz2Sg+HHP8sg2ZJZCbM3Vc0BN0hOPl7
XzvUnCMUcuYXFHxFM59tYDItir6wCrntO25WsSyFHr6STnSNdl2c02tbgDTb5AQI
HSjA7dNT8CZ352uFOTR+0MghnLfL/ksTIc1Cht+irl0kXqHLuGaSP1yLIUwBwuj/
qTaiBEIjh/MleeBtQ2obo/QvYkKNf5Dw3bIj4uQ8LgVSicbua7I3gjbKk0ca+Cay
rY4pPpkfPrD8vj7M16UOug/9GEopV0UOxCYur3sen8rNYxfNr/8DMWUiA9N5fLhD
O8e8s5qNT0yj2p+ZjnXQtut7N7LigNmX0nUoqjga58jab+zt1rHGmm9Ro2Rqbb84
nyHkkxHAjWF/Aq9nSYmPVxvhxrIAtQSZm5YtRupzfAl1N41KgJ0xtQWSOJqcjLyr
kL7VZl3FiE72XH7SxYKhHcDNqiYlJfIi5KvtRJqncm9UpdmZxDSVMFDRnNJ4W5BX
zb/Z7Q4KQLUsW7+wutJP1jiPSUv0mUO4fWXBBFOJOvK8xnYBBEyqw7PFgvveA1Z1
5OwnLfDDe/z9C3B/SY3gRkMeSJfeIemnKcH34HIOGzfbDCM73Qof5Ne2k6SYsKjP
w9jLOacWz2lrPnGd9C/4lPKP8hzmh6TRRP51q6RstkcBET/O6VE9tTSmax/kFIvY
Cl9zSYHcDC4+TXTavGCPLg9zMWT9xXe8SBjEtrTOToJ7vJjkIhmbppj3C6I5ukQB
I4XiaWOWKdasWUfyGmyiMRPOyAGXtEy/XtevyEWzuzrxxYbR6XnBzNdAi9osj7Vm
G+rwxEMZLx9V0Bwsp8U9ImxlHYZk9PYYsxpSuMk88clKRknG1GcaSF6eDVDgdLKU
5/HVfIT2wXxNikksGMWyiistp7Zb9aSlanb7qBUuRqtaylqC5R26ox4V4D6pcu9Y
6D1Ci2wKQQFdoyaHM3QXTyeL3ZcWV48AqHhXBRnbQCqpaAFczEtXyUzvehO7F12k
JEpVejO0JnNDi0EliC0f78fv+9RgxYZXGwHgR1qb8s84pC03XtC7S6L9gZd6rGaQ
cFJjv+nTJFiNszIOOhJIr4XseZHda2vM4RxYsfNANIQg7jYa/OcZptbtwMhKaoA5
H4CegX6MOpIR4DjKs9dC+8NC+5VcKxt/AcbgpdUJD/VDlN5wvfGaIq6Yz8Mao/UU
H6pBCPZnJcJPLPZ1z3Ycx5uXUuwQVyjsJAZFM2yVmIBfHwrVcf5JhzMcDG9ZRBD7
cchxKM5j1+JD57LOz9jrFgFNF+rQymSUgZWx6zxfqDtDPeQlIAVT2c9/FhApFgJl
ib3XXIpFl/6p4VAbHYHxqp2nScgRl6bExqxKjQpOJwXM/LZnFctLWeA/PRtOzgWM
Bmi564MzDoufPCKeurG7IU2nrtziZviCLp8SAAxASi/AgfdPOWyuDgzD/K6gzcyO
Z3YRgSsf+PaPZYFQ1EjBY9RaRpl8r5CwyuWiPmAZRHkwGselSj4R1gP7oj+b4ltO
Uza+G69XPpRCeO7bCuYA2ywRyqremu3EaXALpp8IIq1IUw+LQ33eotJtZ3Ii1l8/
lRgLGZ11DeSvwos8rrkTDdp7ly8dLXTqVWwqMI9euPu6fewb5TUpr1dzE90PSUgt
SIRaL0qAMLYN9kTJWVMWeg9tDnIq7wfv+eBV+xhCDtAwCLQKyqQOGCvEp7ICudO1
ynzQ+x0+UmbyyxTAFKFjwalRkj/Y5Y07nzzrpUX9626pwVqyqk/H+Vl19LFh/WUj
j/K4Yds3rPsN590yuPelkhTtPugQihEyIHtEzqxwH/mOnEwZPWFRmOc4YFfN+oSN
SKLSi4ykOgSOKwZ1O9PdofZb7mdqIHb+rIlRm6LggKBE7fqDfRH/Zos7LusNZ7yg
BdXCy2hBj6JkPmmea/0VC5XyM0DiKr91L1XYNo+1hbBzt8aiTDhhSY/WpdyNwbYl
KuiWO0xqv1xdfndUcQEdmrk5jio/lzlqE7pRwuTxeU7/t9iHth3QYqroeC/kwFaQ
Nq3moS4/dqmebwZ11MYOmygDf8Y552Jx9mBHob3guQuXEgfYfTClU2WFYZbJaeBL
c9b3iK7YgsRj+zNEsJkXAToB0zBuJx+dMZHhF+9t/u8oH1YuQPotB86et/jpE04f
gfiASJBht+incdhNWNlEs3Qt6DSyMkI9GyqkLqVRVZWHLfsPOBRO+PaFptPwBpK7
iqZTY3ONi/8v3sON6EMGdG+ng3CxnSpptwYqhYoYXvUjvlTWq14TZDcbKoMhOytY
ohba3QDGKyH+XnuH7s9L+cT1d//gDAUosUfN4GfaSwelCSHPl9RTno+HulvCG/3Z
8EX+4poausm+Xi3M9YE3rRgg5yDlBJv2YuzLVZ+C21g2G/V9tZJEVDxnfSeBoGPp
j4j8n8X1o6iiSzgE0FuysV6ITvlZQizSybDIcJsk+jJrp0HU1cytPDWkgRMLrAml
fGAa9FXZ1kBkpWKdWeKI8EYWDGUeWM0jecQTCcy+GHwfTiE0D4EAWqf4XJsekLxj
gMQ1V2vqYYFO8R4yKtD2IDVabOURnpyWkwuIp1oQVKOmFsy39s7X/DfHm1tWYc88
GJy43li+9gnBn0ywQqxcvsJ/MQ0IZpS0MZpyU+6N29ZTo7/Ds+zejiVwP3AHpPDO
q/6yWiZsYVoAx2HBes2Tp3XvvVnyRKvGY9GPT0V7aix+eX+QT4otfvFBYQpDyF3w
8Qe12v+6MK+OsgbQymQ4kqYTyNK7Fk427KnFA2g+TEsRIzGFPqm7WudoM3E8HWi6
LmmhY/13Mk0L5axP8Dblnvfd5wLRu6FMxENIMZMHsTYuk2TXqD3WiAFZD4hP9CvZ
JQcCq5EgXOR3ktLGV9995vCYfLN9kziZK1bKzSu0l/C0Lf+OfgpAjXyItstWpNZA
V/k9RNEs7kBdM+IN4+EUMDt4rdMBD8yndSe/NdRvIC4lkyKCpg+unMsqvxS69XZl
9NBPfk1PNT3V4keXbN3tp/jf8JyesYptiPYzP6XB2y3zBpneRxV1MAUdrGkuAQyv
mQO3pU7VW4WNZNbO7mvIwy6XexLWd56Oq0htmaMYnoPVccEGOUi7tV0dGUWlG+mm
awMr6EyziQ3oUDJf19mMcuxycKNW/Y2dR3VbP2qOjS3SIcWPqr0pBlgqoXtRMroX
TN77S4Salhc5/dxuy8AP7lTVrfYMcvm/7pU98Exn4EzDM2Miuo3m1rXAhFUQ4kPk
E9eXkYH+0PQqQN/8vj5eyxBoCIO35vVPRk3Bvl/ALrl6m7pufmNWM7sHztagQH2B
qMDvNUoWE288AGrCCcvCd3eXopmp+xNwsWeStkP9IrCoKjXE2Ws6JcrKMYD58/9M
ve8pSH7UOBvs+Y8HeKgfdVnfdI2yYrZHiqga3/28bR6XSbo/3ayzB/HduOWaU2n+
AvIymN0AI2peclEMOarWPX9uGf9d22A5d2GYvT8OIDzCXnuOTE9n0eVv/U4Q77Um
gzeBoBniVy/1MjRoIAMlOhJ72sBVC/SNI9hu5AfqOVndLLQiWAyss5hqHT5fZ/+N
Doce6TCrh+OfxqxVDmEAGjHwHfmjnfm7vjY6RzNLhPQAG5vtmuTLrA+lsHjrq64G
DHnTxjPFC2FoQGdbN3AbA4Jp1gmYSL6V9zJwLADz+29eHmKhe+3lEdHa/wb02Q9r
x0y9mKhSCFqggAIbSanLmbXzKmkv7hM+A9g8V+5Y6u4Q2x6c1QMwTj9n6MlDlld5
C4is3rinJ1L07A7n7DRz0TbTdTTFxLYzAFV+hWKTz5LrhwGwv6UXb3oD1YTf25I/
fbRl12RFteoZ0zBYNVV3FFNpVdmIAGaZNQNj/WLf7n4QtGfSnHhSfe5i2fg+OHej
Oe970X1SvMVT9f9k1bU9+/rMxqvArz9Hx/uynonb002pEO5AcRYTcXy8upjiMc01
txhXK1u2ax4WFAZA7QOUV9IqRMI38LgZmcsMxXw44JD9kH9a7rsTsAytV8Tnwav8
7aRxXWFXBfLhq8NaxaVQ8xYLgINrX9O7wZ4M1FLIOMv7c52Wc89M0jnjK6U3IWvh
g2eZHtIeODvAgvPjShI5Ix+yxOSvH6Rrjs7acuvjT7I0+9AwjnRQke1J+tSMNYqt
jLvOe1a/65DninVO9FGQhgCsvvo3OwP90mDlIGdRwCzKB0GnealpywBURTph6qa9
/7AHMhY9rrq3EKElFRZnWFnNwF0gEsZ9NIFHlUyL8uRjSpNCnjcQ0NquNtLpfeTQ
5UfHV8Q7EjSAZDJbeb+gKG3Yvv7tT0q4EJ7SdgycctT9LggMG4ade5JkZhX1705l
t9lUossvbZziwrZTM8yGfkJ7VT1t7HmlyTKLjcffvIkpD1r/+YTkYQItlEVqZhSN
7OeeLQUmlJXEsOYRnkE+VDv6td+JSyMQjNEY7Vb68e1BrMWSAnzKVZcu9QmUrmdS
V0ObkbimCiQ4cM+KN8FWDYnf2uiuLTUm5j3CJWU+YKiimCWtiuh32s7/NHmvnla8
v00AgbUyzXwkb412cwMk14OkK6hL6aFWvPQOh6y/KppQVOoW34qBAHDCr8h07aEl
RKB3wEMYQfeUlr4jbV3CroacUWOBGkzVB077quyRH/LBPbzBSntlXJUafoEnIxM2
Qw2XhPdn7eJgJ93vdIObUYRd6aDpUXk0SLt8g3yYwsVDuZaqaLwiLhKxZXzPktLt
lBZEyL2dr5P8gJme+YEG8QNY/G+Y90KasZh/0FqZMb4R/FLNRycTNkEzWdwhenEo
aNrrERUp+IZN8OV4wmS7SUtNFvNYuLgjOKqDTRbsGa6es0LGLgO48ohjtF2IIt1G
Zinjau+rHTUNWFKgjVRaW6r7UMU85Mf7p1G6meZqjmP96CPmDg7Mm6PTyPV2i0rJ
27SiPQhPAqfnNV0t1KUnXAx5ujbFFVwxwoegKNdPC3mVSFphPNVJI46MPujmIUbX
jZ1Rh+boLygE1ZybSrZS3+l9jKP5UQUtLOENs5lcyufu/OLWeAFuPxTbwnJe2FlK
i5ywHbNEhuaaqDdj3Gdb8OyM/GMQOkfdNtzEHALyPnUNnXoBa2U/AbQlUSETVjQu
lQqs4eKNvQALXbCZKonN3+U5o+oA5folk8xxqpg4n5neCpoQJWBKle61eX3TceoV
cCW+7IvlMg4KYFFrhrt2571nlaCkN2C9PgeqqFU9/U8Lf6jUYoUOtxSs34XbJR1W
BIDYDGT09Xyd0b7KGnoPic7EUhef+tR1Lps/LWf3/CPSPqk9RkqV7hnlxLdEl59K
mrhwbTpy+KareJAam3Wzrc6KOniVl78+hOLZrVwafbkC5ZriNx27hc0FKtkR9vbt
SJ4EBvRWHj006GN+guPF9BLFU0jF39NhMiXberxwn/d6T3+Hp/hXthHl4B8EmwfU
/ez9TTZSZdkSJiYy0RHJFXzbSzixXat2ulDca9MZmxK1Wjn+B1c3WLY80GUvD7SP
dDo7Bdrm9j+w2rNR8TJ7lRrUui2oNs6sWPTLPTROoOz+LpsZePj6mgEZlZrcpJKx
3jEYzaTiI7jDcgDEYHS4lZq0KVAWbSTyT4nY+n98eQGGC2a62ibfnCusDfwnGABN
ZqGDJ+Ev8Og+usOD2HElevIXc1Os2O1gIiyXPhw1+rDtjCWZUSICUNoz9+eDhVgJ
X7Ryl6PMkRcVVwu4paSwUd1T9DDBqnZ1MZ8VvgTHAeSDdJeVowzgIoSVPF9u+IOf
F4PUaoSbBweC6Z5HeKaZx1zZTIOchhQlEQ2Cp3EpRE2cDqJMKLrGTBSTsFx99MTB
cQ/tmk/8Dzq/VVdHPL0ME+dmSMwmlcAfBnKqFbQi4Uu34ICXBKaGsEelE1JV5ElM
wPKxAApTCrs0ZoBdkpPpNdOYezaeQLEyhJsU0BwluqxJH7MfQtDbt77+HsV4sjpy
hRTrUu+Ly8625g/9OfSO411ZTJVTAU3DqXurXgR+HRrr7wHz5GbfM7dZpcoa0k/s
+oHGdIXTbyhn5m7Hnh9vF8MuJYKz3no0m/CNHcSPmV7ygCPlIM7Go//XLvcJGfnU
ZDsc19+a9AJHCt10rDFseIuG95Iy7+3Q1beTC7y3+S73PX1IXzWblLxj9I2tkgU5
OPElVAnEby53rlToKlRkIOvAtbTOWYosYns0jGw5ILjBpO97BbafaskL1EIwEPZV
UThqcIqnXb8aUvCLztpzGxdp+3LQYTX4b8QAj7LvK/s4FV0u3J4SaszaYpMr41AJ
PgLamHbs3R8drQovvCnKqDG4oTw02EER3qlSE1PpOGXkX1kYWufKWRp7H+M0lyLa
cy5rQcfjhfoxK86gcxfR3L8v4Kwfyqh/JsNg/lUlGenmpyfXhu7l5bqC2rJDVDuX
qfgMiRJ1VsZGJcfjblf3zX2pmnWMdtMV4YB2uhgt7QxETvBFckTVInI/8cdi0arU
L0N+3NNSxzaZ8hIpjwCFdSpTRJ2zGKkYCkAjLwTy8yOxH5wImkRAX+mZIj9D845X
se3o4XmL+cSjrSS0c49ZBDKqxQuEo+O6o6szq+jO/nykGnuS4QPLeZqI2z52QkPT
H8JayiyvqPhXehWL7GyzD+IDx980BxewtFcpZE0X0NFDy+JWjVRDujL9SwRmU2dM
1hZ7BJVJtPozWAPX2wpZa08ItV4BYBMNc/MiEGSF0jongeJliWKx83Mzb7SXsqVK
xBXTG98QvUokUTdhj5BlvHx8s/I73YNOCbNHWqacawWUCnI5tQz4XXlLV7lzfRQe
UFARcZ6qlFeZPyZfT8UInC5MJTMbEKeeqkGUuvNV0r6x9rrfzZkRVEOKUwSIDMkz
oo77p0e9f4UucLtaDYK58lAqa3y72/iCCCiEYZVYbbZ6l2PwwVR0fuK7dGkTYyOz
WkjHJuYu4XaV7LVQWXjDX24O01L8aMYcQ+LBi2o/eGSDkZPdDI+GTD6fMOnDqDV3
Jb/hqHQ3UtXCyewH2CQ8I9befnc8S2A6rsLwe8ehVH4PG1GL2N8yhunB+MPWkxKF
t16xJBTHzhmWc5yeR0qjRl7IRdU4bZPK4Uv87jKVMc1lfZEmb2eg0vcwA/Eyu12J
+81XLD97JK+CQ9ftCWSDGpyFFT4/zTAaPlqEl7bS6eN9+NEInClb5pg9PeqfCzPb
lVDSScyGzAztoByHKl14JacPgGqeujGjRfjhKiwLR3CLAYXdujlA92lJ+efVaFyT
17uDLW0JWh7T1xcZmEzBtU3uAxiI5fgTQCKAXV7xcqTiE44XHyOiknsC67M4MPx2
ICC4q0IF5xy+24lYOADRhiLza5XeMsf3oq85m9XHyUhyfka1c0S7L7bR3zvXFaAg
m95q6kDq83+r37mjL89mCqMyrOFK3pvp3mORQqTtFekE0iwZ/fXjEjjsY6BratMU
zkvFShPtUrbQafSy1tGA6hsd89haPthk2lx9b+MnlWi3GcjOGHjS1iAAt6lWnKn2
cvm0ci3QB5VjWoL4ArW2IvoUeqGGMd+ZKSrNv/i3+vm3eles3J/u/j7ICcpX3yg+
MwtBgPc+FBMRaaeli5s4DniYZj2bcK9Kq2RMQU1QNQjnFi2/OwDGdAjj7UVnZx6O
KORNg3POsqYoMoezFyvkRFjeiEjmb11hdLQ91FSYxwWAjAtAx27ufu0+Y+n/v5Lj
J+f2v6iJBnzCcZ2wfSrfe9toGRdoZoPg3Y+DivvIkGgfwdOtEvtyf9D5FrJytcvn
x4vW0qFKmh0uhdKUDZf9itBs1v8t7fHqQVSUHG5mfvaN+HZ2S2OsI/e285rWGqaF
HTq4AQiE8mxhsfu2NbbytfRCswogLSITZpdTkXt345BDnzpm8pvpRUrwiaeRuk3g
3LtUDuGPtoXVLig3BNJcY4/hz6+Ysm4QHpGA/fkPwPmSzUYou590mzCViOcFNi+z
oiucB5PiAZwnkvwLK3en1tnruBLZIMHY5kgynj4AO+cdwoLnAPiK+lg8iZOPBuIo
QT48TqJ91DhMkPnxG5hypmYVX3qTNCvtcFXhZZ49T65ttva44hDIgtLiKm/ajQom
4q0jYqJ3gnXhjZ2jz/VPsIPn2j9MLgt//2P0w1FWZVAZ2CgIFmpyc259ClUsuEJ7
Ie8NsKhtr+ybXSg5jWxIivOvFfIi65Di/KclOJl75mSybKNGrkElq2cFjDUviaSl
NPM0DleE4jVdiH5UT5DGV21W+Y78EUQuAtIAUa6gfOmuTu03O/Ek4yXin8s7xTqm
LwplJpnzQPX3vrIRpNYGbCMf1+F8XstOOQDDfqQgt7yW8UFCxpNmXaf0TT0XuJx0
t3P77cBBjbZvdAwoZVG33wm9y1wxWG6tOcpnGzaXF1pT/aDu8/TW/0fw/14vp07W
FLISAkd56PfRWYjjmXqWqQAFQImBaTQnslp+6vLCyB3glUGhvAGXHxl47Wnv/FD7
ryTp0Q5MNHXaDk4Fh07/YX2YYw9KvVrfSsU/ZIl4n1xs6AyQWiFaxcQW/RwocsA8
z8wU7dd5ji6//ckf3K2b8ED6yPSRHqme0u9Kltfrybb+vteHJ86O14TbQQwbW+Cw
0wE5G54EesQmRUqvkJACy5NSXwdA0ABBm0slw6W+s4Klt+JPKqOUVMUknQEVyvsj
ub5QMkwU8x+z7vQXVQCJJjLMeaXKaGaHATVOp/qrcR64Xg00khAw+YMwfK9A0+t3
4FmcZobp+aqE9pXIzx59yfaIIs2Ow8e4v7yTtHLL8EB0kGg8ugvhuRM2XqLLurDb
ZY+ztegznAeojSKNW79SArBneJPHk5YulmW76AUpVnEtNM2c6Bg89WKqY0YTVTWm
+3NgrpmK/OrDNlV3pcalanpYP+Q3ogywpJ7Mk5OU3lgHe3o1tbKcqmz9pzamfZOi
dO1a3Fdhg99t6u17Kk/aW6CtN09MhAUAmQiW4Gkcrr7DtWaFhcijRBQOfzRrkyqa
DPLOoeMKF+VDQIcR7k82Uuhvq+p+xX1ZWO5XObxs/tKolizdR3YAa6UwQmc0FLLz
hTCUy1/RWMXPQLNnPD3b7/Iel8dY69Vn6MwEwxJD0ow315k1CzgYslL+MVgBoMW2
hsL2VX+Qka7eIWaGgPYvOyxKnOYU1GOsVbZwTJ8A+Gi3ZV9qUhBM0+eyTpRzRMaH
SeqsMo34fmMRb9FIA+9GmNKy9KdLGA04BEhG2t6DT6KXw66EMbum31XttsaziaGI
W3wRkKpIIgHkWmHqeHx30fwl8uLdKceXRtpGHfSWIGihT8R/VzvQjaCGf2gLWOqv
3Yc+bl/jO096gnZiCfX0p+VyQ+vaQdyFNuAWGxLD+w4KOcyTWQlvsguLXBK27fTV
mz0KjCqF5tMhs8KQV43g2645uY/d+iM+1oQk5EnBZwJIeZ9//64EJsN4YU+GuuHs
E52dzdAy6tAWZbMOlmos9DUF0uezEFiHTuVggPUyMU0MuNzlW6J9zWs/gX69SZw9
66agG08orGEzg2qAmIS5qxlI69avoyDIl1foypLD0Rd3reL4wWsdD+VcbIog9sVx
FjFJkwUvaPIN9nSHQC9i0cPPKc3hYSXpSTV++0/UdQp1/ScBWqiz31Sd+PwmNCwi
qIoYQnXScC+wj8I0BqZRjdPs/UY4iqtMntSuH5q5NKfu9pg/I7yi4sDJKeuCth3m
qp3IarHdDr4SQ8PjqNphyiQN70YlSLPCsFIo1FSFZkgLF8ICjgPiKynD0qEMqi3U
zr8/IZrLwvE2xBxR4gNska1fTY8+1ccS8ePiRelm5OcOrsmA0e2VoPK/4/YcCdbf
n4r+Brl1kDQKGELEFCjOFSUapLTjBFCZ7ZmphsuTe0uoKeu9lgHfL19yhAOj3wXI
PK4JTrz6AsORy7Mp970ag5ZDzAN3+PzUAMcAifU+tP0TtsUuwaeaOfb1o/JussLL
1ld5g+v0kz8jDj7mRKd3/fV8JyacUqfJOY5LIO9/HGzK/oyBSf3+uG70Umw/9i+e
eqqLMCzl7UIbMWJOO+lY/DWClW/lbi1xXuMJnqL7mSDm65BQ8XQVlM1CXYhf9Hxi
xhj1L3ojrDPNyzQy5vEPUy6hq3tY/hiUbtEpjV6K3EngbtAf7BKAEYdx1Po9OrUJ
Rl+l92fc2V9c2JD78XBMGGc3RYnQhcxLKQKWpC7/L2WhpO2e/pr7s2AhKs1XC0Z1
uoZgztzgaKZTKPkWJvL/iB9sx4i5C5p8/+09BHJGoay6CAJmLd4s44Wi4n1aqiUq
LSgsuS8pZq9cCAvrJeLGj+UqOxes88AEkLCwrr1r5z+9vuS8HOBm5jelRVRmwME/
ZGxWI3Zwtg0SKK9dqeQsk+ehHCgQ5yxRW5pOBo0goiV154ry2qrl0APkBrZXLpYw
ypNMZFvuYrEdhO6behVCdDxJx0grcTSxxa59sJ8jWAj23Ir8hy9wpxsscLbFKsoC
WdgS7iGCExepyeovH6IAYC0KMnbvJ/u4EPAEi863iF5V/0VwcYfpZRVhqXYj51FD
0U4oHncEzyJQeIoxDj+egXRHaX5oNJZGoAmdDwPatkWG/KIIR85SzOTlxnZuBLfd
S6Byw+WaJPXvt5/ow5XjOTawSRk3pMHqB6MEVQhysiOUgAHnKbAEHeS/ZRIr8b2T
+8oBBx2V4a8S8Ye8YsjYYurcUaXnvUc7t8fi0yajuI5mtMI5bKo0bkiUfm24d1nC
zouzf/ISRwr52PpPzOHaXkVFXWw4gw3af9jROO2cnVEmNAXO8Zx6WB+Ui4MIWvfr
UpCtwH+afXr9BtQN+2lFSTyDiJRjbGKO460nrIMPIqS6YlMcKUgWt0v/WHlO6SQ1
VVzKTFqzBwIkbiaAJ8OuqwmgcBOyHvjQES6IO/tsMl8b9MVHN572BeqATCCe8bEE
0NMA3CyMdrRAbMWTUY2vYWXwMTWPB0A0ikw2y00PdLSSJm/AdD5B8HN4cv1NBeRN
JolQ8C/FUaLUpVD0wit7Gy/fKlrZsZqnJxIgEddl0QGrCGqg3uhlvWUK8F+7LSnl
J1SWua4UUz1mXlajyfhd9ssfjdfWSMcfucRcUxDWW0BYGsv3cfy9QEZpv738xFko
ciuE7yM5PR5d4d3lnzyNTxqA2ca6VY5aIeNGbe+oGxDlM8TtNWad0dV49m4PbGBJ
BPSogDtdqlQ+wr8jJc/KgwMfslqmtfjU0WHNFSSc0TmmMW/lOH5fpBzsDsLJUX3z
7fRzNYmaXcR8ki/gmht9oSwLypL9QvSrdWY5fEQbeQpTTo3dB0P8mZnUycKrdZ/d
UZ7NboZNOJVgK+3Po8PfogNJw+4txWzQh2CSFSa5+0wvApy4bxF5dx1mJVfKc6vB
nE0iO3rf2cWa7pWx8zN5UwFh8cdZtDa6r0/IzvbwLDFEH7zxqEb1nn8uRmSMsl8b
IslhfKMLabOvaz9L/Ubdt21NhwJWR1hqM+JrrxHOHtWRUtgCuF6TFhvF7ik9QIkh
GQPV4yH051pC7CLyU0X//7XG/HprGtjhZw0H6TC1E2w1wIrHkWLg5pjA7wHn4L1G
WM5AEvm6zioa9xZXrfIPkNeTnZfrriqin/ZYnI6dF22USj0wxFkrqnvdw8WHH0ra
FiiJhrsjJbySG+XgxDUZRRJZE497D+hEtF/J2BNlr8t2IbMGD83UWPBmoIgYqqfE
UgoncnPRYt3i2Iki6D91T4WQY289GcmrumdtOegSDCUvXAOxdgROSlR3dIq3yiDt
R4pA0NuLBrg5EjgseTPLTuXIDeH5c67HYFp+8IlGxZL0LXksbtms5/j3rWkBN9FO
2ujAHlRziwYYidMoGwDAGymvwGo9RMkzQwfJGAySiFI6ZvWNKf9n39rJt0Kk7bnt
dhTTipTT/rxa9BrHIngH1E1RHL1ir8uyN53O72IeuOI/B/A53jFdtlho87czIZFI
fkjqvFIvcSgEw1TUEXGfzH3ySvB5RU+MpYFGXL6t0zYmkHZ/gW6ygrEfU/PAiKn+
xlu2WbPcxL7+EzpQ5C46I135VQJUlk6e2tUuyBOCt0WfH9k7zhV63CFUSRkpNJQx
UqKX0Uu1ff8z+dElifXeSu/9bb0gdwSrZu4JfjC2GqE9OFeR/tVGO5RuDwqymHmb
M7IRFdr7by2DZ2UgFi9eSXxiklD6JDKKtEhLfoGT1YCXVWxAqq4fN2+Ox0v7KQmo
Wz5PuexAEIBFka5VV1hVdQIgq/W65nV+4HWd8Yt82xMbvWE6fXGk8K66BQSKmOok
L1268Jys/gTDIJo8fsF+6D4Qah1Efh81o3cqM/BomYc1pFZ3gEkkNf0tocYNjSk6
TGmfNJcm+3cjdc/DzeCnMUvGUZDBHNefqTHmkvUGrshQnXNIMH1o5CysmY3/rvz+
h2ombU8J7pWIYOwItPrQVPtWyOwknuKyeEB84gQYLWgJyuUkZwOmH0kGuoml7vkE
bSrmDXrQIIowIqFKgxO/qlZrRkqr/cf2753ML53acYAu5gc4Fi/iNzb4ApY9wju9
kk8bGW4kTpAH3qovPPWdDNo8qSWRlWeghtGcK+M2iL+XPlP6OYdjCsBu0JRdptg1
7pzTEwZ/KjIw7GsQ9R51Inr9dD4aUPxDZN7RzdBwMO8h0J3+6WxnExdAVqvarXWi
mrOSruPAgmMiMd3VzGFqkhBdIj/FbTbUP8+z5Eu3rpANu2LT64koXIYBtvNwkIs7
Ap35cgM+OwXgBYG9wEazhSApdTsWth86Hh3qFmtxPFEn7kjsluAS0ytNEmYfLiNY
UcTLjNAy1TPHIlp/dw6bKAPC+wQVzfKlTVY4wHRhovm6H6jNEsoexlsIHjCAsLoa
lPPdPs5pkfc1l4H/DtnFBcj1t+mxbJRGgZfPfo5GHJH4JACo7ou3DPmtWZCyotR1
YWqN782OT036i1tazvg3z/xWOxi+5e+dlY82mkE7ygSwBb3Uh9pK6Fomwo93Alyt
ywKzf9B1gWLKIueGmuj8bly35M7ejiAjgrR6ty4xG2L6AGxfXlFXnMn/Y43w/55P
JSPHYen43LwweU/1bMn2QbTWOKDuEiPeF5ersXTF5P2enODrr1RMFKJyNVnkfI1W
ytjj6hnI0X7kfoS0RC0vDGI2pvUPeU2n27+2jScBhCMhRRzn5n0FjIRuJzpinI3N
2S1OQvDAT215SeHCz50CQP+dEyra4eB6dX4ncnhWIEzdNiVb+eNRis5Iipge0q3V
bHiwur03Y56pHQBYC08GbaJxE3KN8tdFgscdjBjD+6gKFoLiMgDs36H//lVFxy4y
uoqzrDVN/SjsD8T6k8uAwWwE+VplFHAMkzY1V53zv1at0QHx5GF5Y+MJf4nEwCQG
wqDszS93qymyVKJYg4qQv0vxpfVUF/3TnnURXU6YHpgF8XNgKn+Hy5qI3pN1xDet
bEZk7HKWujKSnh61ZdXnyQ4Y8Vv4YtNCx6dqQy31BufSlZkW3xIGOPQY/jhhcZuL
yggxEY1Cvq/e5TNQs8ifd9lJjI4WpcWBfXSCytDTv0I6S1SPiIKAtrtBR8apu0LE
/dhXJB0eTZ4d/+u/6RW+6TgsYwKakrLVqlqzXnbO4JTrzkERvmOUw09l6ma5RS6l
tDHzrX/dmHWe1wjYB7UEFO503B3Ck5w7asAb8p677knbP2IV+HurnrAkrxp99gdj
sMMQHMZLMKVojhfYnitTGS7UpfaSx/eOesNJtknfiZ7i1OtXI0P6HebINX+yuKQy
v3UnO3YpW9b4s0DTHMMKy8dTsStkFW0rms6YfZNXPZNAk0E6ObKlvH8PBtaC4tWK
P1FOJXiMM2ZtOp2IvzdYgCEAOknjNNzOqekbhkgMe6jgIQhR2eeRRWOUXTgfpKTc
w+0a0qho6GBIbj62SNxqfDB6q8jY/2PIGzLXSkUllWdfd4ygAuZh3f5hJ++s/z3U
8lcaVRooj26mVzkQAWYJ8bRP96pW2f6QnkfHM1wJ3CbY60afUQji5zJH+nGRNNMy
W8vl/ae9uPt736HLdBcQxhPw8J8gMqbWIt1IbRBhvamjvR6fLrWDtSdbdzk9ErVc
mkl4+YkoTkr4SqNz5FZfkZz19WTktgQb54jfDF5Z8X29W+l3rEuAjbc+NAzwei/x
Td4pyUIsxD5vtbB/dfOwwQ1QDTTpmvCRyDe1UsKh5nrjtBHtxxbyUFa8/31X87RD
8B9nfvcoDukRWPzBe7VCPWyyn6XwjIxyeR31DwIsrFJGW2nhZDOvhnLeQchAxrC0
1Gozo2qDXKC0XILps4V6z0YQHEBfoaNcppYI3HsSbW8icD+pTu3P+pFHeRKsIpAC
0dCTGs5ZlVUg+1feldsVxdlooix8VZ5MuFJcTingwVf/CPKNZsRDKHICFEuiIqEJ
dMTcxM89ZbKgRcCGrlXFL3aAXIIR/ATnyleqMkvXwHGNVh9T/A0yInb3tvTLNyuY
cT/IxeFS4lKf9Z7h4iRAOwcGyBubsn2bHiA9MxIoBZ6wedwkkLwcbraTAVPIkjsL
BgvMOfU761VW8D/LbC8WlUWIz9di9xFr5UOzg3x6AZGUrzoC2K/fyrtRGLS7J5bw
xtbyy+Iw/ZZfKdFJVWPY0Vp7HVgu0sSf2KIOSXJ2aozePbGV/FzFvOYJ1IXjEtpr
BXIa8aAYQaDdA37F0WVvZI/qnGawnjNue1hCSQyI62X2FOefNoQluN8CHJVKwfUz
cN2xOZVQ1TcbeMWXs3OAOyisR93Khtd9GUtgBcTRV8yzkPq1CZpH74FoVZ+0wPgg
9O6cVvj4IPN3AbLwxWzXAp3/2ei//4fP8KDtOj4WTpF09MFYFEQi5jAMd98siHv2
LWFkvagwBdf49sugzSBUKkBaz5JnlgMcLcFY46YSGXjpKjpgaoIemfTyjKhRkgNU
/Z5whpcfLESDh2wn1XjVkKTNIB/qB56mudrKeA7vs54royWSrbpuq7uFYyT/qhOI
Ww27nVbfnc9X100P+O46VvSaUsKcYVufImTnuDazh1ZnrPkEO0hxobQ2p7ApI7U1
XIYUTfGNGKx4beME+lVgRj+M74adbP/FRNlBjO/2RK408plmkswsUXHebaEtlJE5
qy5oRKiCwj/P/kP5wIFL1mlZAES2XzzQj+NCZdUqWlqq/KA1T2SWOfYnbbNWg/wd
1uxgG9PtwjOcp8UqX9nXX7gcUPTpG43KRE18jocrG8JbCA0gs9ECmQv5swUtS3ni
9saLhxXetKfcnMOODhcjaOT4FhcOYHeUE06kGdy3sdhKqRQ6BmRtI8CmzMmxJuAU
mh6AmtMJI7dm0Vjqz+jXKgg4tvvaSuBoL+NuTPQnpG07BSxsMAT7KuCNvqw5SvWJ
2B3cmhDNfb94W4ip9z5XIYgmhWfKFe6uTh8DRE6NeKDH7J41H6oePyqJMKt94bU2
b36XOSdj4lvULF9yvQDO18Y/Ay2tiHSrodOdqjPFkLBNR3vAvjW4z6GUnMHtau/X
SL1ABNWR5HF3E4IAPxr6fFmltlTjpPIwarJpqkfl9sMkqRNwgz/igNQi9JB4NIM7
pTOcevNQxx/3V8u//HAi/gLX/YgVFUoG4Pp/BYok6TeIvTt71MUCM9HJoCK762VW
VdOMofxDyu9LtX+9NTWs6rC4DHnhyz3RMSgZaYgscDOFU4K4j473spSgO3RIt+P0
7cqoMpeSwqibKog3RHuJoD21qq2EaWkf2F6n0UA3sdNO5yzqHbPgs4F+jKoJ0zUw
j55rQ7/UWJemRGlwaX3dwpKNzj+ddj6cntZDBndoQW/2tw+/XaosEmpgI5G85Du0
VsvUO2b7CrrmuhjRdrcrywBExz1m5p8Upt0Y5nlm82+PB+Ko/4DmjXeQbYNcqieK
C6QfG8Nr6iI4lyPTMmcLdHS4VukKRBlN6fzAPcdzMRtW+lKf7p4GZBDbiAFa7vdl
eakV7OVTeq8pjdSJHNzfHXyDEcQFGtmFEUSazFGoFbcVHCCfq70OXcqj5yoMtNGt
xpojuviadrStaPFuFQTPBOKH95oOx9GWjPXbcZzUqj2urC36L3AQH8PLYp09QEPF
IhWhNACCjvE9SHVIjYocGyde9Lf6OWkJXGR3lKiDrl3KHUOMVFAlCHRTqmFt0q1W
UWq8ruwfgjbdBzn+bAr8dPJOACRlATMhBbIsc6dp0ldJNcxCU7FTRxo0/7Kf61oD
R8lwEjafhmFKV8BtA2uCXir4ZGOirAwJ0rPUBhb8Qz8djDJ+jSjS+nGL5KcOx9/X
lrAs84CYYseW5zoWP2zJQtKopJQqFrvViByrMIuFrvGgePs9mI/AZG0gjF9EEi0p
K/QrqRfGFOb8blj3BA1VfdR4C+yl+lETB+QsvVEf9Py98l4+01BJTUnrwtk8D8fV
QQY/13l3s/qzQSdMVZm9HkX0+/8Nf3+0lTtsAt0Iu7hUwr14okPlylq7/az1j/qQ
PgaJYB+mMGwqssuozrQOzf0zHAebE4SBLTzVS2xk1ODYz1vvzFAefwaPvL27GZ8o
eD5FX9BX4UknWOSEDMFXhNSw0XoIWifyrkRlSFrbgUvXEobv6SNGl37JzCpsJJEV
Ah3XyvTXfarAlGgfbJo/abDLzf7mIa/BKCG8jbZBZnUOMYEZEodU1enlTbQNz+oP
WT7RkKBkx3R0RDUeh/ikuNMD5gTh4fBM2QcjrKFVEvjSlA630auwQ4PUC92O0wNg
F2qtn7rynCS/NmJRE8ox/0L4PJ+UO22v/tOqHlvqybpKLcTKIVubZw0LAMi/EOAu
R2fOdDKkhhLar6TTm25+XxoO/yUGPj1E1McmksBBFiV4j/oum5yyfJ5gO/W+0kIc
l+OZsBIEPjSv8mX+M9dPo+BqxXmx69sHaWGZKb2ENDD6y1fFb00vXfTW+c9A2jxv
hb+mCcjCf2RLnci+apZDag8dRbdyC7g5Fd3eBlYOMFvPTwytUMC0fIY0P3Hsmhe6
e21/t+lj9mWJvszkeZZn/SKXW3RaKzE04d5oPI8nmhJzC2YnXsmagvEZHlbEshrW
FeyzmTPCEPg3dhgwdaboCz1Mfgut4qsLOSMVXCUY0jZK4WhjpQsuu4vGhPOsXyI5
qPnf3HfwhTPy7eo4LnJMU/7HbZmp57pHHou8gskTz4phZV4C0dWpu3v9OjmtzuiY
FQrWNFyPCDOmwqpRQgYqsb68xQzVUYle8kKkO4zWc0tUKBtvFT8G3akLLUs+TYL7
NVkXCkpQy98Q/ODRvOqgqaU2rwDSduUUHd32tf6eqHzIJebvEa2pcUtHnenqLGdr
Te4Sef1M+YzkHl8EdcheSx9NX/FG6hGwcFHgYSJTbMUN964Q8C4f1g05j6v8Iju/
mlOqYol3D9N8bnVbY2B0sZYGgBwqgWdTeX9Dj0669IlbD+TIenJDBYNHx9E2WHA3
rLhLKUBs+HFQ+Fwhc+ohqsmUnoK6W2Oh5L1apB9iyzy+93duLHv6HzHln000RFS3
dtnCKcsuI7xYN4Lt547YTWKj3Qxr8otxOFX1lj+hoMR/ywR3ofB495ISE2ik2+/o
Np+kQpdQa/misDGQ+kBrNOpvgk8LQl00l7Z6H8HR46Pm+Npquy0iLRcLuu/7QIr7
L0moO1KFgHnSG8quBihRXar3fjShpiC5kFGvNd/JRL+0Ih7mKhx7Q0LwClet/olb
AdgubGulZCGip0yzYhinAZYqAbg9w9F6gFMJYStwhi2AmS698ppvtDL69yacMv2R
qpo7EMtZfxit8em69nyUbZsnxnfJoZ4ZBWsWa90mxTzDux4dH2WN8H9y6ChwoF5z
r3ddhOcCAhqitFSa1l3j5POIYLjQzE4DqZmL2E7ziCCN9W3lLcirqIHPJu3NgTTd
V71xDO9JHj2aQtbv5NKXCXdfR9slgrty52gOoF3GZe9PTTJjNnMLSYqmwh8lKdjV
oa7SObbzVUNa2PNjSvpfGfEdJSIUenjeH8KhE0m9RMmWQsmsmDNoA1pbvq+h0ATj
RERC5XzJbidJ5dXYx+KAVwWx+Y5CnWTPIkhF02qBrLEhxmkQ7Ul/VcldSVjsQa8S
bVcN/CxrfAq/I2cLB1tYRc959d2/Me0F2KnNHuxBPjn+psKU/qntbDofuesHPWpA
8z+u+NJfkKq1wfSaiFQjuHLUgR/UJErLJMFGB94YfT9XEHXeEFZfVR/IBME/yr6N
V0I1oBDuFBadszPZvZVXRxZdlbmUhGFSHuhy7RdXiJQbukJfbwEINpH/PWNqxkIp
XkT+pEvTEebopCNkWdy6Y528CakyLabfWcD8UsqDm/uwPb2mq+W7uSoNiYXqDbN/
JzDmvWeijwkBk86VmyBPl8RequWzqpEiREfthaV60oURJgBJZpTGJ2aSTWV4HIBI
pDG4pfTO6FxUVRX6tjsi6uw5PskiidzHiAVgLiGQIOwMxalwNv3GduCmW0+KQMVV
/HbYMRzi/YDH/KjENs82jmyceMvLG5Ts8ULCHjgD0OoTvAUsDDeHranu4bvRwv46
PyVW9GCM2Qiqg96smnTQJJ+0I9vzg+eOzuEsMTePc71snqy4YmeTYIcAW8509on2
75kdlcFCil5cxqbOfWsxjutLIJyGaAcYogOyi/SLmybo+2ODCpvutAy9uqn7+IlA
Pfalpj8u1XSUjrVx59oGKdbI+eA52qATjqpXKEYE/AF+1MwGa7cJPbqTVC4dHfNi
DgTEG6um0UZlw9RB7ePXwlYjsId2RxDh6DlOII3AfAzFdGVDFS9IW4EQe/EDbvvO
VlNsk6OETQMvz+v4EnXVEvI7+Kj6Q73wC6Uof5o3hDl7jPE5QMi8EgbO9LWaWzbb
w9ezK4jr9vUhxPQmIPtrJBK1rls/+F+DqHQTDw0HQxdG95zkQtpaSFkR1CzYZ3Ak
5HpQsUPnCnLw9Y2ZqBYcQDIkem1bNqMAPlpgnMr36TxOd29tgM+ldMayFR6UKB78
tKFHuNH+5O3/vFxL+ejiLWKn6x1yhA3gJxHMjsgnMAoW1p54xxFYykUkXLabBJd/
nM23Y76Ul2OeaZDn5LZ+eo3tsLf5qHu9Lp19KsqGJJ6f+NxjvCau96MdOZEERmJi
IAPU3br1jNSk5dm9UarmUBKFRHaA0GHAqbgavMrCpDby/uV/qFBEAJlx5H15PUwv
aVuxwbAK5gPUvdNzAe3tlGP56VGATYB7FCtgbpNMrb8xZZvJaLdlJXpcSwM1YJIg
ASmAuZbDtv0dBFi0Y4pQdCwaDg+JnfmaiXrTzTFdGmfkIi+XZCLu42re0hju2aCs
9YcmZCJ9KoukC5fc9A78rqD75Pb4lSaSgrPftjAwgk7FfAaIfQnzVzCiQnIE5GYu
IB4GRWUD7LIa/TO+/GW8YKI+je3fm/jUlwuPBKfSsTzkUEdnyOicvvwinyyJlQgH
Q2BOAlWyr9LuDtUDhnjG2FJFV1jbmeeIBIowrmRtgWcYYaH2aEq0u43Pxf3k1gFa
XMFH87ez+azPjk1vGOEN8EbvLrw5eVfZ+6yf74ygjm/giIval04RX7a/Didq/P38
s1DJgDJgiJ+582FNMOHiXueX170xt6/VEbpgCRJuzNCAbb92INwgvIl5bG679xwd
DzKIaT42bT8prm/ljwMMos7qt2P1GnWc7D/vHLhzLDvK6GuO9zdY1XymvWLfONpb
SmUllPkaggtTeTACYIAJpml322f1VwHnnC5I7wo3mLGhurwWvBCYECBjSFx5jpxg
Vak8KQV4zF4QZJNVPEsBdmwMd9+XtIkJVyvyBUHZ5vXbZEtdpoZjfPSsRnldB1AX
78iHoEErBZ3EPuVY6NPXxc5/9XKnUIC/51DW3iTJ1Vk/J57MJ/rW+vK2YGJ61yqt
W9hnq+v163xs9J0k2/NtiBI5MLTdbvoHMzDU4lj1ZoFuPd2daLdh98fn/hFPsZ6V
K6TSogpjtN1zh9RPu6ATzgBsYzoP8LzdaKQSHhbVLMOu0HZfqJ5s1l/bweoazMU1
0WQ086Qrv7MbngvZ+opcqLno7QAgkuJX9SzQtzOzHlO7Qg2iTt0bszdd8aUubXGJ
lUru3u1ZVCs/DdkkQxg0nPRECOyO4FQY+Q3DxXa392m1sIbFcxA2guSYcKeIU+BW
nj/2SzQyZlIIryqTbbqRFS+3AWJc7aNUxt+s4yumeNU1Ded+KRWGCfuv+1QPYZVy
eYX7uwZuyIRh/k7BrVvygCr+4umh1wejfz8yPT98c3ggCRqv7cMQdkVEgF24ps3r
BN5uAAhYqGlCPemhaeD1LvzykmuRKXcPf2xv8uL5abPHfkIWHUFlsQBjcUBV1mW8
YUVz+naqsXg26g9xLD5LmGq1bPOhdqDn5Sx1l4Gj3tiZuvEH17eQC6IwCZff0p9q
IDi2ML90E6gqENowax5M4yo0jI/ldNQS0Y7LzXojnBDifEj+18iQm2wf7KIjMhPx
56A44wHFLSGc5QyT0a5l2PxZ1Ee6w+W5/U5pS++3TiTP0Jp4LZJZ2sMRvU7elQUs
ksGuT7Xsz9obfrSKk7tEsfV+qra2VH4IzYBbPAwhaYDlwbMiQ3/o5YMdrcErjget
8+QmDN+9uzw7KiagaCY2WF6g6ylVpPkIYLzwZo1sDOyfeeBXpX7AK1m/KfouvwI+
Dsrre0BCH0DuFQix18AxWKTBM5ALGgtMH2lzrtwlZXsYF3z2sbW8BxA+0nCz0JSG
ZllgJc08WJZ+mr11dJimPxkWysqcAwMZsjv003gPChVfZyPQ8ci/tmqQ05m6Qzr3
Y3RHl44jHfwTD0MnHmAp35EZvQUR25jxEMoJXJArpjezm8RPfQ6p/szOPQO3ep4R
Tz9a+Dm2lkS+KFajJ0eZOckfYZnvXF+lE0XRfn4JvCZAH14by04Ny+7hEE1iYdPB
zuae4ifqDEYpH6SehjZjWxUInYLsWSRdYHiVT4nYcOCj9Dc15Xf7GlkaLtpuL59M
SA9FDUFrOndlv0aSYZ4cjeWrNeqMHq+UdgCpmwfu1h9dZOXx133Nq3lN/yIuPWTp
xKwlDO87lOvlftMXWNHc3l5XmlRxRRBG0QmWuqCUI2mCoAOOKwQmKkPP6+p04dva
LkkjMOQ58Mfgil3XmJdwcKhSY0gEy9BgSAnO1Ch9LAG/KATBTBBjjeBOln7iLNl8
e5zKfuoQdu0D0hr875W58mg79eSu0ChJlcrBkZjEUDChSdgG5HmmQqB/pROEy0nF
xwyXsCIPKuoFLiwvua1u8LGkR6BQeNJmqDBDAIJ/ieDoKpJvST7Gl0oNE6oJW5Id
/6EcJTKyy0e8wiG7zAcr4souofd9DqCMsdOEamBsBI1cxC1xlUa8xstFFjKXOToS
NwaHtk6nlGkvJzGzaYatXkSC2XHqufL4aRPK+HZLctZITbsKsw1JSketKXSmdDX0
N6fQ6tMfQqUIGa1ksI99rrWotDgShv40jDZ5eIdLafXT9twu5wzor/dgis01KTd3
VOet38HJzwqvbrWsrHFCPS2uLak8GCWgwhn0ddMERkE2pKQ7M77DvANqq4/UIfmD
BRZMi/n9lQzrgID4OPdoDhgyeVBN/nl2oVhE6cI3FRV3qW2NOZ19vNYwED8TWmpc
QitWa49KVvgnclQWFldFbmxHklZj6Ctqcz1whv4Zq0zjTnwAqt1c8j1BDf/nupKu
zsG0octRB82f8lGVNsc9+LuOxM7G0BDvfUs5VbAWjKp21hzX2KHh/+RGVj93yJFN
hiFvla0uZG4tgHzR3AgTEvKxrCYemtg10RZ0EcnVdra/gPxGiS6DUyq1pV5uS4Ix
Ns9d2LhZIki5SvkDJziu4zF60L94UF/yEaKN+95ZIEZMBuhDOQDHdURanpVzAxhW
3gpO5Y6IDdLvQpGk+LMmCMWbK9VXZGJfv3WPq6FRYJCsTfb1oPaqZmwLRdfVSd9O
O3cPKrfBHwytIQJELrFsus7cMFk5dKpytoZrTdXrSPbVgUUJ+ZhtFCx3p7Tw7YEp
hgNemzfbVzYccH2rKD56DHgMyHJJLQ+iapscuZq++FahwtrAuvfMy5cdJh3MVoFn
/ggcKQkuSToSlR/EBELJ0x2fhlEdxw/+fBIYICY5c6M6ZQNaTFOZF/ed95oGnFJT
aahDEFvXVQpHwiKm7jJW/C8FozJirMjZhpssOyaOAizlZkT5tHAQdLH3NRArf0/w
ZbUmmG340phuKb/1/oR372jMEenDfA9vWCZ03aluQaUhf/uEsxoyGXUMZ+6ZQGxU
ZDnTcrluNTudyYd8mSJcUSquYTFbYOgJb77wE/oxse+zCrRoL9IkhAvhUL1nAFXw
Q1Tj/tv9aX/4qNf9HyFxdxg65Em3RiCYmYAscB11woV+ZtQDF+X/3Rg4Z5vjf1jP
PvbQI2SX2+4+6mi2XZEURy/pyFLFabQ3YF1AC3+Zfjd4srm5BoYgzdvjvQFPEBEH
zjZ/Zduuk/cttYndp1IIsb7VJpS0gm8aTAbgqrxZ2G69UNVXkNqQ2Jp8mksmLCcu
qc8/YMv9LHBXcd79tGRc3JadFDpHbCeMAoH0rdUPY/BwQKoq3dHK7TvVZ74QfJwe
kRTYOwzb7L2Q1DEykQ4zVTGjQTSS63+R69ZGPNyiT8BfcJpgedYlXJgMTg8o3F9D
sIXhwIbhUNksOmawg5NGP68gq2SYkfnd8o5jKfLYqgf8qfZqSc3tkjSDWPW4jOLC
ee6i4H31qXXKAaHIffqcAvGy365muUlEsDlsznaPmt4MjQUcJLR+Y99FzSKlr3UP
3a/PqvqdJs96c0yOR6V8oM+vvDDZkXk0NVHKG7ACh3ncZYSEmMXI82xg2Ztr5ZWE
Jw/C0lxl/R6KZo5OI4dsstP+0OsFINxbPdowhF1/rRj39bcYpqT3OrtLTBiTDfUp
4d03ZPouxao1nFmZj/VpM1kJn7Qv00vm8ZzK5/9dh/ZwhU3xke1cj4Q9Z7Ub4JEz
sQYo++lXkbNFsIGemurbZx3txNB+Yjj3L3DSyIhSs60IkYx14FumqQZEiNjPQS3Q
glDH8Lz7hPLuHiwGbzkDjzLqheZbfIzwCNTSydJI9Ssf0BfOTj/CBSEks3Jb94Cp
pdqBaiPH3OxkLkW1iRMoNBDBxLNbP1jfQedoq6/ZiRA1mwIGT9PM5pW/xxedpNQ9
B/4dHTJW4BK6gm6gXQhsPtcLWMn9BLIkuDNqhMK5ULrA9FCnzwApjxxLAfuJRm+1
99TL0yXEFKkloKNzN5EKVqKrZGXI0J+TR1MWlQDMR79Vt8T8KxUQrYik8GImB4Tf
nQG/pYRlLYeNhVVpcn98Q1C5bmrAEYm1jMB8TH+ryR4y4YqcNvP7u1ndyiiV6Gah
+F9fNGrT78Zc2pOrNhhvkKJco+lQFunSJQ6V2Na7yaGzwtyo7tACt+wzxSOHvCTB
nSZPRLlvnTxSpvQKTz2zS3EGB5Q3jLUW/83w0ppcZD4vqSYX35k6vaSN+FZBI0j8
dOQliH+ddLxyLNNXhK6KOpnFEXRce5qfz5rciGlfiYjSnuuT2HvIH07kGeDz9+Bk
YyVtrftutE0MTYHxdA3qUilpQKQZW7195e2aFIMRe76expBB4KpCFwx06BhSu5WD
u+1TRrAyQWbcfJQTeoMfSjr8ESfUTfWVRboX5j1Kosc5ODW6MMwzAoReQesJ87LD
/NGrTZBtHY7EGPAUolgEmxhDWxWbMRHU9gKU8rP8ab5H1NaeoxR/ASOFZPM0bQkM
RWtzssMLRxxlWkm2Iar4q6MsIDf3t1p3DbwdCayxL9b/IfS2E2jnMyvzc18U8BvY
cOw8uuP9yKv57a5Z8QsB+a6Iwvz4SMN+mKTmUsYFCn3oYVejvEOjqNNxC5M74rZM
UFm/n5aC6x+9LLIxFmj1tcf9O6kFH6+Fv3stc+SD+dXW6HRhzr8H4M3Smk8rhEig
MilhtL5gSr7BEu+dd1Xh0rqp9dwvTWUwv4oSF1QJoEeBl/6GFWzSLFBXtn/gnblJ
RNT/yhHesWbSfpcRoZCS6mMwX+yQgQPnW+qV3DTSJejwoEbg8b6XVAdRwfcUzrEn
NtLoFKDZAVQAm/6nY0jrSHxDJRZRFa9HFl+2TkSbSITxXJWqrze24EVBLgxDg87s
IPttDF9grDSutiZDJ1MYEkqzfw7oVThW5NmkJzwcqY2616l84kf5R5dLxhjCIImo
QB0PEfUSJUwvNmfIOonUYxZpA0+qywxYH/PqY5T+YsBuecgDebdjsLsiHuWdgK5o
vt/IE7NUrJc69YEJoC21pYS/KJeqSdC2kx73eSrAPn7kkKJsoTIz3iqNBJ6XKFIS
DKc32tjGuUVeKev3nbrWRX1q4212sjedoKPB/e0kn8PnjvgUhmb5cz5ZlpSt8xWt
Pt7SKQUtZMB6RibpylyvQwJD9lkcjVWk+9Iki4zJV8t6WGkcPb9fo0+mZjCHr/C0
lciGKrQI8Hkj6uCORSQvuXW2fic/zmrwMAzPmGqonSL4NLcMMlFwSyFLRQW+8H2M
WU0Rx8qmsgsIN5EjY6qhsmwd8Pqil2FQ3SKfZP7N9pFzFI3YbRNYnIF9tDDgLm4N
XVnW6noNo3zJKIHvExtgt71B7xrTCNGLPYvKHvdvZauyWccP01RqzQbwmMYRp0Xl
xgXWJxOqRFe/KIfDOFONABt8l6g4RYVy17vqg+di90H0hRaIY9AxKgIs5rXucYTJ
X9Mr4DMu6iMLsO8/5of+cLWojUZXt9RuNmrVHofuImImlqwzWT+PVqrsIiDNIg7p
TidjGYaHC0i59XEvOLotEqb53aFVueaYQGTBTVl3vbL64rRuKCnrmOFXhc8ZqFzi
shc96vml0R9ANSYbN3+bzwKLK/4ryBCqrSfhBX+In/QoFTokioGIyDuuZinC8his
hb1HM4FCEHLkWgSoByIN5fgKuQrVQndP7GN1V2BrjfbsOTv/k1XDUmWo3X7ssU/X
qf4KMR1ha3bU2hPZgnsbVl+YwUfvqhxIsSP6CVM7KjiGVubW3SVk6SNA70iKIbXe
E2pf3eJs8wYi22ehP9v5/Vz9M7jppXAjDznFBpAuQwlz2JDy5cY3Qa1V7aMTGvsv
t/CfkvNwMIE2px2mDaD1MKhDH3/Bkhp4g3YlLF5SfqmOu9d7FnkDy9UnhJDMBEEy
amzF8q90qJ6fqZnuD3AWjN+oDChLxy7QyWD0/gnxkCW+SuwivwRCbCFdN4LtC1mm
ToSPovMAIozWY1FftSBg2NDnhFxG42jl8FTYcuf+aEN0O4+IVNjKrX05KnBq8/0J
EHXMe24ArnhzlTBRpK93kXICSf9eWYBtZjbsDM9KZRV868jHa8WxNg27f+esX4lk
B9XtoJStxyhsaikFeh22Y7RzCaVrFjB9vip0zB2e+CPZRpTs744nGU/ajB1afiXJ
PMCk65mFUBHzrquqTfcyouE6DsaCgGSU7gdML1o9WTcqA4X+GGG01dWEEr+4xpRN
Po5YV7TxFjRs645JOPFVx67SqrbmbraA0ec5WPwrQDG3YgNDbeW/Aeq8VY4h2U4e
Tp+JGCw1VgujxBOxF8IqAzVUEnnBVG9zoG/86J4FCoNI1u4vfbG/1Mp048A/Am6e
E+c7bqihMXuzi+kMn9qpiawwUYLJGeZjmuk1aX57PtaG7/FpuWt/glOcpMLCo8Mm
uYj37kCXouOoIVssOfD/nYeEsXTV5PdwGObYyazm9yVz2QQCCmpGR5sHpuHnuKLi
xdB1gvZW6PE3VDNo04K8QwrycJOwqaGVxB9652wE9WkAM8loJi7auwAtZgWOqEKD
DmZFyYPDSnkcznjLloUhfkwRNrqvucWpHI4pMwUKaY/SViHmBcssbJ6RbDx1HDKo
kRnJFHicvhLfIT5sn9qfHD7IErdBG/c93+gwlynXV0EnMWak9INoHzUVI239jJaj
OCAIKSRvjVrjavVgvbeH6bIoVGyjRrU5QVhwdoeh2w/v8Bm96rSmhCF3fonKrIjo
SMfU2I7ATerxyZLew38F/9QTuzOQw+0J7Df8OxrBOcQVc6iFdrmsPqFmsfyrG5LV
qvzX4mSvG3Y8bVlZe06U7AjfafePHVK/osIAj+C2Zlm+uwnb1QtY82LK/y0qxe0L
DJMa+ncNvaY6Ly9ectpLyyOrBVg+EpBASh5NyG8JXPB5CCHU+MBtKyfaSBIxJF+i
0JVbXyX/FzsCPnWaZOEJgCQHrf670IPaEycM5tNp5gJCyrhKmlGkFms6YjXroMQb
h82LiXrhAj3KM69SgyJ8lypDyylJNSUTVx+BgYhla16KazbdApbKGl0RJsSIrXoJ
1jFglEINYZ3eT+vWJakHfkAjz85CM+RQdpOPlTm3Px0czq2c7me3htJdTPlD+XQc
jxTEWg7yIW6v/cEAmXDO8fWyXCNRNMvEuVkYb/YdKkuiLai/1siefgoO+orJrmDY
suebNXrgBtDZFYyZI7pOyy2E35zx5NuNJ+0WPFqZHjQGFbDA6mZLVu9ybTobEQPZ
FNKyrRpFYWv7dTEpGizOUc7LuPyVGpgll//Gwj4CntuGtAW36irn5Ov6nz7gfjjH
9ecupjIETyGip83tSEz4AlWA8gHgn0GeyU+h17zCwuUAXept76ge/BbJ3HqPAk8+
jjZ+MY2a9E5HXkm26jVLHK1qx4KMDScFh1KtsSSqB7k1Qj9Qj7MQdj3Ih/osNSUp
1svEVeloPI5tMAvZbeWJXPHuzFBbSRFFby8Y450QyWTp9JhgPS3dWOZEbCrPG+06
vhUKk2kuQsDD5/v/sXzHEN0YOK6TPQQAJM346AT8Ra6LNJ+2ywGRXeaH4iO0p6jK
kXGpnYmY9+q7a6eco2w/SHnq4wNg/a4EpPGdm4AmvBR6T75A7KEpX7vn2LNe6DYY
Y5IR/O2om4f+xVrFO9fIH7J3mHJon8sFMuBtwumXmjhwHtxzrq/cniDnR5kBgk1k
0SRRc1dA++VdKpWC/YMTkJG6+ronDW89cvRjnyLeu5kh4Ul0uGv2fHvP6O6GUdbo
pSPrrhIl6Q2AT4QDg0wr8RLZqk1RUczd9+RrTErbPY+ahJbVYLqfky4r5zi0PAJT
+DJZSKD+JanKIXmFzGgxwDwAhga6fW+uL4Iy3cvkQOoNolYZTz0AYmMBHwxvC5Xj
Zji77BEtfpoFN9/rNhpbbBiUjukN1HNNJ1UDOXC2bgFUh7Ms8T1N64FlpTtaYRqe
/J5tsYZNQbP3ULK5KVHr9AqDKdKqpNWmxGvUpNYMY8SBInM770uS/+Qa3K4o15X2
XvFEPBsCCFDsHfvMe9za/S7wSBoqjC7VyE2nynaBk0HFJw5IC8D61imCGouIiW0b
Yzg6mA+DTHItLZMT9f+o1i8l7KDk8Yig/m0TPzgGrIhAF9V7JRNM/7GScn6+Zxtu
VXobD7COYRERlP9Gq14I/ysaVTGUbvilZZsZWAafDYEW8VI3rgmF44/b5DUPfYF/
M9DLRBZ3CecaOOkF3jtT8SbN/mtTggE+JpD18UVD1LKIcqfMz2rU5yZg0+Ypc/hI
9uQ8DkblYxZaJ6/bgba9f/oC+Np7R+FcRLjsPM1j8ogcbu0F9MI5mU5pYLmJwbAG
14eYVr2Pt8pd+vF/JeDOka0HqsRDVEwSJBpQ5OpP1wM3w/bFCrr1Uq0o5cqNkc+l
sZyh/CayfT1sAE17dSmzzd4XITAf0aufB6YBxBqEAUevBGF0Z7k++Q+EJM6TZDRm
wwMlef6WXP0FMaBFUxD0jGemq1ff8CNEnNN0UJFgR0j7ExF1eOzqVybF1jbRd6I5
pLMJ2zHe2g3tNw/O3aWEaOeY8kn5HasFxEvVKdixGxIJMZ2GXd/F3dvcFziJG/oO
ivAkAPpAQLc6BD1aiAAaxzWBAc9S/hcTRrcTSGf/0hNbs+ZXPX9VBjLTyiHSjir7
JrfoGbdYonQgFi9IxepeZyEuP3EVJhPaF5HZaCh0M79Ieb3NB/L5qbcXTFL1jAO/
Y+d9PhhmcnLQeaPnZ0WjiqfdYOc9FjQ0QM2vdB2WwfCgnhWhMRSMBJRENxvdqug6
19WNXcjjy4+liECwHKd+gDSSKokDncf9r8Xddi8dFp5dujWnkHLjbWymNipfjey5
1QwsY9O4L9YHdYLxP4icO2zOGcQ1c14qx6SVElMU5o/sFD8vM2E57LcNvOl2NZp8
ePS0DMTIV8+cty+I62LVse6+WwRBFse9mleXmrIbsux7z8JW8SHtsc564dags1hf
Ox8BL4I557GQ55j3J5sz8aon+zSwCFIghGrzJxyLTFRKmjaITeRleiSS7FIXdius
fjgVFStmaJfYdELByezKHXDP7PN1rmp78adSwLRueEAv9vuB23OOgTyhpBRceqbk
7brqi/kh7Fwmegy0XaZMYx0dxTNAwfXizUTkdibJStNnjfBtQO/cW0DdIc/1j3ro
ONptItI3PbmHW1KVm+wHC1fAI6EFiN/v80VwhygK9+d3Hc64vI9iJexGEs4hMW+r
Tc56KdjINqivOqNFp76Xa7Wl3AZ3qy2YK7jTaIjr3MnaX4E4IUbfdmhZFL5Evd2Z
vFKcwlbbkvSSwIFj1S6qk6O1T5jXEE1X5EifeBVxgzAbJbpLhtkVpx28WHaSNrA3
x5wFU68kozK3SUt1uuEWoc/E1hhK3gtGtkuMDtZIiR4UMT4UxzFri58XtOpMOew1
2zlOGOQNFGZ+4gYao3CI+rnOc6hxrSgYJ5O4faTjY4iHjv5tnXLvVGbbAZmroVlk
UlZTApFAIORvWNBAe28ODGv4Sy0l/WNZshp8GgN35/t9WoVmuwufKvU4dIpxwA4A
Zb+TU2ve3YR6SvRcF74o5+f1Pe3NST718Xu9aiS9oHQlpl/CEcg+IuxPbNpvVdwM
njDCAVnqpQ8ALgXLc83rCn4boVvib8MHIPpwF89XhnwWATC7y6y9LEz8mhHD/0Cc
y6OzqEeI2kkJVRkwyOoHQ7AFgbNK6Q4vwJcg5iyBBLbetUwugz8G29MAdEJ/D4j+
Pm6SMISygkFq6EaLELXwrKiQz/PqUNMLud4kzNHp8aT5Eeh6GnCvQBpwXpSWju6F
9LoK7TtsWlcu0U8YFvEslWKhsSDrLwO062leyphc7huxBEOefq53YHchjPKf8P9a
MntsxGm6ObGbW+veIAg94/IADRZTX8kj0QHTVeKeAakWnEZFLhah9cWetqLv+KdH
yrTUdoXLjwp1/j/Y8lCQTohCRgjndbtEEap0aierWy6A94PbJLECh4NYKBe8xakN
eyZvU9QqJKLk+sKJbBst6AM9Z+MY4YxYrHq343+k4V69N3ItqhSA4ookiGp1tkJJ
KOcDyNiLIRPHkYsMlLbVSxtKNxHCMdN1Yk22wE0MuDFW+7iGgRjsQOLhBfk96EmF
iB0hdNb/dRVwrywjDiHHtXxZN3OwHEHQYi0QodZiPTRopistgsTKXlBuO1/8vPH1
ZTkKV60qPpbh89/3+6j0rJLD3jGtppKqqHgI6dhxO/TrsBxXbQ/5haKbcRq5CEh4
YEvlNvy+ynYuySoYUuWD+7jUR/f79h4+EijjrgQxH1BSQG3xRKxZ6G1pzdFO9zfX
2MeZ+X4GXYvKBGJkaAjeT1ZdZs/Wo/gcm8hXamNdU4DxyZ1K+iY23F+xUAFaevq3
t4cbNVZzACaYNfiZtDSBWzbFKFAeLhnPwFJfpHx3wm2FTVmLgJFC5Fk9QomGRlbz
0thjtH/5QwAKoXjwCdAJZ761uDYgokomnylaabjULIDi6iHJv/UUx7MoeILQ6pQ0
GChGqStF0FvVg2D3S82Jl7YWzKDt3aCsgCOhSKtHHHHZ02HNz6Es7uS1iIRYzgDA
wGBhPCaYd7RcAbu8UXPhpKpzlljpF4fbck8eh3Ms0OnOCS6pNAuL9hE7QITZcpaM
N0pFXN/kXKBWK9a3IOKKMvWhvIyCtCeLmloAqXvssqGdYgCRx20tl5NhhqJd6vNG
KjKW1cFMNMsS+ANxbfgVszz40LukAiKQymnGYU6dakoi6Rqt6SH3DI9QhwToc93j
zna0qVRMTiJWABAD0SDPJOlgebvJS7muttRHScF4q93fHc9SlnFFAmZBqd3jl43E
2HUKGv3UJhZa+4HonAUiNS6H360JqVHsvDm7tMwG/7p2UaY7in9AOUxlYUUnoDN7
0HxFWfnmE0WoGjeNUbTYhWgp4/ZN4leH8x7POz8x1jfqZyfbLd+kwdiphdunwp3z
tP698x57esX6LKUZnMlWpmD74tT05WIlpxLPrSJTRGbNU0Rb/OGB+u+lVTGHWkCB
u/jwAvqvzI8TiRKubjsUH1mYn/5fT1w+3qpfV2tPT+OWC7uowRKt0FF/+7c3jO45
P3nhb4zOkoCuiUq1E+otZHOy0hl8g6mjiEEHeLvwl8t8hH28ssrKWtL21WvETJj9
3Y5t9uTHv7xfl5Uze7PpPxF1TfRDEvzlKJGvAR4BEoq40anbe3nwpfBLaZYtb9fr
lblc2gg2QNVxEUR6bFEFg84i1f21IcCUO2k2oyI7Cc1qT+vCdfKYyS4xdcn34GhJ
rQ/ZsWzKHzJQmDHBq48F4opMp2YSeakRMb5iNRGIhpOeNzZHH16Q2A5pe6L8mE0F
lKSZ+9GYRN43UhjXX+MhVZNzRkMUG3FQgXc8ZC3E7b7QT4Zj4SW/x5kmS1KoMQh1
+2on1ZfGQ7Fsf3KDH9Pask+m75P/NXkIEu2Rtw3Hu1vVGpID+zrp0iF7kntkNxXa
tr5uPi8L9eCwqdaoXt9QFgvWj1sHWf0DXGh42HQRXHT8CIc3LW7SbiwnvcnIJ2To
voheJRjKQi46jhe5LwF/3jQ+lhPQcO0LPlRAeWfnNICiKVEFayFS47juQ1xskXG3
nI+Lcksel7H+knq2CtXFRZBzOQY0Z018G99o2U58wA1hj9/QxhMHKt/uLiio4/Y/
4VpSkaeRDcmdqd+iO/1xw7s4HESf/NFixEJ/3wYorBA8tEXrepM0lirz5MuvqwTe
h6KYbpH6cn2TYkkuHZx6Xj69tsXq367hbs85ATDlM4+XfMbjEAkzgkfJiDMndtNj
mm6fAMxIndMfObTRXncqlT/P+geNtQLqAQMRoMCPV7pOyLbkXk2+U26KfaicH4qT
ZsWsaufHpAxEJZTXYZS0i36OjeylE1QYv5BvtIr+hT/tPtbZtn/DsjU4JRrnaOdk
97U17bMZAGt37Lk2f6+LAffWQaZ70d6ybuJrUWjiVbqAxlfvYf7eXMNc9aZQSh/z
hmGZBkY/fFCeoHeE9ZU8rbas31Iw9558ORV9fzorPA9rPjnJkl72Azfo24Ixe1QY
g09baXurikTBVrSC8kC0wN4ZGvI0Atuy/q8+3yqY/9uG+0rNHrs3acTw61/ojMmv
WokA1qHCeT2wjyonopMijITf1eZJjALtIFnb5AHNLFp1lvBLBqKAQehyDFXtTL3P
OZXT94PA0m7YWNY/aRavPOhzFiketafWEnI4JVrGvlt15Dc8k34SgGkkDbFICYBb
glBbkGlv2sm5KEI0IuSzN4/1F06MSrYhCN+fUT/bTtMgt0RWqUjccHKfer00canv
aecAFpj5xZnB32UWK436hT0JCBaeNWWxmJaV36OKLKGVZ+HTfDsUpHTC2HeQYt1r
dUi3625VgewwIPBOVDMPbLiMIdQ8kpWhKy6JrML7JjY7JwfUAonvMhEe1dL7T0gH
U5qKEDPuz08+pFZ+EWX3esh80KoQ03GFJ610rnK6t4U+Ik/SebxEW15L3jnFlnOb
eOmxEfdTcGhbu4cS5Gn/6UOS3VAJnXpZGpZB4HXW1qA6umU6KvqWf5YH0XJfSRQG
n4E32SPYclt5XnljddvNvFJ/i4TG14ObXBNORh5YoLfOCOn6BszsG1LFdbtsALqc
akHAz3wUdluhwnxWcJz3SvHGPkCT0NvmCTkcm1P95N2VjPDtWq5Z67jEcFdx5ezw
tao1CN+7glxnoMyd/5YDJ6b31ypnI6DK7CIVHjs3y6+aj3htWc+bqDtCqfXkESwH
vA/nf5E1HL3q6zmaDEYvLdf/73ML3uz2stlv5pSsKzm7QvJxL/QUcxDV15SNk9vG
0ZCPHdjayhBoGUE0Gr+05PIZJ2VqbiyHd+xVT+8m/S+dCaae5Q5z8UZDL5csWnyc
+gOzZH8HqJyYiIs3mMT+sFgyND3Gco+9GUx4OfLg+hlzSCoa4UD/WyzHaiIrQISk
ImppXyaV3Caf1NprMa1fLMx5Emb/+mxlTmNxEVv24hJy1o7DBGBZjs1MCeHb1hmh
7SyikjnoRuQ4tKHU3khm/dwMlSCQBliuB14IYBQ1Hqv6zPZXllVYvVEXBYEZpB3y
YOswCXZRFC/iRpQVetv7fATx/zHX/SJbUEmDrCpNF/tTJpji4Q+338wzAGEAxos4
oCaou/q03d+WO7m+D3eJdQF271ZuwBL6BJJWYanuXcodlqPKvF1Cs0LUARXVLgRF
sEL/TncFe9sA2Gu8PFtv61NgL0dQHtm6wC/C1K6sQplHix+Th6uGpjWQre0Xw3we
mz5y8QHE/nvX/xpWgyo+LqQ1xzlReWfqqOwPqsnii0SVUoSkX0RNIGSAp/tMGAQL
y1oChGa/x+GUasSRJNimAyI0FOh/G8iO72HkAUqhTogQlybEYlMEOSl/pMo+TWV1
HXAU4o8Bdk9sZY3Cc/c4gujLFuLUMYuqBQZWRnaW8p6aH8HOQOfdHECwKlPR2g09
zAhek+gzsz+F9LRv82D+GhPsOM4rpKLCdcV/JoVm/w36VU7Llm+dPlnEq0lqpCRs
KTlHDYoOjdiU3QSLrlaTpbjUyO3oc5wml6aUap5L2BhyOCiv4drH+mutfxAIR++a
LNFgBgM5uqqGBMuDbNnBmib3BH/p0/dKI1nzpFS8KjY65+xPFhJd3Fnu/JZRaF9h
bxfA0A7xE5OxVmiyom9zVT7MNQMG4fXp/lThfFE7oAdEYh9TeNXKMM4C/ZW32ofA
Wo6oVJz6WUOVaAP7woOMflJ7PhE/qeysQJLgmOTPJ/jn42OwNzKvO6CZTmnpOlHT
AKdDbostQAqJN9IqgtDH+UbWtZ1qVeQCpk+Q3fN9bZs8BHeKqekjt2jeszOpupuy
FWyxqivCwWA6rokH26I+vLHyrP7xfa7seKRHrc6IDuU6i7h64dLskhVppACeYXgo
gRYvC7qHalZorPk8fXevCI3zE+wgn92l6jxQtDW/t4s3eQp1RNhbNW/PGhxCpQcE
EVY9+2Xp9LzkMorizR3DqmoLKhfyQXOwce6Jzan7Ntj2XC6EqePYEDLzSeQ2Pq0M
WbNxlfXuwu0Hpq6uTctS3Qa/0rTyydmqqqFy7TVAm6Xlqf5SwY7KxTtXHUhKC/Oe
SKpGiNqaH+cepnwCO+F7aHW2z7zPgFIEvkuAY07lI397gHMXHXM0kYrqg6RgOQ7w
v77tU6OBIsexwbBmKMT88lSS+Ao9zLIGe+MAJ2rhOMNxY59KFdcwFqFBmSExiXpZ
ZPVig+w7kVjsMGTF1raEVDELmyguqAAV3zqt7EB0ZqFoJhUCpUvaTOp2jvgxqwai
QTW3Ov5mMapW6FcPF2xzYoK5tiqzqBmZseLBLT3A+jbbNj4B6fSfNrsRdO/LYuog
eor+6YcRO2VHhFo0zWfEcwwj76Sps/PDfwN/uNpbVsuB5nO1vD+P51Q5skdY0piD
Hf7NXmXcGTc/9D7WlyRGrYObjsXMPghsIdhdZWvDZxTg9kB/syUdeX7FeCT1lV10
xus5PCROyk7DCjlqxgrC6xFCkBYCmoTq0Yqxqqn0FEDhVHldNNMSQJORWteg1EGb
OeMPVTklFFY8TDy7rchAEXFC6p8+z70afS4bGLoqKtR1YovzXdEp9W77US9he/ES
L1I962hWgPdOwajBZd5slFtxIw/IEYNk7UiWa+nGMFhmQbYm/ViR54JECQ0IYyua
/TrxQzN13o2vC1uA66ji79EmuvPiApe/IpzukSmT4lXvIlyDCE8HabHRXnEancCx
YEmmFhQ9lE+X1W+MyfzXYiP1334WUY4/sKwL6IX5JA3s4C6GfWHyMaVXgaWiWsF7
W5fYbtAnMNXL24vhCKG2IimV/hAx/B2CCwpezCVFFARKXyeWN0i5atsxDviQyTkQ
6A83rFvVoecwPk0B/Fl0ZdofVjZx1+y3pi91FjWkgDZln1+QX0XtBkLysdnPB+rm
sdp/BwKTEykZYyubW65hbE/h4EfdrAmBoZvF57XyQIrVZYOxzbGZuuerxsLkkHXD
uuAs+O5Izj+xbxEfPIQ+1IMGn/TpODjQznG4GOnd5+547EvRWBvB/cY57upFlPEn
5coHZt2xsfmEXoZCGzLEHSIQZ++Yuzl1BSIqgRuN5j+k9TzMB7oppsCvltQAJaxq
6wtP6uqiQ3zsNhag3+IlCoJ7C7IMsgXxKe6qhAmVp2016g4uhJuCjcliM9dzAjX3
D6NRSWCdeXpCDOlSOU8wb6euKbQfokhp4vy9Iz6jecB9m/KyMAksAdXa/nxIBGlN
fGVaqSj/maG4R6ajnVfa6P2bpsj5Es4DO5rIm6gOYAuc3tK2FPacPNj26/yu+3NU
HBDdDZnfeXSWgpA9LYThfPB3iCvch2IpZ/sy4RmxBxWT51bVI/uSfvpZ+m+Vc2ki
JwvY6jM3fp6pT62Ed6H4bgLkhcH/Ff0CUZOPtR038u543GLI09qIbS4TIAT2lzI1
e4rLcpnV7uN8uzx1YW8+Zx11ZEodtsuT9Lf01QKpx8rHl5aRluhd0qNur20iGQuY
VK5yLbbCG1p/JNMk67O4cQYZugJG9EzYDqUQoEyD7kzDHqSmCCrgGlaHqlMyHRAP
QNn3T6+zgxVb2qODQn+8hnZaBQiQ8zvLsL5QzMSEHNjuu+l3tObhPKZe4nXYZI9V
A6/ijFEcjk47XSsC7cDTcK5hMfIcLMkif/mHxNK73p1Rwt5nYd/ZDTIMWt4n/96O
A/XUkMRdKcvlk2BNiYPbz+KiueAaWpLNjko2Blow7ja2pDEccpwD+QKgbvSocDZ3
xt4lStrtZ9jvDJ1JcnkxFY19d7NMh5G/BDmpZyX446uQGoVMezZzJJqoecpxTs3J
+Nh1i5dw2davHwQ/kohdyMCArqHxR2cakkqIqVCu2gxjh49P3XIP/DG49V2WVXXA
Bxb31JSoEHGZtnkNi/6dF0iYiPsXAbFGxXegLdIxlw4t6BdLRZcwz7mnUVsnLBpb
D7IUmoIZnEDqGR6gCsPs7UPDkG0dqSuN6erS66XGkDKd9DrptDOZxNkHcbXJ7h3e
mKOXX2vA18O3WL5RSw6P9uWlVf1DL/a5O/Mgu/w0hhFAtpBpjhE/Dx+11Mp0aa4J
9jEAkyvWha/pLWfi2ua81VHfdE6Q5T7KRJ0wAHPcQ2Yh4roQZtrVbuDidCn3PyCU
0rmQZJ3rxvZGSOWbPd8h0xtK3PZx5LEl5o9m5frgul85MnWhRoM48Q3Ii56ALOv8
nZ1b0mjjkefwAcht7M/AM3dwwazhqynFfLGOtXpzoRJsm3lHokF2kcGe4gsMoVfB
PALrf7jYLKQM3b1St1OBh6YN/RcgAzeq93UuRPMfbzv1NnftYtKM0dJt853aNvYa
Ku4asfqshbPhCfMT6BxlTgY0JF8j+/Cu6h6zcvgqJTMPFrcVPO1WWXWH/Cb1uma3
lG4IkVlLiQFo2iVf/qcW43Sdk5r5o8O9b3MMSJHFwH9xzEJ4fq3ydpjwY8YKVKtB
JvhvVZTmEVypakzpGuJu7ms9O7Y3Kox6JIMbpC3kLe0JKrOzVByay8U+OP0RkaaM
17lXAKb0oGT4Z+DyZwRHxadZqejvOTyu12j1knAryoegGuk8Az9mRFgci37OF1kk
SB75ARUb6HWTrMKq3N0vXov4ToxM6mR7wffUkz0k7adc9CvUQcCxSNMTJUJubYob
di5qZuhOd5+f1XlgiV16tMZg6RMOkqfFHpK8f5bsXJU8eTxhKaN5Fn+unBWEYeg1
JBY5xtN5Vb+6jnp7vJVb5unX1k8hnTfVrhy1qBYxfZJKeoGBWOMD+ITnXKfKS5wD
c/UZz54/m6zLBqrKw+qfva/exsYCJ0ibc+xYiwmWxWBNu7VtKSi7uZKKdQXDjySB
7vT81OVfwQ09OciUuAyOYG/LFHtAAGxObpBErDBcAa7ZGWTVJSlNL2ZxabcX0ySn
ia/bnBfi2+KhPu9hG3QH5TH263iWQejkgVLmh8mp4p+s+KGn/pmpXF20O631/0gN
DUSr4Jcz8EcQyuXIyjs8h8IC9t9+7nJmL4s5VirkcGRDsT7IMxrKCovDW7CUKXVx
K3gMCUJxOico1HS/ljbDxvGeb1R+c7Cjt6my7x46kg3ekNTHy2xOu2FRFCJk+y6W
4yWjz2H+EVtaa2eWglzew/81Z98vrtCB6zz9aG2HBD5C9dQZs6ysHsVsKlDgvb6Z
ESFXnT21gD81+5WDcYlUr3tzXPidLFWSXm6Sro0LM/KgqwV0pl+yJjOwVLbPjbHu
nG3DwtfXffj0MQ7jnVAumlnXm0NpsGzHnhRqTY5G9VqI5EqjBXOTveN5sGI+svUM
0d5ILf+ll39cTjkjfRXdc5SWmAIxU9JglkcSn6iU2bvDxPb0npcODz9XD+QqRn0m
Gw0+RgiprSvaz2zLGAMYID3AwrQ1Bo3xwoMdcJwHOD0MH48zluC0yB6vbPXQjUax
09W0YWlOXeKrILazwMkBsa7aJBRet8J2CFlZ1SN4CTBWub9CY+rBX6I0UetR/ykP
+bb6IZDDLiG/7iNviX7R7sx1IgVMbukqz+Qhp003ekVkTbjOoWC/61tIm1yOlc3Q
Mg6ejnAvcMEdQNSgR5xGsoL/KCvI1nqgbyHC2O4WDEXY7fMdNb0qH3aXIRvAOggZ
9f9YPQD0lYeL7NbYgr4GOVN1o1/jK+g2nkpvksx+oRzr2zr+D6rK79NpzpejLJTy
VWXStgkPA18ks6M/7zFlSVS6+Xemk8pjP70AbYdL4elHEB+EGDA3FvdWOUUf15dh
2BSfG0dWw1dAhJ1gVA1xeXTKta2KnoQo6zRqvHsCd62zjlVBhz1wm/ZlEjQ/fdZ/
HmhXlD/yDQnveISb4B2ZBsHF7ONt1HLDzlU1QUeJ0HWnww0DINPm2fDPq7Lj+dS1
IG0FHQhktHFrytk69JJydffIsIxQ4pYvenPthRZqP/8ImkriG/rWSt+6Y14+Qui2
pMZct7DwoR9DC0efIuPHVet4/BjWspJK6RkbliE9n2ilkxk08Vxp44cq7UuQoS75
xlxRfXHsuGfQJq+zZiaVVlWV9LxG1u8nB9HpVDHwHpMlXuqDY25PLIeYkb+0YCXg
+Vs+prq9oa3yJSGMQMouQThknJdc9ba3oIM5jMtlB71qh6q+eml8/OpIL5+uHqnk
ZAMyH3+b3l7txqWzkhjfLINeOEL+v6rTxNidUz787NnIQ2G9XJjjxfLcMJgzgXr6
hPpuk96CzlsUx6zOI6CZ6Qy6+2aUe9PqMBNlR5TOAdY4HUeJmoqw2+gxKbuDTAiL
4E9oa6KgpydkeRGOmwWRj7C30vvHe/jo0Ndp4eD26mXDwJAwx/m/AdPPXmImExV2
khAqfb/ji+HJiM1Vd0+heDGerNJEuDrkT/CjCLk/cOUmW7LtAdLChw9ofeSVB6Lr
t+rQaehVubmq2Jdavb1SxRtRAXiT5SlQbuMRGkRpJmwSPVQhVRtRW98ELVFQFOAn
TYYMvmQJBHItOtYXM9Qem8xcOb9a4SnqCPGIiSHc8NDYIk5WAdIHWuju0KQB8p4S
pd7jXsHF+KuJR5xCTavUBwX4nvUPDULsyBIP9VM5qQlMkS9UoAsRfG56hwVH+YpK
Qq0oMWLHTk0StK5MxfJ6IwDtT5EHUoRzFtbxxhtRRM0OfxkFQ8DAGoTwT7sW1ctT
D5NM1YDxoZIuWfz9PwQ/B07I9Ygls9gWMc5TB+NaXi9f14ywvzpduF1imZhnBaLs
BkULyrYtt227vfN88nqs2BvPSWl49O/LcSv2dNGVVSNkmjrXnAHort2342iBidWJ
JYHbBjD++ECg+VMFtS779l+F6pm9WS0ki9bjBMU7DxP+Y6DXQD1F0KRu0hHS1yyu
WazyZR44Mswh016rmQCYoldKgDcesHt8qa5s9G9zOwj/fEBiuXQIvmosBUmIZ5bY
ZiYOfpAoIHyBfjliE8wbOMq0LyMONCPpfjOvDfb9pk2rTOC0G4QsRTdKCNMu1bOe
+99DmX4vO5EdaQbU/SHEzha5/gB+geNYFR4313Okt7P/uGVO+ZgLyVjzM4e76/mf
wy/nKLyxNMNzvwJ76+/YlT6skFV9Xh8R24MyxsC7gOtWOQ7pN0HHdF5eWyOkF82/
8/mZWYj20NK4HOHO0CAi28VHPkE7cnrWIPkXStQR2IKSvq5caEO4cLDs29+i65K1
ZHKkawaCq0w6M609aGQEbm7fwUcz77hEbnxntVyZ03yxNdMaYpS7WhtuRiGakBcW
RW8oDo9/SO0GNy1tJlPvqnFKbhgMjWy63KAR2yeJIq4WtP3sDxvqfsca93TcCi1b
oCjmqK/o787d8gvW/joPTh0aTl8gByhkr2a8Z0QUDpavjbTBMC2ypugjnVBlG043
GGU2he7zgEHw4H3a8Zf2USJSSvHry3OHxSh9ItM+pkV9QcS7wVIeKADnLhZ7EtMx
Y7DN3bNoyRoj/Su44Hf0R34zQXMFu9KQGAcJQVNZIeezGu4EA9L6a8t3ieNFGFPr
SvAxESfaBZseOktDmU5Zyv9CXxi4FhG345jdyP31hObhgHfP2VMLjFRkSYT27hz7
nCQbMUTaFWM2k1JKu6wsUJpSeDOGk5VL1O5H/tsQBsf9UOoGRMT8h7rbH/PWxo05
sDPbjMixYaQuodmC7UNnrTubPNTFrZwcPnKNRNHI3U6J5AHvYdwhFt0tGSz/QtQR
bj0U1EXOfnusz/Tv3MFV3MsSTGY3wZsv+HFJPbM/m+fItgZow5gLzxwhsdwi7Mvx
OsHNsAjkbEEiQB0qj7FUvJFSOlZeHinYg2w2qrpD9dGDno7OOUepGRPx1lcRNlgJ
aEdk9HsfFMlJG8FqVZivQE4pv81u/ONTh7CLvg+2xPk4L0CiNlqVTQy7lGFJkDPz
kLqfkNzEjER3G8dvI8AcwzRZqkiIMNnAZwr1uLqdvvnssISScFWL/Wh7wuLN1fEI
YLQcvMFifRyereh9I6EttIio5GTiXaUQhqnbOZUwuywrpFCw75BhheBPvGot+yt4
ByhLckKC4BdDzG5Y0uTz5YCp35NHkoee8oFWDbaEJTg20qw2C6QG/hsYaBtPYDbT
YWnhkAzL5vRyrlZ99CWSVI8VPGhV8PR9Z5UmVoAw7OBTg/w3qVeUZAShySlqkGVy
wcr3uGNVvHUtoH6DWKvMvGpJInjlztQBxjr8w27wbad6O29BH+zbf00V22QzYPwk
n7zoYQ5pgulfUJfUjlFnp+LbYenMMZ5EXzwIFns4dd7LFi+pCT2LfVC5GVE+3aiE
wUGlDmawiLJMoC/IxHr6ERS/l9NBQRGe+MzzBUxJNlqb3C3KnMXAX7G7+fq5qG3Z
Nmv8TtCg2nHQNbdwFshttCySamYkrTtctoisoaiA3QBN6FkhV3rSwzVd0xKAiBec
rHNNJpuwPzzXOuMmUeuAwqYc0N/4zHRoT2UenAK5bQvGXzhQXqFlNjzqM9usRDIx
bD0GMmtdMNvypYj71DVNyTqIjRH2ukVG9yX0fs7IOa64llLsfldHqhs63/cVTPhX
gh+RMjGpyO0Fhox8DGIbkrMSvF+L/EOON9Eah2Myc4R+xDI1yXrSkj0svqH1LE03
auCZKUMnH/xvXVQk4+EfpZuyOweq+Koixegk59VB0ScnFxbrqpTExWg08VqpEAUb
wrY5ACwqo5akhxMCAYvRygztdjXkv5s8ecTz0C6x4awIss1xNXYlqAKAk804pxnV
0dtf417qcnDEHa7RDGcxe84H8oj+hgj8dqugxrFe0gGf/DtrAu0Rbx+Iep5U2Xxp
1GROxuPhycaVNFPVh9CrbkRt+bSN+gUYFoAvdr2iCwY1+m6cJiUFzQfJGYw3G7BZ
QVmJOqgJ0Y+rlxyuwiTtXXiabCVquC3QboWklAls9Ro6DFDecHYDEGNirld2EKDH
9lWKW9O4ZJbd8a1RduS11sUrVoGJB4n+bFWO65JvZ/hbL5hLfURdDkZN9PRn/Nz0
v36WJUyuI3NxwKBcUUkQc9ucsMF22XSO/076OuH5mDt+HpVrpE4k716Yp5HT7LAi
XOEH38jcC/IQ5cVdx89EJfKZZqHCaq0SdhOmgWElG1TQOXiXhP3uN0TM1C0o98Kp
+mYEB6NyodpCsdO77wPFRNnpfE7IIZuh3vdFJk9zddG7tVZ+dJ0Fo5akEafeNDga
b11aFRCr9vZCOe2ixkddOys2iu0bDteuQ4sQbHcix/23NjJIobN6Vxe2ovwT+uZO
o3kEDhchGvhDh1MxD9rezU8+5tJRAn9Y1C5bs8bNs+6FdRX0d1GdPiX5kQ/HZs7Z
DlYrE9c5Cubcpg3GvSwVB/FheJr7P663HnolCyMsENNrL9YZfIa53yHVMqhitCwY
cFEEnUOjpZiA7wzrfMfjlgo92pa4rYjH3nEDaBzug4cA4SnMADjNlY47LU07g0Xo
qzVBHLKWviJePXTQAcnNiweYK5mW0qoSyVnwyj7aTQEuc11EdLIWfceqyU2d2ZXf
ayQLrjG2CFLOggCnflvFWW3jk4ZT9WmLlaW8M9k0BmQtexWebJzhoqckS9EWyx+s
rowITyYUvPmrJy8CIr/t/9xblq2LRY5yuQIqEtTTs6Zve0U8/1DSrm+hpkBUH86H
P3RYGyZuIhwNfaeUsqRfYkb8motEwuCX86vezgxDxXWllZQXgMUkLGISIpIXVb3R
17wvJz3fJbmo76dveK9XKXYbNnPfH9ocYPsFsQdB3CXBsnFb0zrnyetoPWUktaaX
xe1O640cJ1uV73HQR1xUwYcoEKT2xuNQMY6HUCYXI9wAw5DzZc+KMNjTDp9oLPTB
k39qi2hJUXH7yVATxeHhCtOKH4R+2lz8siGk8tvT1tDoB7OVxqd1Tvud9v9+nXek
T5x/2bScdfJXj4wtcKA1nLmi0yaxV5QhCidfbiwue5Mod76a0OjwL3emSR35Ef25
2C5RW6UdR+t05dPXqMNCHW0LviQEhoW91Sy3DbaLxoKVDH3J0wI3L2iA5RyBnpCa
41Lsc4sjTwqlbuj8/MjXutMb3e2d0Ipp3kclgX1igqE1ZL7nz0IiJzenYpweNqND
mE+pr2LsBeTGq7aGsKBEqI1WeSs91BfMGnf2AnBagkcyTQcb+T3PNzlFTz8gEcWM
tw11HtLkoNB1DBp7ehRK0/xdzlX2lmc18bR6cKIZ75TCx09R2Z0N0ieKejNqun8X
/9gSTVTk+24otgtroMA+EZsx1GVPICzfZltd6dcG0T85u6/emZffOhxdQqL/+mK6
3clP3UlrNb8MWQjVAz/DRXWKt+AmmN7asfpIjSygv3gMnGHMmZ8bykGOiNRbf7Ws
swrQVjAATBBinNvmRvvdIYRQS7w2GmYXc44pI4KIqO2V4ZlLx/NWXJvvZnzkWF92
28Ixqu5u80hmLq/W7zF+NpPponX7N+5XDjR0pQE/Eq/9rHUB4lqSoac3HKbZ1l+T
RRX0cKt0g4Xd7Mr1lNGonBa2vLlTDW2K7uTa8HTp3KNj0zgIbuuOPYeW+uJMpYdD
bC4gixr5ihAJctnQ1/u9fmitP4ozarUQWwCWCuz5NHK60AYhQ7P/Rf5v2uqkzDCO
i0g+CPvyrN56ogo/IEHSJYd91JeibzkjHjAKz7oDbFJnCPLVoWfutM87tqWz8PPt
5RSOtCrnb/bUMc0kfTDRYEQiiMzalelR54sREo3UoTyeVVQWnWzl1YYQM8KEKHaF
XPcXZlJS9U4PlyF8QfNEBdigdJMkwN2OUhR/+rob58wGyhLOV0Y+pR0mXs2aM8Pa
Guols/QMvM47dJb1o4ORESVqoIxr1w7vhZYQY411YEyZMOVW5ejo92tlFKDvhDpp
vZehyXZRdVQf7io4D/OHOTlZyzyjBje1MobHZV8QlJsv3RX/BvoiAqFep6LMXfHm
Zvu1tj8RYBv9vqFNwj/zD302zcD7Y6zmb4vgXHqVgEfCW51F306NaGgkEH9BMZM1
u1BnY0eSBwC0il6pDDeq+9xNaA6PRddDlmMq/jpJp1BPbDSEw2OxbMDDOhs3+nQE
iAWtZIRAObqwAGf4VkoMfYL9gb6eqhTVaoGUjSSh5YU9GQr5r7sg9gA7t6LTMLzo
YTQKTjPR/LhOFGkOP6Ts4y15OJUCr+YkVJqfbYiDPIPzo3jCXpHL3rbjIBTq4gNV
JXRgqSbT1pYoDRI1jjkkr/xltI4QjqWtm3/ctq0CMO8PTDmXG+42FLZTCcHZAmJ/
ZgdojkS/B21AtAdV6RzdaM9iRUSTIIldPJbdyvWatHACeSgz626FjDusQGoUMs5S
9MHC3ZO3UFO+91w2U9ESQhop/s7B03seGsscA+4eKWv+toEvZFVP73DnFiAiJN6G
8yCwTqLxqnA4InZVKQBPfGDDfPF9T6AUAf8OvULw/auyXAk6+LC07rRxLYnfd77P
yg1V9CIRiOXmV9XUg+erQN1ihTwsoVhLn9iTMFFeJ1zGbdE1JValUZah/tOJKPYw
SwLhAXCvrh4Wjvmj/TuNQYY4m2aBtNm4AJxyGZEbbt8dwydNt3vRMMHc7/OwIKSj
CZBfn4rnP9Nwulq1K9QaGFSwq2DyPb8v0Mlkrclpbpu58y8hLXLnaQNhd+n/YRgD
Kytdn/Mg+mEiRM4gljz7YkvuQY2PVsvpgHAzIosc0u6rP6z9M/4h3LAmirsiSBkM
6rf0wESKgDsxyH3L0TTTeE/FzQl9BSFsjGIDnCbOsDzk9vHSxzygkvD5VrxtKBdq
wXYkyzOk4aVJ7C4H1isoJV94Vs7TvhWMmm8MBuGafyyMkvD1PHNYBju+FCRCqoHO
xiBCnil51B7yBhCkDg4HhsYDdkHRvaH+SRDu0f+dxRkfmp+WUw1XMw5/GNGoHSz7
XBSnsVYXaZG2S/wTqIIllaAhnqnfYU2UuMhIAGLI/9eQI+jr44E0RrWQrZB6eV5K
AJ2SgB+ap3JyPoRED/F81NY06kxE2fj/ZhTmxLX16gShg+z3jCiDZTIFb7JRDwbV
EWq5FB2VmHIplVkr/deIhyCqZbu4+DYSmdx8rsihNj97CRrkLaUVgeOqoR8GPymT
vcwp5WlCGJm9VkS86bJ/TC8YlgiZjT32e7gSm/Pgm8U+IR6z1jhWxPqb19HRZlL9
oqc3ooeWoQcngwR7XNQxuuqlp+iMfOHYPsX9Czq06HEFWO9nlW5IhYKqeSuvl2NM
gA5hUyKeCF0h7+15Ocrvi+3twdCLVj97JwnOe4KCZgcrazAEq/v05Y5oED1yXwyl
2vXSXNmrWdXywUjoUhlW7f+LggUJCfAvGqKKrpJjFHWkqWdqDv2wRTeIn8UH423w
kXIKpNsEGm1KtcJ5Z06GVMjiMEunUrDKWhdsHV4B5TLn+rQ/M5e8R/FxQEVx8hgL
+ih27CpslQ5wyNKwyVtMi6873tygcy6CRjCSidAVWBKlLwWaA5L3iR70yD0oy455
61XBcP1xgTUbpZdqlB0L9NKGBeAkv3DrH4wk/MDuHEvaO4KObR9lszmDoN6NeRiB
0lKVA6hhxQ2Y29PWOLm36L/bK4LzH+Ywevb0jp+91UeyrOhAQqBBvN7zIW/jLK69
RqzdmXcELpfQj6o/JpZ2eKlS4UG2vPhemXXbGeB1leB+eG5IO9CWILMLjyMdmp4M
glEOHKRUy9jY1obd2AQLjaaCsJQcXJQhoGdB0qwHnUrbCIOcTkLj6NQicnDiAFZ/
HzBH3/oqDVUYgp+wVtd+3i09Wi0ZwSis6SRZwO1EmLzmcS134Jd2EzSoqx1OTFAz
KV7wnqzt3uu0iIgbGBf3JGHx0lUNUNQ5TpDdoDFDXei25huHJt89sGfya06s0zMe
OHKJQWd0/V+0iKam6SsHOeLTx2w+Xt4BqL5XPDXyh6ttLGfQgNOtDYLDf+TglT22
LOFUgfQLa+Jj9hH+7e7TuX0xXUCiRk0+sx6id6GLJ6M9Y7U5ZGcNP4+ns8wWDfwY
ETQfFFahoV0cp71eGlPr3k+tScHupqdstuG7TslEeinyLV7RPrrVDy2YrLcXvNUE
4SgyXGuFpjSeV22HgZHZ1+TiCPMsiErQj1o+jYmcVKkto3FQS24uYtr0CHbVIK3h
P73k8ZDKZZEUc56oVxMSg68F4Ouv8ls7PW5pgS7XS9tBqBdpEFBssU6RRNPvkT9Z
0gIlOQ9Kv2mw9CmOrtnUamjXO92o/lHw5IzbNh4R4OnXJWoZK6p9fWv9KpLsw/ob
xbCScfNm1n5ByYmFSMZM8oFy5bwp42rkVK3O8MJpHJibJZe+qdhwmgHxeMA4TkYd
50J1ptmv4FcK20UY6rhqwcu7hngXrta5waIonfr0qDZCsDG9mH005QIsk9LmwC0I
NQxSQtO3YyXAG9qoAU45svu3wew+pQcbHG6s+h2vx55nTwsB4Dz+0WgsJoCixmnx
CPRewiKrBqJkBduQ8c67s/rc/MQuLrONn0AmvTiQzKjWDzWi4Gn2gKZwgkZYZA5t
cQGXIHQK81ooVuggkgFD3uKTuUOf0Gcu2WWYR8Ee8BzuyhImVI+kvGOPFAnqaU3g
tTa+UKD4Jfnaa2Nhf2wvjrycgcTyc+RAp02DEGn/fLzBQ5X7as0Hv9ohwtrrpssl
T+3lRpAG0hJho37idk8rhuqtGBiUdmbpG4ivOqzkK43eqJn5f4Smwz21P6AIv/OC
HupyuBXqUPSv5Rg5ZBlyyIgSaNfsSn8oXqyk99aSo3iWul/QTnCpYSO0UBFXpHMw
Mw1sBSvOF3MHnczA8K9EX25J2L90uj/6X7/xwrWi+x8njHEHtcvECsQxO+Aq0YTZ
aBK4b4ioIzslOKDRwC8xH3C7X23MRJ6XYXAA47IeXIP30nD4VDD7u7ZJ5tRt+kD8
faWnovFiiI2C8XRAyHJ6r3q60rDf0EtycmQuHHHIzoejdprh8s/my9fq0eR5yRS+
CDhVJ2W9CEeHQ4KDkO6YSPkr61oCUMXvqjzKC2mio30E9ho/fa3DQ8bDrPK6T8/C
iUsp3xMy0O5RXYXX/ovM7eS4Dz0SElYxGuh0yUn7lrsppZsgs5ciCyOnd7WAtL+d
SMniGNJhJIvq2ZTqYh5dnttRM9WjoiVdPPGKM3jMlymhYV84Bxh7E+uzNojfB6sb
1rgOTkMmBHT2eJSnLdIFbwZhNvWM7jBTz+oPQ3RgZ7pcqYGEgj328dLzuLhm7r2a
icYyJVgZ0jGYj386O/WnQHOWkoycqwP+eJ8jFz8hSGFWsE4IYGgOqJNiFRVDxyxs
5fLua9eXW5cyd1MeTY4l9vacHgZBGZzsgVr1sTaAjQyrtLj8xaeS5E4NSbRCCi4D
GSHgWOd4jCRAhCyJ/6rJyO4XI7EfZiBYoVQMKfwf0i8JJT/nsuGUgxixGbNuiMX4
hME76YqWolMSyqfhy+eLfKO7H0y27VdRjOZPWVFIv2k5/eBEogxbk1yhQGgov9nZ
U9ALRcceuAjwvKbOwrRHwueef9doGkRvYWafwArAqljMKYUqBpJlb/Er4336l61T
rmQUkix3tgOXm4E1LNTkM1NBbMO79SgXvIPrbZPnCfBSPSxOBq+hQmnJNahaz+DS
TTnjB/pvcaOZ1sOW2gKLJf4caqLsPT/7Srg4LVM+BvgO1fBMpIDAqs/exYOeru/0
49D2sYpMV9q1E2yyBQhmE/fZid+NHyFGAxsSmk0kaZEazBK9gj8jdB3IUUJ2bFfV
+CdQBgszje4Vl+s3hcxzy2UpbN57bzFcf6Ly7CRbK7Tefaj/TkShPGpAZhgVQx2j
5PF3Rdwnh4Dk0pqJbCoX2E9K9BL0J32iXm42APtGHGJe5AWE2F2p9SwAdsACfUF6
bPVckdCmGkcNoXgC+RBMbXNLpal0UQokR0nW1dYc4B4F/uPWY70O+qAfuFUNSKxY
cZWAZwcVm4JVSzo3j6BwIL8F0/zgupu4yXT1kOP3VFiXYF14WmuMH0w7NEUvrFRe
1B+2D93mpB0ii0noK+2yRZpQjSmHNVnk9iCgeac1hxg2YcxyJLwAcwWVnlpCl2iz
jkutEWoAXfTaLf+KB0yyuXw3MOQAN39nPbauBMMxiAIa5wxb/cnevjssheQ16gkm
2DVN7vfk8RSX5pvhhrOeP76ZiWuNzVF2MF8Nm5jEpWwT/AJDZ3UZzDTngQCBK2k5
cpvWRId7Wz/W/3cr8uJpRNfWFvvDgLNJAx9J0WXpl+sJV2X356Ow+h3idwDmF8eO
7Y7pE3/1VN4Li1T/v1zYDVCviBjP3iFR+QOjjdocRNpMokHdoGf3F1xHQM0ovZ2w
EEZbmktqhkH+R3w6ORvgi+hJTHaBypmi1a9R67i4FngjLEZsyZLbpCoG1VlG/K9C
8Z1UKIsWXUicKYMz3Zk0Bzx13yDPinKp8p8AH/ZnrUUt3JGXPUmk9qEGVnlZEbs3
6CI6Y3tszjE4s3yAypAjCJo6SLGFCZ3xj63cMXlHzjBnEeLgSzQbhUh8iHN8r+4o
pIgQ816DfM4HCZUboW7QzLYk0ZNEwSfwDDgSo30OjeYVuiLTeEllLXqD13AoqpPC
gCnIwmusnp0Ks6g0bKkhEXwbtNvreXh5FPHMWtiEf6ER7DPMMT6HMRo49ZGHWIPr
UiMPakKVxcfhviG6ty9Wak6Hd9rL8k2ZflnFKrYpszM8oqMyBo5HjjcyjBY27W/Q
D8Ar9LImYnRztWPGZAsX133zaG/taZc4N6SIL2HLUlWnwZ7Zq2s9XLoWDFMPxmpR
K48fYW7V2LBjaCrQL+tWnd7OkJlhFR0RZzlBpJrZeQhzfL8PuY26zyfCnb4O6zJU
YX7u+zZmholGlKcIzSVa5s2UazAcOFJoz+2qvn3+SMeg2kVNx8Y+PtoqP1QvXPE1
p/MjpzLQJAb+L43Cr7i4F7MnimbsQ8abo4jOTeTcIOvdHnIbCkhAyKcBqUcb9ryP
RstJAc4EstF4FpgCAA1qr8EHK+Bt3q8Ewy98EU+ncRp9+LOTCHd+R4Qu7M8oAmmx
1zCbtoK95bYbqgfyr6Ryj5ukbK3WLgiHijtSvLFMZR70PK/9n3gnZ0UX8677jCEe
T3nsL0MSD25DmhyweX5IAgSfZxIV1uWePg8sfJXS/h2FR4kIkcpeho4ysnVf8Wm+
01NR2LXYBjvmpjrwr4nEATEYXv6tQcVnVgbZy7zOJC7Atqw4JgAFgCq7iCRIBbfq
0x3bevYq2hybtM3eg3ZJt+ahOIRtztXgCGiW+QRpRlB03T8Ea9aJ+Ptpngq0OT+B
cAhpkU3abyNcbfEJLIK7o0PfJwNBRxolPPWJu/QZk/5ILRaj6X5FUyRXX75Xyn7Y
EMjRx4YCTltjebfFAWXaqTl6+mZefksiKeyRWsCl2eflNhbFBuiA2IgdsUeqsW/J
hM9SfHcZ7qC2KATp/r+F9DJNNyluyozoJS+rbEuz/1Bv/k5Ko6ed2ZZwiTAlROCa
vk4cYM5eBdPLLxNN8CDcLmhOclmaggrLfLEoAwnhKGq4at4pLNoitmioIO/P8xuL
vKHb9qubciUouIjuF+Bea6PULL7o47Yz6bp7ixf1D1f4HJ1sYmfmU0AU9nG/gEEk
WWifmGZg7Z0zHrb0MNENgd2q6IwH77lYI3LAAyfqmnxzO84dYnlIOo42tEjoEcoi
2APFCV+vIamBlsAHASJgS6BmVPablnt/q+FFPdlB9K2sCejQldYV/ObqkxJQ7xgf
vMib5miWCE5ZLlGBsK7KeUsQe3K7Q5P2enkJIF4pBdXUCzDctuxKTDEbAxxTGiUF
VGX3nDkwSRY61KOzXBSwqq/sedEgcROI5l0s8rFrG9QbChMMmxeptr/Ki5rPe5k8
nAlY+sX770jGxAcRW+LXUjzlMOPFEOxHmP6Z/ud16pUfa7xPvp6XMqEiCKMNKJOh
E/VOEe1P8ZcTzJo4QgUBzzTmwkaHeCK2fI8b8eROpiCZ/tXENvflDyyanYET82Se
FQY7r9f91TW1zxBbBH/4jnr3DJs29uAKh0kOLBHLfbL+BTeMF03v0gjVxYR9sTZJ
ck+3jf7Pev2Z1UZ/W0QlKOIl+A2i9OZQA8E8/Fm1i+jzihWeMb/TxkgsJ1TybqrH
SOfLT+sqxYHv+eUhhwu2KTK+CHcO+4+St9+8dfvNZk22+INR3/dssrFCZy6jCGoq
irJiE4433vclJm4DYP6CfRQkB3fZUXWx7yDdceQygqO8eRseF6hdJx983k4HCioL
BLLcbPYxUK2Z+r8L14p2re3eMPMjImQXJW1L2JLaIE4kBArtdUA04FDbonfwHoyT
5KPUE6vGkC0vKRfyGpPM2eK25IMXAyMVRitt+U2Te24lcoYplUXoLmjm5LFWE6tG
d7v97vsAQDtCgOt4MkMdVVnUoHXsw85R9KCwI4wHQ12ivqUVDD9c/vbhTnKGensv
BCBCwJxpAc5gV8IEDJwcr5yO+VColQ6V/HC/8MP/LN3iA6H3syWCIoE+8sPcghL3
jOM5aEEmyFy9Gg56eCVV10pdXWsv89OLmP67QhwsEHjWbi+csRLY9W0IK6Xo++Tp
9LS5EKDmEe2dKJep+ZgCcVWXn5yiNe2Aak3qkGCH7R6DDacbBwas3zIAmxq7/K5S
ta+882xNSn89241fDgFauuUXXGTgrODrHETxtXiiJvP21eA0ZAadyWKZtnJIW3Dc
Ach3fIkrxunudJmcnqXc+fmUVmaFjVVR3lxM2aZ6FHHaVdARrwsqCCMNDQHEb8LR
mmh9OvSjoPit/xGB5hsXEAJqA1PPjhH/T2SKql3FkQcDD92d1NvV7K+FfNFQePvb
8jtfe/8pgx0wbIYglGzOXPff8Wr/tioPpF04uIfo8yFVZolg92dvsnWP3587154w
gC6RNjwbnEvpMxKQaslwUuORZrF0Zh/CvzTp4QsferWlhVWYGls1QXrf54LJgsyn
sbooQN4XAVtkxJPMendkzzpYIWF20qKPORVGmu1+cQolLMTXyzZgqP5VC4ERXFww
cR4GvK2HV78DNXIPMt+8XvxUl2toWUu+A+LivGkkRA/9HFD1x8JpBePX6HAG++Vs
ea3HfcOmFJH8Rq1OZxQJQpbL24VLGWqQyKSjNFoxwYfqMX2HYCERQVh+yNXES+Tn
Lgv6Oa5rWS2I2gQVryq242EmcJtDGKyjcnvEFdzED9PkpWqidjE45koA0Wf5MnIl
zUviiMhacCy6Uq6Oc8NzV1t7tS2czRAvO8cxQvlSTPap2p4v9z7apQ/sEsboNBSH
1xOu7gHBSgaJlCheVkth+FblHVsik1h0AkSGX0steKgdz9Sml5m/IhFo0nNGWWn9
fJQ8N7ApFiGKLaka0RG3kTvWRcNX0xDHMaLJ09PW+HMeOGYz21d7Plq6rXgOVkh+
9xXpekuChXssmN5n6715vMc2UjzmDSPKxZawaEZguF/+nmuxoUFYkkVkSGobGaEj
Z7mVKuzSDDIUEcWFBKbQcX42HKYJH+4BY/T17+EUn0OrmAhEsswoyDTsLW+4LrPH
/4gR7GcsNmaPtM0yad9dt8g4QihmrIIVRudUoCRn29v1wCfiFpQEo6+vDfMaCXBZ
y4PskiBcCpD7KEurh/wfp+HZBuzkcNHwVEdTy9PIkayX7+XD31veglq/dG847Uqh
mhv6h5qJ1dMcXoxhW59Vm0gGPX4oZJgemiXPOL4ulJEgtM+j8DB8P49/NHy20nkQ
AVdRHwwp/NeW9Dqnfwd803By0pG6WfEfuY5hMepwW7qfV3FDdbvs25lpe00gNvLn
DWKiXwP5rWxKbQ9KX0ALPf/aVRtzYrsMd9Xnvo9e7Fab8yA99EMK92GdKHac0/EX
sxPkPkbfIUUDoNKtGsjjpNZLLr/aWSIdVYixtMNfEa820v8rpZEnQPZMKZmJB48D
Osx8gQa/sGnh5RdRInM0O/oEwwXoHwOnbevHdg04zZWbvb2jnshpO4o9OWkF7/Qd
8olbPiih1etShQHGVqUeqH+yS0+ozZ4XQ3kcKyAWrhRre0I3zrkcmIJivY83jrkm
6UdwpY2RjdiPfOH4D4t46aC4DRKuWERnr8uAthY9xizJjvcTdmT2qCzS4DD34LH6
TmmUYJNIpOTuW6zYnvKLy+Am/UC+D8Wr2MXYrbMabKB+z9KdLFiocbojTkJBobfM
cMps0lQvJ3oRPddG/guizslJxVUTxKLncOhjtTH9QiqL+JmL+VADXcH4S7qonilR
DG7EYFIbTTXUTrr+qXfOsnXTcYosNp4+9/LeZD7YdTJsH5nw1wPp0m7Vp6hLHYoy
UmmwFsOjQHN3n/zMDizfw/BZfusZlNpn9AOAXXMKPZcm/8xru5YpSgqifuqO194m
dG5M+1MdoRtn24B1P8ZQR0a0X74DEEzbEugo5JTWTomeXm+JOSOWRPheDPnDq55R
xIUAiSpgpsx5yer0XSZjbfGbcTaNXCtXe9oeOWvjNfRW2V3nH7H5eqcTVObuVJVC
owhNSmzi6g3GZp5RRg+j4UEuN7bRkHHW+gs17acz9UPx5kV7pl5YSHJ4GKUhHj44
HD9r0mmRs8eA2SBR9qDtZGUMDRqbgB4FEzDQ92yCmHlVlrOlKr2xO66dG5fzCetN
B6fy5Fzm73AlIipKuEHvJ4lsPzUczpM3R7h7KeA3pDpXOuTvmxFf2ftUYNEQZ7i1
HEvqYkz+J39wQrLhMyg7MQ134gnWxISvt5ybCo9+1qENps2EHA+me4OC9QfV+DQp
2xSxRMtU0mOOi+YlV3BkS/szVubARjOFplhuFRs/cYKsTYH6XSNzS5ZTeVHfzA6m
MgzjmaiTcrEsP2ueqXhOZAS0bdKS6eWXchUCf5FYIipNwD8eTKkA451b5rQo4Tgd
EgBrsixt2YaF/ZdjaorGNSnwdh/53udlHX5CO4+fXPsHSxd1rwaCCI+ccJqPqMVC
Vc5DtaszNCDo5+vTp5lLFwD50K3AxgjUHmwtbo+fueJ7uA9D7myOvaT//7jpql2i
oVtHpU6ng529wVllNrAGNuSs+Istrxh0YII31xL9ougTZ8ZUGJzSH++1zSCeJszi
j4+OrSe9kzVGpLwstejdjKzUoyji69pRzpZDO0e43p2fgZZovoTaZl1wC1uM2CD6
hMU4HeMcAoyNR9kIAL4TreI96hHhS01FFqPbOYfraaaOCCd90qJwRJ9Gi193wcEC
6irH4AX2cysFBa4ffSQDJsSJ9b6K4qrHx9PuIIdN0XxmsKHZ1BMkEUWbCrkpmVIk
Oi5/4+SThS4loY2HlDKHJvyKzEDaUGbxTOcyJAA5KQfYs6NFqYbN+dXnDVRufIAO
EyWgwzimatEd9AOisNa6wbsRZYh11AOsTmu+0QnlOI96UIyPsrC6vehMkdr0Ozn9
bwxHqjeuB1KYltNVF6DqTgHQby8u4UUcDlxcf+96VUu/X4yHZLwaxbBRXRU7q3ef
C/H8bEFDNMSOgHuavPbkrPAEahrSS1HbdzjgwFzO7fbPqRlxVxN2KSRajN4Ya+ac
AR1HAMWA1hFROKZIy1WJerq7Qbys3EHA8SqwP8CJ1BD1AU2ZDXOVcfLr6aTAC0b2
u6Li59ZLeIWk8uiKvUAAs237+6O51WUJwqAodJTN3AES3t3iDFSJhQD/fC83i6Yz
PBiEKB8eTpzs+xS51HT2eqMQhUoUYbPGfs699Oyh8YSdqHKlUCvABIlZJaxJgTHS
DQjFbAXWsWuywRpQnOdvCDUw1Y89IyF2L8p9wFf+cat91o1NBe5BsyhC+U/kS6HL
kpCR/DSIcumzFGRaTlwM5jrVsXjUkFR0Offu8kzUc6khgBEc9s34I4lxSKJKiKbM
0qS8RXbYwBQuRRiiZCTWCoam1ms6fw4LW4cShLTQOr/I4dxBrAddT2VxsU58En2V
9XhckX/oSolHzh/sz/est2mxfSaJVF00AGEWG9gSN1yYwcbaJMUi3PRgOHZuOUeC
fEHkWUoPnJ/zwYBMAycIUoVv1mxaFC7EmwhuZAUfezdfm7kfy3OadDuHZIch1RBD
P9PdqUnCp1gRu+b7FFLxnWT7n2ROto/vxx4cBQScBwZOXhCSQPkbbclJRfdCcfWq
67HQjbO1tc96F0xEXtOHZLaigKKXH/01vnRCWp+tJTIktYZ5BA66aEFQx3SV+RAL
0H9sqzfZKUVYL5FX6si8+HCtTySu2ThinQ22Iw64wzSA5JJsM2ij69wrgAsGZhqr
6hJhIUxVqm6OCj9jn616GjAbsL2hMHYlo0ygE8Ep+vrhcy5rqgcg4yteoU/QL5PM
rA21cc8gvJjIt3aLCboY31EJ561mBfevKlRpL0H5yO0PkhCCr07Rg3UffHQ3gq7+
yYFO06nv5GhjJQnTUfJfXh4LOXC1/BXE2GzUJYqwnnlmzL1PQaG2Bdfcc6h4SPM5
YyE1DOE3h0lNwdP3UZh4K6w/ragdpJlH7U7DIq6QUiQwGL9RbeLp0vThtLRAI0jf
yTcoQyWn6Ljf75JMT6WPBXHVMqBEw4do9hD+FXfuP/p3G4jaXWjb7CDhe089zuKn
oZSUXukbETJpzBa0AWYwxm7a8AKXzMtzRRkQr7O+jHv+CDDbGo028KjbLlZs1Soo
O/OkrzTu5oAY4BFDTBbywcpUbi1lyWM3c72in2GhWa4Bq1jVOG6OMX1wNAii8aXu
a/ZhQ7KM36nQ/ine0AjfiHBngNavjAcEfA8wWcGaCjBgLCsc7ez86r65lH+329Ko
D2nCWHxMyrhwh8NgRCaA5wvZVvs7x7/lBSKs2gHaCo4eL27MWB/FOWzkuzPOdrFi
zx/a+rZFAmJ5AMw545xhMtYl0nH/5ppC6pwqfrPaBwguwJMksrqIRZHXQ+mgFYoI
eYbW0JPGRMZiyysRJPVquHfpiSpNwjpE1sL84hAh7JRaD2aFvCI6/ut7hUelFVBj
5EKbRvptpOCxvT3ndrXHq29ppT2li+4v/NSzRrMdmIub6ONroOs0XqkRpG32hmLe
MIswcavNzts+5H4W2wS2C9fou8+tWh6zeQ/YR4Ww8jE6TQ+sXmQv1rsJz0ghDqhm
yHP4cJgDHelQBrS9mEmu+RiD9d0GSBWXUJLEUD/DPAnIgZSZCCv0NhTk81KXh34B
KtD0xZRZGUr7ks6EpSU+8e0fvIQqCUwL0ORWAEOQ47oaCCom7z2JCL/0owUU7HR8
Qd1iRHWFtzFoBtKEGaxZQM4i1gAyOFUktaWtFpPql9fHv4qDz7A+YFLrP2xCcytu
fMQpi+f6o2WROH2IWF85OHkuBKATAVvFXANI76P/IzyuPP+RcClwChesV5fRXNKk
boJk/aPdJs1c6PILz8bfzh005KVrU+AwKxvCSmGIk+Gysambt9Y2wzeRMxxkZB6G
LrG4Olk2GsNHoJGa3dtb9BtX6Dt/c3rlNT1N4BVNpqTAeNBfV1hnwj2poUnMG33p
P7utqcK5oaEqGLdAx6g+H63YolhGA4l/y5CdkdjESxWTQf67dlXmWytFl3G5fW6H
EHG2ERWdntvS96sp3xKJUF3GzP0svTgWYmS903FW4++6uHtZzPhWGtdXK2+CETlY
LCfnyddhACy7f8pl69jThU6W4QabDtqYrHVxr+AHtbOTv1hJQXRfFOojNvz7sY86
Bzlg4NOTMnwscXvPgWg31lQdV+dVOXk0ektSttldwHFSnBAthmoYsUOpjTNJm2LQ
VI+LLCFplrq6REcXKOMpfZhjtzq90yIsgYYg14AryVv9NUZdv5LBJlPiYmIt+lTu
3vBrgQn/y5cYFs6dY6mP7GmSPn+daNoJxQkVckXiNEN/4Mdic4P4dn3+LauvOlhS
HfdW2Thq+eWUD9NK60dT8RZ/spXl/IY8+SFDzvJnbx3Jbtki1m1zEltMHLuxxkbn
2VKoQKgJYfRxU8P6CNa1/KgqGkpeYFFSElWq2YxXOres2474LKuPvSVfy50eOpq9
RBxI9/l+IJYlB9vU8T6mgkNhGH1NgJnxsKn0qzGVJ1+hdaySmMdDzowuvuPfRkPE
vaTozboM7VcUE0TEopTzYFEmcEjNU9lo1iUGYl17Ar+m8KSOGvGdlX+EBl3ldirx
alBoSTcK4Od7tDH9P2dqTLPOCtYVHhmhwZVGa+ULkgA51ow9qRYxwfHVl8BwVg/K
Pv5SgSD0WrzzMKs3aiD3nVbzIjmDVpig+fCz7JHy4u4RxRHp1klIU2TKWYHHxsTA
llxsWceg0QhKAdAI7oa7h0oVgJR55v0RIsEaoJ31qkBbDdvBasvzz106jf52Meh0
oQdRL4bqltqwDicCBTa4KkN+vCnl+EvUin6Erp+F1+6cRB4TiW8A5y3OLTO9af+p
yX87K99mxqbxjQWt7pEfvnVFhYBOmVmQB1t7Z5ZnsW7te+Bgbb1m/P+/o+uVH7GL
oPSYuZao/3hnJFnY+vXleM0D9vk7WJNo6Ad0z94gxOXU+8GBx1IOb0YqChz43/0O
IWbAt/SvZtF995tXAXoUgGztiznpQfExmBIlbkC9E8Y23C6PrKz07lYLaymSTiM8
EYH38dh/0pZmf5lXshKl9/s3q9OJxEGPA12gjNGQHYeJ57kvYs6Dd6dqQ9h3AeDl
ues2nUy4sih/BiQxhKmMUSR6X3QyYUhALQm6qTm/4IXNGMP+5LY/PYOffoDv9fH+
8OMgLfEdg+eti0jmdCHaZRuBgvTqcUz0w8JwL7VFEWjaZ0+To+wfuD+G06CBByjd
gxD/xOoFqr9sGwEeVG7Hn/VIJwu3Gh/atstvZdFdr+Xv17gky7ik74stiWtGeVV1
OS7G/iO1CKASMDWnxQWrghUF0YDdKay7lAoP//iFeBphwMx1V1lA0a8TYjweR0WP
nb7XW45efcT8ubn/MMiVy3ZIJAeF8Ia1T/Z3jYabRxqYe+OB3tmIBxxDuHGxY+iG
53P5jADyArH+5nfy1XmRBAXTwtfrVlJaRue+7DEm9h7cyz2O848JH6zTr/daXyCS
wfcf9cRWjAkjcHqslWF0dOJ5lQPazF5WkTqDjRH/SaWXwip8HYt4NzbcyRjrFT5l
VooazuiPtdAhEyfOY1+Pk6yAx2/O2dxQgnwnI9VklrG754/t78fqUyffad7Osl1j
JQKeKk7rWKTjQSrw2rOM6dJEmxA7jSa0DBGEXQBfCWCYUxt04kEiuZx2gvlCEYFb
o5R3UBCpCG5enoJxElnLK0QAcG4zn1lmz91/ZaoUDAtWHh1fnOKnGOuN8EBHkJec
UQoEo/5AD9Akvtr33XPIssxL+eyupfjcxj6uI222MxFfzOwuGro2OWJcg/0b09Vt
sGVi+cexHVE1JmljIl37lSu3X+lZr62OcI6UQbUqGXu7FkKf4aHdPbyfpbDV4LaO
RuVhzyIacbhqn50JJilsHfNEh+h06FfHXHdELKs2mCqDt6XKe7gH+kLixgIwhBt7
K/UaTooVYydR1S9pNLKY2SnTyuHmCod+SwEe3KR0F2YCvZE6ecCi8xX4CLPkaGwS
4CIrwDkoNaElEt93YNmrwzFqFsAr9qicS7snV5I2MmgdqMH/Jzw4BP8uTC34KC8M
zgzOZJ8Lq6uETPourTDnQwWy0+YncypFHpGbGqoQo39Fz4TzClW+cspwKPTo3bxM
s3nZy3hBHeCdhl0jhxiOlrxTuA6hfJ31vi5QzNzWWIpo3RXsfDuf/rmGG6ZPGtme
QEm0doHgEbTbp0PUncM/oopwUHCAP+wwc9HnvDLHRXG6AGuBNgUKpKimNHU3Bijk
CUWCsmmR0nMuPRCvEhh+u+RktoYTnx0lLrVmY3+j+RNpy4BpDf0cBi0Fw1IROPJN
a46v3k1XoBMbB4TJfUf5JTFCN+CZrlmKI0D7iUaIZdKtZB5DLdTTJEG2ZMca1anI
mpvEUa6JYagy1/3JweVe9vqVcQwGg9lDGQ0CoAVzzLKU+XfdaR841zCSJqIMHUzQ
6MG9X4ixCOBj4iZwZQUnGSDuqViIZSR4fx/DXa1NM6aCZj5u/PQiXOB3rTV7NE2Z
w1El5REZOuZfGZ61BclLQENt+ex92L3osz17kI3DKpqtPcYGlwfv+uo05/IR0rOv
BCAyjRtOoPCnduMV/HU7ZFU2kaxfIu/azJzl4Eo2Z5T3Uo+yaVCXcZt1sZ8ID2sr
DqV36TRHR2CCMVlexfIG2SR1uoPZ880Y9YnwPMH09um4ITFxinn28ORsS3GLuG4t
Jf5p+2el+dyG4QahgwvSULnAu5wwNinXNMO4rt6UpqkAbf93t0l4ZuItcp20Vh8l
bFlcYNvvwiB4VqzgJ409hhEUeccrOcp0ePdnCasPwKKD6LhO3JwM5VagIS1nbhkm
/nD+WnDu4sOnirHEzWbcfpu5Gu/gG2WHt9j7AtqGndcpms16inCH/B1mdYIcL3iV
NPIrPhip9jHpdvSjerpvkyjhgMzqosgXVoZQtMFxrEKHsdXoAgqpS5LXK4wDHeYh
OElOBY0zoYMnxZJu+VP/XPSIrjlnJCL+occTz2+xrRpujp3YNppBuZ6vBa0yKhzI
jUf5GctK0zmJYsowL9cL5JRb7zsA2CrKf8uuk0U1JRRFDiew3BVosirByK/cVEig
iOFvLgjViGJ8M2aT2rARwzDF4VdWFsuV+h/CHCJGIgGI02n9kOaG8ITI3np4g/Oy
uk5IjY/9xRXRoJNHK1M8QoXjXHzWT+GwsJwHHw6rBb3v9SGTiLv0LppqGmlrqb2a
qK8gYK9a6W+3xdDw4aiX1QEQNUxrm1OUE3aGsAxYZfUAAO1LjxBjtrqvPO27FNxb
fJ7vUROAwezMwTSxQkuEcEii2wKX23PageYsVWgH9TTptCC9qEftfQbIk72ZZc93
NL62I+Z4MK+qStIwbw91NqhNNtHDWruvmyeKylW6F3l09yaT3r2++HWZOAyKHLvp
OBi2N2WJX7aHSW4Wg/Itb+zUq6GFOaJKeXNIUFFpWZ4YiPlssvtH9S5o5tP7Tzkw
1oGi7UugksB5WPFQW3YMq0wxfnsxSbVGZlQ8GT+9487y5P+1X8f4e8k3hv52n3bY
T7xFb4XAyn2T2JBNq+QAqwSehQDuthQ7iQ6xQn34GkkZxgkg0uab5birb0YANvQk
k9Eummi8aV0urtpJ5Qzd/q4WgMl2pkJBrYfL6ntmr5FbvHiQgzuTAIQ/kzuXdKWG
dkEibU0rPP+27LfiU6LWTwx66bxPM0tiR4DijVOnGQO48EKowMUOe8q3YfidN/2x
STI7ppdIYZu7WosgPGWgXsq0bVyu9dzt/Qp7VXjJj+ci+zNfvk8mfv6KOaaRTxI7
pygfonl1hOKPDtWVGQvBrMxyuxP+WndC0H//DMbe79zX1SC+SVE72qme8AHNCp+G
ohLDUaPg19MjzFUSCS1uPFMuV9rGTw6D/Bv5Z5YoklhZZ5o81gRx+l99V+oD7vkj
5CgkLI9r5a6m0E9NsZ64EzWgUztwhCS6n65T0O/boKQOTLv5i02ULmGlKxZeJzXb
V+RkoShS76fxqBB5axeji6sOp0M46Qe5Mo0Fea/Pwx4CJ1nR3sCKeuMLmidsc5XE
LY8ojXvK4Qo7H4kCBdxrR/SzoxlK0mMsKpxEkE4b2xIrdbatMwqBvidfwo3ab0Sf
lg7pBknvdDQ4R51HbFJiHLEdmem+8zaJXvfLMQmIBlnWeJcb4GcdavfDne7dHAqV
DahvWpjTsbWaXXwHguAt3SEHjp0a3wz/4ZoMFMWZJWq2N/lgsWx6tDbgGTe1JImF
U0PU7hoqnk3BNqH5wJHh6VlX/vd68mV2YUz3tkOypfpqAzaSaoupxvb+C9ilkLW6
Kw2qtBGtlNWyGtJnJTAVdMfejI+4ct73tU2TVtIz4mw1XHfU3n7cSssFw6bzTILF
fA/cofyfbxQctH3TAjUkBxOdNd6Anjde1SzPhgUjl9SEUWtfjLndfigG4+op8MH0
Ny3V6nlM9wqC9tLUcSPsFvYKeBFOCKqndWQGsbRyg1LpYBl9VzRhxxVY79/MT+SB
G6eXWw1iVtsBr5PgTAUg/cSyGPOGZ7ksRCAhnWh0748XKA8bR1wk0hOkMbvc2Dzn
PoNXK0rVwY96M3kViZeRAalElevqLXfiFsGaRl3CaYshDlFRMTssGQHZWhtQWGaE
9YfZwTADZ28f/DRirmFUpDJhVmii6fgUqZnyoAKKEH4pTGElYarnSCIE2loePm1/
LR7SqQb7DZFJ68gacaRtN3ZwEjiyoX7dATVgDXDFedRD0xhirwgFGciEGtTjQT/w
PmxrfrLoZ0cn87sko6+7lCWjp1k3h6m/m0LZ09wqO0b1gSJjmZtCOh4IVh70TTYI
5W8sL+KTRJYPWpC1giEnt7JrBO6B6lzxRDRn/KJ9uHv2pt6sTD6QHpUfyz+281I9
vfX/9Kq6GbVUpnq2Wj65c5NRlUXqBz4w1bP0DSNkzSIf6HWBgNACmNSK+cRROakJ
NRdSGC913wJIZw5cci0gSa5Nw82fnakwOM4zr8H/XEccdqUZUzJizUvdGqIEQNbe
P7N5QwvBn4fXaKgLSTLoQhA2vOxfrhn9byZoI7QUDmN++lVwJnPy2ee8Hn/S4rH4
aw9n8zICz9hRqXDiACWA9K2hLEl0RAsW4F45hSvasSa/5DsCo7I2R729H+87FcLo
XgLzVixvJTLuY9+5Nc1mDGQRPHF6VXktQF0L+3xpVqHLWYg7vvv05hkD1PWpAUNz
NUz+WSmpBs8ATxyp7+5d+nPlz7pu5Wl4wuIlVaEzN+VBHnICD01/Z5iXWcpt8dGM
6j+LrLXp9LQiistZShOV552G+XKJBSl6L1ImNJgKCkwu3SUMRxmQnKfGFfw6nqne
av3WMfGB4t9utg6oZNhn8dPT9bZxejGn+0JR0IOqByCKm+M8Db5JY7aPiMz2aRDO
u95P2M9JMw0rkOWhGSLKau/JdMekwZJIWhjwqn0ko0d/6CzyiX3t92wCxLVwuNln
cMJBAKQHzMyu/whOnT/oItIrVr24s0R3xRebNme5vLr/nNgX7L/U+YfvPvkyChSI
SCyzXmnD936vnATbVWAK/hRvVlHfRpbThAYFzyasinoAv6PHYHPE/aDd9GHep20l
H6bbQ/prcmN8Y2DBIwz1nYXX4GZ96x+epnSM5YchPm0KqmbGeuAcmtwRlk6qKRPg
EcNVCC93DVvELz3SF3A5gaeuwNoxUJLeQJbnyFyfCk3/F7nRJckqxi4zs7PbUffl
M4Ssjf1RYUcNCfDLXK8XiEQq8HvFNfXXeAS36olZ0cB0fhl1JTJaeUl8a0ZYjI+N
yWz/ZPmL9UAXH+NIf89QuaoEXGWOgH89fKBUbLyB/WWq2P6UdAqQ/R4sLdQWUOw3
9zXGFDkXuIYICe7xP9U4ZiL3cAGW0nnE4y3isfRSJTZQRaoWBum/ZxFYBOQ8Tvsy
P5Oeiq2KXZgjmJV5Pg1Xp5dazcYnj2ZaYKiecu/KqxJryJHCbxCOzofZNDgLCB+e
z/quYwxnSJKv7ZLIXv7a3pRaTfRYeX+rcO9Zx2qwUPe5BLvYoNEy/+3wW/ykP9CS
37z3G1jAH5mAFR2UIupWdq3K+FV2y3/iM5PCmsCH3rRGPpgjiGNPGdIkuz+rdnyf
quhmcascbC1RYhStAuWdVl0UaUaO1Mkk8rTt7TNQrNCCrc+PhSzhSmD3xDVIoepd
RSJbziWB8Yxk9t+WN2a9g7HbSivO3F/G6x9tMqdz/DFdZ8LOG/9y1VcEWkfAJ+ZH
JgcWpaacK9HFiWRRWEmiWTFCXYDUERKXyA+s5kbTtbEta3KFUiTN2Rjylan8jXi4
fZwIZp+QH0dimR4HQu8mpgaCeaaXEwBZAKJBFIjtp18JIgnD0UHm6xDb5pPPgtiy
ZdXgfU+Fv0nPbdXqXc+yOtjLgDbzMcvqHTeTJ9EcL5f0sMEDp3LDM4hItEUoQvxE
UlFOwhOIsDJwFctMORSBpdSVU9w62NG9Cf+efNWue/1RuKzk5wKieh4igROZ34rn
lzOXbHXnn9vmwuif3VfUAqQf4DzKWkXeBub7ZRWUm0yfT10VRz58Y87NhvlnvIb4
wsyUycAsoso5lSx2Tl0FaYJdy0lM/r20BIBIII6JtZnnfJrEh25evL6oi9Z7QBEB
cinKZCPiI5kgciK1XOERixJF4r50PsIgT+y/ctwwDUc8Jq8YZWNHt/XV8qPmDvGO
9Fr0iJPN11RUCeG81U/qrFsebTe00WrT2U33ce/7/GLDyPgA/CiGc2NGMQcEkYjo
5IuwQpAcwJMLQ/5Hh8Mzq4BrYf5EPL53dGaU7QlBQY5IPcAmH5k/wJflWjGhebI5
q9flKAiw5jW9POQtcVfF8H1EpExApgL+Caufy63VM3kib0dtz9rnveYvoX0tGgal
FzXgRWcJN2/jfEolVcB2nFBkJM3m05W+AQuLM7jhK2MSLtQEPNSvFA6wWQO75vLW
9lGtm06prvzRMefVzEKAJDpOhkvSnUq5FXws8wC3kR5paj7IaSvf85sDnB3eHmoH
rMRdF4F32EBy+P7sDCOTQ+rN589SSRhZkRP2n+hI9+iXB4WgKPK11FLa73f0NVma
3ZTfdLwJN6I/3hRgBuAoI9GiOMTHLpsgzeYZ7Bb8hpUmpVdciL/MOMF1/76yaN5h
08Zc6zPE8494QIZBzKrkU5WPVDL5SofqGR2ulrh+2YRugaF0w6TY6X+tSZAE7o0U
NeqdslkS21dDoRcG7VQKWJEJNq8mkmg7XCH2EN9jD5yH2XotqbBFsSmE9eWDPXwS
CUUOKn+sK80UU8HhsgBp6J83B/X6xGj5Tf9wQ9EOWkHrcAvr5ta1JoZDmF5HJoNc
woKo3vjloUX1CgceRlMqKgl01ZLj9XoucWY6+gbViea4ZoFpzr8jz0M/1Jjxfofv
3KoTTuSTjfAIdYck+hxwZkISU5vhNTwQlqAiSmSurXQTvFzK5aifUYH6h2bsI7YZ
DUhr0eR5oAwywavR+hoNIN6iCDV03q6+5wj2sS7xEO+GIekCFOS6P/h7FMZeWLiT
ePFOlz+cnEmlCBnxdzPMcNBAs2VL4hmrjBvdm8wQrzxf3p5r25O1BuAfk0sR8dtG
ylypk6SZTTeyxkBIsJiCyoGcWDgCO3erLReBtn4RvKqLtXBaz0feXG7k6aE4Qqll
QfwOO8fpHDdVQPAbsrNQx0UBDfSj9yU/ZdeH2jAffvY2TkPzU8Qib2cFC01Tcwmp
KNXXYpZGVxgGqiwwRa4u1jt+BX7IDDUnocvTWOIHNhOPzE8uXGI5yn5aqSVtPV7A
3b8ZZ6yXul/wIgAKXuT44xWeIdXIDAPu0gpme25tSKvdYvI4U+7YAhbMZb7nkntI
3X89CiwyfE3f0SOVrvuSoy3X6ZpMtpl3KWGpAMWmmBiDaz/tJrhLuXC7VvFiLxnB
JkYhSg2ZM/49I09xhSTzODUXaiHElxliyzJkgc/IU9pylWA57bLNJeY+dKazJF3Q
pAcs5zbFoqYkMm9G4PQls75kNC0u5VeW/qOym5KmeD3lhncbpCU4hjsuup26uVOd
pQUBUpL6d/bzQ9o+8POKDMh8/e5NAF+ayh47IbMdHqfOvMnxsSkbh1Zhbw1aJ/km
P0/BTaHJ1vHlIluAvvkV+pNI36qGQQ/7a9avXYSj0MBuLccTC7pm06YRg4NHi/mQ
KqRDQP9rGQe7QCoSi1mtXMItbLbR98X4limqW6US1uX17f44g0PfBToxS7z7p0uz
4pqPIEBx4O7TUOL2rR0F8CnfQjctMn296ClsYfLWXX6Y6midSzJcvK9axwcMv4Jo
KpxAZEPnMEocH4V6u/IG63ebqCImupWfKWbry9p8k90+8RLNxqR/mNwOlf7KdQRH
9+c18Q4HfSx5+q056ZC1cZXXyAW2L1GhJn9nmDBV0eZlcbN0athmf1p4ooRIsbdn
fXWTNVYRysi37enbHlyTI77kbph0CoxJklbhf/wvkm6VhmTS8gcO6uA+zyF+RO87
EtvetCK010BzSlHOG1RQBT56ni1yZsmxkazXk7HIeZy764HwAN5tf8yOG4mtEXQZ
DK5yqJWYIsyaDB3Avrtpcz6l84XD0Mn0BH5TO6zDhR+Jzy7lEk8erL0blYba5aZv
BvcZ66f61fyWzAtYzF/KsavxHmUh+qtH3Y4ORUG7orsLxTv2TLLLxdIghogHo8vY
Ce06jzsvms3a05OJqKQah0AjznxDJE+9AUu0OhOa0W3aP1lDA6pT5CPFKsst1GIF
qrrmPC0rt/7J+sqaXWhMrf0Q2awFWf8XhelnmRZgJJ6MbfnKvEZFZwLNCzTMNEWI
kKQzV5/bhCxbGvKe7EWcVSIbmHfPkEY5Vtignqdm2XyqMcp4FjaBkoYaZPxAWO4k
J2VI8uuq8YCx+Mk7dJOcwigElfcEvyMxBAW/EyfAxl5EhCrKItNEn6tRJFqb7wg1
fQKw4DnhFSlYMX+2IDnCGPQikIwYXPsafisG7vFpvbLIdJzFd0m5CALcm86ZwJ5l
IaPp8Fo+xrKpE9QC6j6lwfCKxl2bfBWzybGvVQyber7tPSujqsnXyf80+zqEssp7
WG4+L/Qd9mpBr5d+k/75S/CmCmJR5Wfi1IeqyI0bOgMpD9puxr775aM2W2xS05UV
I4bXlRuTCjTghsIulDZSQd+7oInriCf4tgMBMgPuLnTDBFDOjoW3DwQC1zTmUMaC
zmV4vwLwaHYYVVdQaCUP6w7sLJb5rEbpt8tINxAcVwC+x1Gj1MUTFB2Wnhi5Np0c
RqAxsseG61X8Pe0oQzN1+yasJQdF4Fve26BWge+2k+8N4Q+rG47FVF9VqObg9cN8
JS0eKpLIDW/CRJXQVjt0FLo4M53w1RP5NuRFaWGG9sPM9+JAmUS9DgeOHvxfM8UG
zMx1ABSTkmaQXWcUFMbA7t34dxTjaPBK5spzNL7tBOBDOtjaqsqHVp5qlUQUzsVJ
i0n/rcTa0BybRmPy5kOmS6V/EoaSyUjNSVMEmdKC85AaMOyUf4cOTwIsN4rQbx7/
q0jC+LPQ/F6FqcqJBUI2FzUg9M0jTYAcsT2RfPxqetAHtoD6zKCjF9VH7/GE1JHP
RLDGTfvtgqnWe4rm9FTB4QMvvST6GUg92z0rZppykEcSN2KTG8bIBZP8TVgmsI5V
TCvSscKwmb9G5SslAukAgoUJSKNNDMleAzB61fP51O2OkOEJ1c95eAEnHxD/oG0W
aR7w9FLcBAexxkNkAOR1OME5L7+/sofXlGmM13dsbXr+y3jIXKdCtXkBa1oIuIdf
0D5hT5tnSIzLo8t99CG8wOInZjcYGmfyMjfWTX0Ci5bkdan1QRhFjVcnyjEtMrlS
b1+AstqldhxfFSa+W91EDFbQAl8dJSLysMWHM2FnkffpFvmaAfyTfDFDOATYnEe1
miM9QMI6ph8okkq5/xRxoSRSP5YPkhwmsOSaYjXyvVF/f/QsexfPJt+D58vU7/3U
MPOmhwiZsiNyYnCOr9pE57Xd2wklheGVksQ2IdMo3nXYDuonraQxi6uY+11fmyfJ
Cs5Rs5pyH9HzaeymV62Y9i63d3qrkAkJ1nw+e+kas+5D6TcXr2MQTJfcuSBqb+l7
Foa7QcnXQdN9qDRnukdevv0qmeGVjh3CaJaC/EKS9zAB9ZlSu+HcnxrYvAhswzUM
6rU+zzLRQQGDwrLjBr2aK03cmyqrRBP4snTwbBd7FzRPcLuVlVBIN0zaZVIwP0pn
RMyO0MS/JG/7sC1KMPqGhA1n0DTG6SlA6TONPzvwKT1i0d912SBo70VDAotMCK+b
nOXLbAQ6Ty3hs2nDGwwk86E4Oi0eY1BH3ajPILNgvkcH9u7LFjoSdxaB4WnO+Vnv
ITw8XLWrv3g7XB3ZnXzc/lahz/GHMoNkdfqgUHJnTZPjvr5IcXKOLRwzB3Go/AED
PLrhuqVb+tWKoYNv3eYGxKO0sHx8Uki0N8wiBFJ1n3gp2Z++11Xm6y/SdLlaL14P
qG6KpLF9QZh97W2Lz9v2yoiCauPTaCtAu/emUF0P2JZfr+5l93oiWDe25cnvK5Bw
or+e17KHPwThlSa3bAAOyIajznJnMiAHjWEMfq14NYOzTg2ZLub+VLXk3qzYGyCt
DISInDUbjxd/56xhZ7TVqXGkRB5XOyKIF+lewRG4ryJpND5u2XHPml9vXYpOWiN+
BiOi9sJUpAp87YlUUCJfGU9rt6xfSgzgS6O5ctXJYP6jRzQz46DEwu+yCYO6Jp8L
tzOuIuODyRPwl5TM490kcLESsgfHOSyxM3FpnWnf19gzzsDBcr0njoDC5DFrO+an
NvB4WxRghaPl2cb2I+tGjMHLQ/96ioyoH9vOTprtpSg8ZJZ9xAFnVRm6tqwotugh
wf7P5omjFlp7AgGtGrJRcC3ebtBZJa5huAbobEv5Ehi9X8iNGHWYtdEYB04EJSDf
Xt3HJ1Y24ODpUZzGvOyXnHMBv8EfhdUzpaHbLG2R11pbXCyMvx8wb/5M00+NC9rO
Kf/i4OusdXCothRTXla19Bg0a5jJ/rc4hMVR2n5wg31Orr4CDjvwNm/I/W0BH0z4
GfU2cbEBWFCtsoJLsl9PH11eLqecJsEs25xVg4FxXi0cnhfFuRfBigoy2JTGh3gJ
XABa84JyR1LKqmTFIZWdCIHM36bxs1ka58Vv0ydrzpUcl59K42sjltpp+83Q38lX
vZq1oX+9vOxowSIPhRvKhzsRe18xDkosAHaqywGZMLmMwr7Os3bYK2Kr1leVFGkl
7ei3xO44pQ5O2NBXg4ibp5sM87Ts/wuvTP3OUCEds0YfaafdNfcWJLVxtk7lUr1g
pUtk5wVA5V6YcPQzI5bv745RMd/n9av2XkEGAnlSZm4EPanUWR5BlLiaZlWASM3S
5Px5/N+NHP4q/nvgFgEt38H5XpBnLXsMDtOAdSntIExDyRfykLpOg5r9ub/kkiK9
h29/D3fJ/MojIIo3s3fgJkMufi1TtF8hHdZVvRfrcaUbZeR5B0ZOo+PtDUYV9GGH
g3cRm7LUu7n/8cT1m45K5v6uQzF+OtCUPlvOYXTHQ20B0B0PRn8t4SzT/rASM59a
CDA1k9V7mmWW6RIJ82KZg7SEu9r8m7ZPEIPl0tCbamKbqzoRVEOTZCsdeVsMmaad
S9Uan81ANuAf7eBLVcLZBN56v70pHln+a74GfkxOk/yFV7sS+NE+CXOe8M+LUSrV
R7f584KpY+vadkGnlb6ORJHHxa+sOBBMuLJlsWve2PA9g03zFVL00eFszXGJqzN3
vg4VkgKQmndzTrMkzvUovhtXOB1fF4gSYzRRDp/zUSBkIyIuCySoj6QTx1FnGtB/
2IZX8fjKlbqlmXL91YlYt72nCSxa4buRHVHOoG4m9zV68YDkUmvEkFEwU3rNoMJX
/Kdm7NUyT0GP8G1cxxc6FYOz4UkzRVHfBMLDeood7lr9RqzSPKCxqvRzRBpg40J6
nB440dg8w4sQrbH2f/8LyS8dXJdCKZ3tpCqCgGFspQ/O0YnRngr2F+hPxUWSe6G8
GVPnOXe1jlbpIXmzAbdkshCXxvEzIFzGkBbo3qpqwjLV5oKrtdIlIl3oEvb3VXlM
6PE2WuwuETJnPb3PveclAhvQaf9JhzHwD9yX+lO0bedOga4thEBvZqqSM6rgH6IQ
zt4K/x7oxzm4slyT8pKyEz/mx9fcvEWszuQojzPTDe5tSoM4HkTCtCwUKFYruLjG
A1dPi5VZA+wsYt5yv1NtCodMvt7FOL7/ZpphyOHRDLTaYXDlYcHCY0w7CLnSsCGB
On813XEM3mjI3j+g/RlMjUjy/2F2GwcrHsXHy2R3sYzvl30zQZP4MaxI3RGVTYiJ
4aI3fMHvsp+OEaHSI4YlwqV+G8jfNDS767vcWXjqg2iGBsn0GMZ7YFmSYLuoG4Pu
R7Y3wHeJ75mKRpZUrXQih9vuZKnYGEhbG5G+7HL/oFdJPubJXWO+qtF2akCJI6xp
WfNHmk2WpcVm0UiJyEVe2cz4yTvi3vQ2l+WNqQECwK4hwIVJxE3Vd2cRAvufgv3X
Awu6fld7Ej+Mxexj+OpQnqCRJ9NGSaztmkEEeXy+9dVrU6tzpLGuad/UXLTqtJuG
/nn4oqIf2G4x0dj9KMHuUXzJAEt490512kjVNAr6SXpsiicN7RPBd7I4VO9Cs+Ga
bj++RUz+ALuztOKz7lY5P7VH42NG14CCmIT/JQIcpUPYWkD2RHr6GNuq7Osqe/+m
lEz8ELINAlr47MfSjqvC2sMiD/hgJBHjtMd/MpnEcdzSkRTrLoU0qE4UbGBKrMBG
bAeCOvAOw2QmdQurrzJlya5CVBbMCyQ79xP7clUhELh7l5ZKUpIzV9txX37LsCPL
8y+VM0HuohwKvrMjMpc4hKoiRZDPP34prLtKHZAwektVB6Yoi3DrShuiO2LzspTl
7OygPDhBp3wG5WEYi87H7yMbUrFednaDzaR5q7hWtb0mokBTcAA8BZM+SJLIVk6f
+rdOZbiM4Ot1OFLCYL+DQoYepoq2tW5Abv56rId1IXBiQEOY9UCnM8IitGUKmYQw
Y26ErV/4q9XwBRDfo6+hCcvDLGFN+VLhs49yEi4KLClhwlMson3QL96VTuuHQ/cL
GxhFeHPHsUXqtq/sG/abNIpP6Am2sg+9Xc6aoCUY61Vl8hgaiwTpPPUjJymeJaXp
ckISxlzrRvMXI4bQsB7lQl9nQKcXchtTiakstZYkRYXobYK8MCK7ePgVMBPEmYu4
/5M0IAH3tMotyR0SpMZzdG1Ech7WdZlP/ItKGNsSXIxVGAvHD+wg2CvHWBlzTJ59
QWF6oTQ6l6WBRsWxkWIgHcTRSMAbjbrm7rwIdTUbhnF9/3ZfwAlQygiH4oIx+F3X
KByY4J1N29JdapQTR7VE6TmzLNi+6GbYHkyncFHhid0gy+5WgGWc/CHqRSxTjECJ
1VjCcCWk58RtGOuikcZ2+Y4bFHBJOhOt0tfRhV3hhPjSiySVUw7GDqVnk6X2TKD8
g4DLvkI4P4ZDLcCxeLCcgVa3gNuxAhKSqjOxCL27fSbrWD3JAN2mYdMmnPBjFqo+
bzeI29HNvdJpzuwKR5iS+Gtr2CPh6R76euUWDAeXxXOg2s6EzBdg1aUrrcYRCOI4
zVqh7SzmO9aedjs72vrx+vpvgO2PezXs/Rb17OmbgM7wyoXRlUu92Mvw3LKqYLfr
vOreS3SSTMPcOmkSuXVsCr8d2+jx7blP0WcSu8iO/89QQgU7/8VR62r20QhU3YuC
9PY8HnnKDm/TLF78bKY57CtXNGzknoUXTzWzqgJ5uuvkNoTMPfZGcQnmqVzP2zU2
6eUYeL7FtybuD1JKzqcx78PBobnY9r38oaYb6u52Qkeo8AI1SfUNKC+kPGrVYrvQ
7ENUuMkr88wfAbDeN9hG5tEC3q8yJ/7E4sZdDNa1Qm/95twnDtw7vknHLH6X0Riz
xGI/h6X4CNVMpLCh+Ml+WKtp5KO6lM8/4Sw8fQtCqmYIclTPWl6CFoTNA6YO/rt5
LliQIS3YTZZ6gawXJQlWvB/Oz2W6lf2scizTMa9+hackrYJbvLk5ZIjTf2JuNzM8
oaidkKHZpiF/P5VJHG5NcNWp7Xut0g2U8J8Vsh1CCqRcN1s7iCOFJfCy/q/tRUgG
i5qYFfsDmAHxTkRYEZjPTCXjQ0UiKgovHZuwhDJ78xQ+5+hCrF8UHjcVmtJObrgp
+rnvBrsOHdMOOvOmRMUZ0s7t/p4LsQulsnU4AKy65tiLE7mHhjMG6peBjGgs/i24
pwqhe+hfOMbSNzJL7mVwjeZrjezl1hTYXdkk9e20GlIJn/2pOf+bDMxYJvSLBp3c
ceFyrlPX/4zJEFISEQ91dUHZdqcPuxl2CKqj4nAN8oty1aL6I5ypw7sNqEF7a9rq
+R88NRW/KVqO3Nh2s2myoiuAn/Ab6RTrETywgZtIu9YBV5hIYlfgORt+Nvarx8aG
L0xD/dxX3jPaqJXYBBn/Oa8qZiZmiGw1eIvc2AJHLoOaE7pEdj/FKYXih7DhCBBD
8x4E/8Fb+NVfIadZ7RG1mRKH/iE4E+RfbHmqVaaDLET1eu4CEa52hedRGDGIbGst
ASqYdSGS94lu1hx+J0hNiQOD+X0h3lReJqa+bgfJVs6x42VxJqd03FlCerAmUzAU
n/UgDZtrqSLtCVnz/OJdMCublm+ldcMP9rd0bGgHiYK5Z3Lb2cYt2UlMp0MtVTbS
j/YxTzsxaCA7T0Ruy/ZkHNCNKlD/c12XLR6tmxIA4DFFUWDjJ3bE81v6/FiVuIvo
WDBVhL7KRwrzc4n20k48kDGraHW9I7TE091VEIUdO8uGJCetRirawfMIEPBP7PL7
wZvoMVavm872GUOr8Og3nn7j/gbQYZ4uioJWYtUDNnm3M6Mt050QGv7xjO6jH8ua
5er9ohQMOvXtnlTmrcNNH922uPxQjB6McuXesKv8NAx9IbKBhgGU440sL/BGVOMA
l6u2ilPN2K55eRuQK+IaDfOmhHoVo7URI+htBnZcM4JLX/diVU/w026WbnHuvFsK
Pf8VS9D/1J4GhIAndoApJmQgNC/fcKEYs6Khql7/tMLeTuvy4lZIh8iXwLzGPUBZ
k3RYhozKsKhzE+bqM+2Mdl/sFSjCw4nMpMmw801X9fJUrF2noervdwGjQX+4CF8s
vnHZaPKbGGdTNMJB4vcCmtay/j4dX7XhX9CsL4i6ax62TKmL+K2bfjTml+JjH2VH
d7t6L8K9GLhkE+8/vXHxjT5N3Go+y0UApZDEd4eybVXjrxvDClZ6WWmPg9lPmsBM
weSu5mHHWHnYJGhtr6rIpLOrgHu2GELAD03YvPb4dGjIp7JjV2S7EW4pbJzgKBG0
sgZJH4Fe0yoZ78sD6At4q5TC2ylB2GXyPpLcVGC/z5DzCGLWe9cTQy+fsxAMt4nZ
I6st3k2sXhsvKv9BguRypNyMVhtvcl2JoBwyv2jEwqyADtcM4a64I+ozqvXkIOq1
sX09icFpi12o42iyeLofVrxZ3MIH/jr+n3Un4jCYV7Toqg4IIcVCjFEhshbneFKI
rGRSdH8fvY975awrwGH42zvTyv66nQhfcXAfojI8ASnRQDR3BV7Xxs2ykOQNhGM9
RDhDghMJ4Axtg6qKRc4YQ5UMpXbOLEqrX7fkb9GdLlx9Es3bjPyb6ws/7zgGx+19
LtffUgvlzgVRhdd9+Zr8JolQAPoB2l2RhYpgwKtXYea5s6yie9/IfMD0uZoFnu2B
H943Vj9KRhu7IDmghRa6uveVso5YaAO+Ct2g/4bcgK3xMqLLQEjqNUW9YkzHar3h
zCtcdpf0xCwOGH3vZ8cIb6Kr86WkIjdqbCsFWwh/WW1l3ki5PE857MabGx48h9En
ceceay9pVbca0MhXbfDlTnGoxi8YukvyMjqj8eKI1SzrTDgl/zaEqcd8m4jDbQPx
MItXgyIxgvdTE6uu81OMrL9SWaGks4yix5U4i5R0dy94IHFLrPa4TJq6tGaXmMOD
QLG06VR3chWekNM76k2ZovbmRVpRgEqjnieHMPyrINtrHgl6NvXoAh7wGNj8Qpiu
TzcZPqTvGvcs6SQfZrOQRbEONUC+SRFHU6bIZb9kX/53vk2eGpVVFU3bRTb1vbOt
WBIdnPkbFtcfSUudnR/VxL8QiSPMy9dcbm3Is3je8Q5qjtk7QnwTI5Fv1tMmtO4J
Wuw1oct81nQ/1uGAJkA2K+LVyWkSqC8Ai4FM+8odvvT28I+NmsCGN8zP5o1ZlU+j
JZfR2TSIHPI/mT1yenoF5fkAhgEmF22H9nhgttpFvTv/eVudAOIUK9TOc+bao3CJ
fKT26TD0h8jIyqdzoRatIwEbcNgdOMn5Jen5PF91hVVshe9xZsuFj4LJFAU7g+hz
C9M5WwzgDGzIhgbPYdBsrAJIuf9HdlzOJ8aW/vyV83p1E3yFICBs4Vt0UjwOgX1H
mnWjwVuSke5qmsQOt2c8Uq/pmk8gcpin2q7ni/7yj8X6hbQXdXZtxrosEWynmmtM
LDQ/HpKeMnqWEJys4i8GwrcJCIFSYuIDkMuPD0tRs/ZOiz9uuOxalFW5sYgV3VXC
1EkY6N75uKPPZylREm5DV2Qc/dfrRk/y1/PXSGLlzBuVAWO6EvDFzSzK3dODenzy
Qw47wb0f2+MyyBexUhjXsYtq/c7t5LaGj5yHoXp0afcxf9m+WusDfY87+Md+Vja2
Y0wyqyk0lsHWEykY1xzjbbrfABC42RdekHCKg/9BpTwOLeNn+VTJ7w4nfoQ6dC9v
i2uoS0hbmaTnxO4BeN+DHXfTsGEdznwbdQcWhoLA9otFO/r+cXIoBAGl3TukBIjq
CXQl4pGMr31nMhpT1CFP5sY8o9oK0F/ue2c8tWOBGDAy4ofvoxnRJYSK6NkHKMO/
9lA8/HneoBbrjecRzeeclaBps2bdOU44N4u+SBYg64eemueAL9sMLF2wnYRW+rT7
5kVdtxhiO+agkes8mrCyJYZTt5GW4vm+eo2yJh1UItuHhVdfvftNnSaAuuR1LBwC
YmSvFUb0510trQ42giW0EqtGr7CmxHJBIQauV8RdhldAZQeWVmFzCAICD5QV36JA
KM9VbW5eyzFm3OHfABdS5qjoa9MpXTf028EHanF/NId5veEHV/eStKA/I2bvhf5d
XFIDooLUpEkBYmNFgNFEZCbkxy7veYyFgXq257Ozwf0Wq+r1Gme6O0S1wfHCothf
QohdPTiGnanptCNLCCgBWzTvVnQRPHpbOintA5MCN/aXup2crJ3P5cPjFQK87ni/
qBnzcuO84ELHHd3dFof7IcipQLZYksolx0XxNVkOH3GqN//Dn8gxeK9rMy1IN/Zp
+TrKB1pMHNBbn3pcGS01nd1+D6ZQe85tipPBKkU6rq1s+TTUcr8ZKG27sIEun2dI
8Z/cpaBNDKWxejTKKxa4WBwbBHKupyoIylBp8wQ9KYtOoq9wwfw5eEDX7GpysFPq
D8jxXyUcpZ8kN4xEgVjrq8gloljU1t+vwBilsMzDm8yTFzz/aEjz/uGIMfMi0EiP
G1/XVVjfpNVZG+AZS+WgzstZ5L505XSsX2KdQUpgsIhiG99EpZBRh9Qe3gBdlpVV
UsaLaSI/f8Qj0retpuN4BU0CiA4GvS91gagpLREtUvoNBZCZhVg6U9xDTbKNUnSy
zpuFTem4mvQKWrWqN0/m16jfFByMO/WrUD0LZuKh0YjefJFasbEmmHypHbPQmbeH
hlZzgTqLkgGUzxbfbs6D/JaNYkzWQ0B4MaoK4b4kgtPNQi42PbJ55tvOnQrzi0x7
CVAlEbzqrM5fOpo+Y3GRqQ8ZVgZLHUAIY9WlXrSr58VJBEqJX577Hl2B3OB4GR+y
JszTi4mCoRm5UYK62BmtOmcXteBtAquZ8qC/3yo2kOzeNBq77fEeSVp+cZLtWRAP
hg7rfDwXALECyIHR5TXtDHfToYKCd4PJhDyX+N2ebmGfWcy6qXymrAeJ9k3I87Dn
a2/4O6sTOh2JfUJ5j9spJTrXOtlrajzansZKD+M7OUHbge0xN07ivZ4wDlE3tYJF
KBAUp15XmhBxfAFEy0iLstEXFz1XfXu2A0wLLtEb481MokdAL8gyrzPhjPd5CInl
WyPb8quIUM+gxYKi3mgcf5kAsujJRfEbHyCvUL+YdbGiPy18qo33kjShCtx+mS9S
rMVLznJMk9oFiPrT4PwGPutosW1SMqSA/YGrA4N084FWJLTDkOhm37ixCoMQnzNy
aSv1HpjKJ48YR5nZtxqsIkRwPXXPEKTPgVRt4/RflZvCigjy7LfIj4IN/AT93Otv
ljHxL77vPtJzbpgc15NUpKyn8tv+pTUhwdM5PHj6s4i7a3tRfN6hg3ekUhcnXpKH
CH+U4gSEvoYrBXcIDlWwxKbqfZO8McooNcyJ2vOp57EjwTTsEa7uK1p71qO7qxYd
LqjjGoIAEWAQJBtqw1/i0u+F715Ld93vyQyQh/2oO1Ud+ceUKY1ExExSmLz0kelj
dsLC6ZRmoRYzqXWb/cxbLHQ1pupbhBbmcwUCaZwHv8Jz5awowQvsO3N47PEnWYvG
UFeSgPMi0sLcsiQageseZefX6DUgepC68jPE+mjgnfxszt4wOLC3DqjkHVnqS6N1
3kFQ1iXP9Ih9K7BDvQ75s2Yxy4sCcvBm0WWLFHY8eq6EvZHPCadtXTMA0tURUhD/
KVq6Ruz4lxjOYuVhORPujl4lgn4qEKXHrHf4I8bXzCDyYuFyMoVg5242tNTyEUJE
XypwOakO4xQ5XLDfmZqT5dcNy/AQNdLrItn/H7A3yzbDmMRgJpit0+U3/aZ9/hRK
3d8Zhm1QZFNepT4LLDpWimTzuTRavatzWNhRLa34nQJu5f1FIXkhwd2JTsF7sa7U
Ntdrsn7r3yPFYMGATtunuhWtet2kJIBO+H2X37vfw9sNQMXDJkoYr5bF7pC+QgJ3
5wV0GutrdVlUoHXkMuABHXC57MjlZGUmMFZbvUL012l1snOodkQJhneRi+vyHb+X
xcUqQsgT4UCfw2aCc2fS5X0IgKhVg8AbbH0GAzyQ+ORqKNQRfrpHAwqlsLQcgs0a
TL0lOGuFn3mZQvaT4+8S0yZhoXRykxG7gFn5iorS14kHpHuJcgkztAGp1K0DLLOU
QCegAEENTLyaPkV0OcG665Iflng0VVYpcljgM73tPesqu2mht1UWjTTFndgo6aZh
Omn7k0QB+Fmuo3OCvragxvyWcjuzFt45xZbciG89jrfl683Em4C6rzFPeVJEYRxM
CGB3MRmcIb/pLTFeoW1DdAdjEzsMGRlKLwpDnwCPZbgafL3gF+LUrk5qDrv4cUyc
+8D155yPL7f4Aw8VEr/YHdcdRMqYqt3KE48cQgE8581G8qMm7OJr+D0imezo/N/v
RY8iaQPd0zY+WqvAyjFkHXpCzVy/3FMGrBiP8KCy4iyLYAbRJ/MMoIZg6C0t725I
9wZNOfL1TO2wdAgRqurU55fksN25/2dHZgFnoLPQkVnY9hjyYUiuPNhs+g/+nYkN
zOWHy21qOmivbShqYVSlDXJ2utFqnp3de20aV2BBltoK17rmBD9kCeuXWYB4qfaI
gnUlg8sh6z9cLkes5uBbOqTXgqVMf2kVjmAKt/Vu23od3UCwFQnflE6zfhiea6Cm
eYuJ7LlIoQk8hO99bH23ERL3JO48+z8etTGVo4VlqwTgrZ48sUaCYLqEKVzQMbv9
4Efu+vxbZZljL47yUwmPtyGJfgvvmKkrCpne9SDjmBiAwkLZPowOSZ1d8ofwLPkW
yEyqsfM+3aUosX2GccNtEhq6ItdKbybmKP2DSji+ZU0oUwh2KtpJU7T+eQIaDaok
gpPXzAmBVDsIKtd407DNyFT0Q+I73ZOh9OIRNhqpx72naYlbYZblEVdtVnx6T+Jd
CUx+fAYSA9eRk8jIfGhSN750gf2j+ZhoWFYfbWZfoyvOd0UX+UQMxFWD698ypJ94
O4jdS87F6AVjL4SJGzAjA2EN1+7wi8bi3HH/B3yCli0dyyyNH+lpERLqkGPvRNCh
T55EeKhjB1JWMvpTE9vCd6c2U71wjfrIOECpjkYiHFNczL/AP5R/aSArzD7STgdH
Zdvo8YeULvIH2cK6vQ92X0nwzatQCy2cRbuxbJzy/3eHkugIZEkoPnWNCP6ztqFQ
dEqZVprjcFmTzKsIPZCHmfVIVijWr71rHoq+AGJJ7PyjdrF0ikcfojxup4PVxtqf
6fmGpnlcJmSA4+0v39V22PM671Cqaei4oIXYA8sCmiZA3YSb6sAl1LALUSHNv0AQ
DIthyYx0k6iH0weM+Cuar62qPiCYaxIh6zm9gcbVfHDbgYxDlc7hrjRfQXsXTR51
HDTT+7VLD1h/E7VeJrjj2FbWpxF5XfoiNX96l/6rCmD+tzYPYAQXLQG2ppnmQGpa
60gUj65rQyKl1SHfraURrVoRn9Uz5PbjD0ztNIkM7nLnikU5y9TRO7XJUsjRlqZW
kl32xalv9Ij+Lg2hCndcbZjExwfWpApXR7gkogi2acLo/hI32es05lS46d7knbjS
+SDdxX0tmKFedxnA5RyB5B4Y11WgtrJXgjbyLk+WoOLJSyJ60YeSP0JKHEW1Y53/
F2MWtg1877tI+1DSrXbdUrFRoCU4tGp7uQ5jR+oMkcUnlAI91o/WPOCw98Kclk3b
NxjEd1di5VP7jACdcLERqlqQkqtZwp9tSZWM1J+KY0zbdEJSQeOzM7ZdllmCGqYn
Z1XDm7YPw7bsZIy/FK1qiZQikcf94138H7IkX6Zezx6iXQW4DbGyjtE6HNLoRDe2
3Oq3qx1pp1U/MgmV81/QS0TrHoLdwO+p3B2lh13P7nSnDaKUlCLAW0EzGOgbbiUU
TPK3THodroaoCFbNCzZVdO1DlSdIuIUDd901Zw2BLyVUo3lKDT+LJXMjGJwfMckL
lhGEZNThVhKkiLbCpVQ+bzUsp/Gt7yl8+Jcs7lD/NO6XMEyi32LCbY3L+NGatXgG
VUG+l1snflSlmpUkfWi6f2bTLU3yjwbB1RYDjvfjDWSrl3/7jMGyO2X/MfGyxQCZ
gTE2ecEZl8AuuCsonsRSRH9RPoGThSEBKAxaFX7fZpbzvoVBOuFr8VEk0IlEgDq3
aGOC/d+biomBDvU+h9+nVt9a/7tHU2JcBUiqs+Mf+k69TQSzYNeylVDIvD3eUT2Q
iCStaYa6v2l8PYKmXZylXb2D3D/aRLz0FWEprotoYUBJKkCnjTlrbgn1mJb2NIXb
R8gTPEC1lOjvOYGBVwJbzE1oHxj+BKl0EbfZXE1Gc4QN2wA8fQTLHF+16pjCtUMy
24EtPFlb0HfDtK3pVuZG2FqKHcRQ/5vAxMYZ/wIh/HKaLf3i56E9bHKITitDY1va
h4lAAUkC0zsUaS/UyFpmegTw/dC5oaJScCYrEwXhFgrY/tPcq7eKOSyOKAM7Odtq
Y+snBoBvlcCvIitrjVTDOiVVS6UIbJ449GfHZVu4Q+olYimPTYGG/yG3lyy2WqXD
YuN/ZgOI30gm8bognuBf6/0TxkZM8hVoAYqmpqWgl+8GBj4jFfHBgTjlt5GeiSeX
S0A3uinveMg5uDaUbFRh/wtKuBMd+n62vg2XcXSvzKKfYEPizPuqrt0In736gFb7
oXRtt8lwsERsI5R9bGCP5eFp5uVMItxJx81zS8KMkVRGfOw+VxCd3VhshRJzioNC
MvMdB28P5BImhrX7o1Y5lVkfa9o8FlNBhOiNgftocpmNBDJWbKUJU5iMaYNz+nDy
BlJRzFJnu6Bxx78YdsMS+KxzBV3kyyhWUWyc1LVYz65b1XmXMpc/yDSwUh8KV8Y7
oyelwmsJjcKc6b6da5xOSsR4sFT8J6lPhpr4Pe6q7OgJkgu9OX4QVd9NCDUfGaRr
GxsPY5HV2evh5wzgDiV/ovxSvExupW5ZgjrYc1XgriQ8hxyzjuwq4f4CR1+kVoTg
rteax39/IX03YYpu3grFE+JueMXQDqpQi+XoUFj13g1PPdGfk+iUVGlhxizelaGz
Xb1pR0wR4Ly6f6vUSy55BbbM9V5eQxS4jNZ/X7yJbxFD06LqLFdssdNJUjuPsD1Z
0NlsBPxR1kLv5B0W6a7IplW2LBsg0bqIqU6poWquY+c5JxEIcb5cqlmZ2xM1brQA
dq+3UXRWz/YhM9JBweHck/WMOx1NEufY5w4EKm+4IwXUiHohC11CrZwNPUMnEh6y
a8oHJRyNG3qO1SEp6aei4o8PpGh4VrkCNuJFL8OITZg6LyYkIPzSetSoZpvahL7V
84I84TjgzE3qbC50hgrntQ1Gv8KP+J1m1iLTWrusEzbDyFL7XLhSmsMgLhb4JbVB
LoIG9fiWdcw937VwgojgD+5LocivQxFR0w4ChCqKA5/G7d5mmJvMIiUS+DhWZmNw
FihY8wiOjiiqYL60kFxhaWcnVZz7G0OA3vmT+1ohyTKcaYHK5G+3mJtRba5aNXMx
8N4x+r0UkJHBlA9m26ly/tiN0E6bNVQUg8o8y6+Hc4EgjSphRymchOiHNeWqSdPa
e8WC3/xzOWISGyWpWRI7jnrXb2P37grefm34UcH+FUCbXSWx9X3IP/KkFWyZvqG2
GikkNxipw6JSe9v2nTRrUkdZ4o4ZHdtNYY1yyPtx1cfjujw+YUuPUN3g82VnoAE5
/uedgb4z1gwK043cwMbYsYfEw9bWSrx6qATD70NPHmVcFX/Gr6mJg8TxLLbQ1IZQ
EhgnaQ54BoW9PzOlUSsOyo44dHDLVhywXUb3qgi3NqmBGKPC700wWv2ZFoJRNGC+
pMhtD1/L5tIhgKIuB0XP4MVT6DBaE9q11ia/SIvOHxowkWKMNeUCgL+3r1sWV9tW
i5SMjfJNv8HXnA8bK5JXZ/OVRmnW9pngB0qMx3+0TMKIPebejJ4GfcRp+3rJplyI
gn1GIhfo5uM9iQNRJAW+3XatXV7zOzYzTMiHDKVUOcc8CxnxCTzhaLkAFqn4FGt/
lCHHo5aGBGIsB+vC4KlDLrip9JnttQPhMiov1OEV07qgNci+6ch86D53wt2XarE4
O7AXA7H2cFH9UCBKBXhOOMlJ7bdKY3HAhFAXCI/TtU0ZO8EAOtyT0ir6FDKZNvze
tWVLo5K2MMZGgGxdWa31Diza3ct0u6CSfhH3x5RoLQICd6ma/sHKresFS3S5o9uY
4jpX9J7pUGTL2AOdLwOkO9KdbpAI/J3L+ZEasO8x40IRwZMXiksEj3mm43FhhMdU
y+qBeaKCiIoO0c5S9FIbVHyy724FAzUA3/HMJlKT+v9ke+M2zZh3vYcjXAIIbiYu
y5q3J8RPsoLwr+orVFi0lg6ybYehnw7U76EkQoUW1pNW5fMVw0apLcqpRLbY4WRk
qXa2UDHOQZ4UX1essm5iz0IuYAeMv8hfSdwmU8hYqBWvEU0LZvmtMUKEvwOqP620
PlAQaqX18Uh9vIrRxnNoKPLoZzR4Z1BlyzBYLxpLavvzfczkvGQJS5dWNsZ+uuYQ
MrLG455HUSiZRD0ZYq5LKu6uS3dCqy7x5JFEUAXNggew8LRuwiyaDeRgdqjkV/6n
toOHgvzo6OG2XPn3Lxr+e3MQ5wpDWLJbg0bF+mWdTHkQX3HxLUnYe8n1lg1MAfzb
d0JrZmlwnK2oCXfRAme1qcgG7y5f7V4AQhooavRu+ChCpscpoZAIGFJPQQoZJAUn
C6yF1+LErShf2liLRwnonewa4NaGtkktxc7nUwGxMgDAOBqU8ZTb7l31dJtWx0vy
mjmYUAVxOHzqBWm6oECLLO6V26D3r2FXwIvnE/vhmAQp3cZWU7ckYdnCv/ALrd2u
T1VX5hdsTB4CK7dUm65sl6JS4xkJbIvWxZMkEmirvKMfKBQl2044KP7k6j092RmI
UCCJ+0aX48isdeuwiMQ6KCIovkLg4bz2WsLQXqbEt2CDBhjt7om+iinqMesSBAts
c6FsVyTDdPujJzf9hoQDNn9XsNICc7q5fepUu+XnGncChSstW48gWGloVsxIh2pE
XXF8mJLzMDJ+PqhTbXY3BYisVWOxlm+z79nDTG1kr0c3ILAyP71LsySUPT/EeMp6
uTNop9eRhG5CA+/CLf2uw7fnJo+Sz+CFtM7XovCai0SAsO7dcNX0z1DPsqqS6pIc
/IVbVjtybpEuwtEtLc/nXcuUHff9ARMAzaF+rhgI/bTSgNyqLtUBDLbpYVQrWIgf
/Ehw49bWcM4+Ocae/yErat0eMHIZCSgdkY0/x73AOuHhfmzXopOADTXVh+FntEAn
U2DG/aNViwPGEQYslpDDdrn38tIojxOGc98h3Ziyt6BLeoXfvjBuf68TCBdHiyIr
p89bgzIxBxv8kIaSp5xJqz16cGgCnYi//lDjPDQ3rTbF3omssDI/T158tmAQANuZ
4R13H6Ou/OfkrifwnnnXxEWd/jkxv9FmnF5B7AHAxPDpZugVVxiaPzjxu/h2GriF
8f8F4HQlvjBeCIyWioZlu3qbaGhXFn1Z0L7Je3bnthyTLGgUEv1tU3Mws1tNMkF4
rHqbI2kRRjsJnh6nNJ5U0Yl020garHVyBiKGFJu5NfLwefP6oX9HpEGuWv20HAPt
UFP+EI+7CfZlU4DKtZvnl0hslLZMEPxBQOCvieqELESwVthjEHmxoFn+CD5p+f/v
zUxMx6jj6bdH53XcO/vc04gifmFF4zUgNce9plasPxZ68L7IoxBHuP4LZ5GRDlCX
Snx6pZHcvc1udhCKpCKdJBQWEhzdxQa2ko4hVhBsC9brq9yxmKK7VjtZflty31/t
Frw7/5FrURij+9LaW+MjVeLtawp1byg8ld9pybeaI1N5+eaG7AlBNbGGQ5gvMasT
jA9x2crmEp+e/PBosk7b28WAfj1gJg4SL756t+nAAK2cKE4+dbu3XPyqeOvvbie1
jC4UVBo12WzpcKpQzhwCrZ9Z1Abv30ucbotPNfEquyWjTb6Og7LN7UYKPoAQlRLI
fDViZ/d+OJ1wmLEQt0HfznRnBWqWm+/5n4kHF2oYC7rnZgwa07uq6Chbzv+WgR2K
aPCeAHFly3cHediwUb6kokUofXEgw0QjXOq/aMIGyimLU+wjI4kj3fV15ixnZrSC
2qVAYuUToUpv6aPigsQL21hGrLyzgQjskU6AC77duy+cTw1aNVl5fvXlXJr33AT+
6PF0I9X8rnquAwaQpG1kRClmiIuo69U9Md1kiaT5Q/GIILbrMjFqpcW03kU3KBCk
yQzigW1RbE4IioiODx3SuabqNGXQBLsIacEiCJCXxVn2+sXClUFjEHxopD/6CrS8
t92nVm56ORsoIEKTCRA2AYZmpBrzUd5D2IHpxNk5pBfiogInJQX4OtafFMDRJmPM
ryqsxNfPxGRsxCo834q6FudrBzDAgnC9YTNagS4JMQkY3MH6JXzw4IwS/SttPueu
FustnmaUD6dh4nINnOZPfkBgLOo/pnGSSX5s3pZ1V6aVF+DuZywow20Wdz4+cQzF
tuoXNAK8znN5OH0Rz2xsL402b+dDzsGWAcBAznpcEKGNzOTA9YPU/vhaXIWuHKd9
+0RnV1HAQy0oNtIdK7i0Lv/6m1Mpfh1JqaU3o+UQQonRH51Kd97Jw55rx1lM3D50
Dx3ouq9coP0xUP9gUirrtVCX7V3kLzXSe/OxJ2KsKhZEYar7QOd8zN7zRTKZZXCx
VhbbQGgkc8u15mpav1ZtQFNEAqCypbu+cDHx7klGa2ieHaieL11dy5U3xNj2HGwO
Tm6ihT3NZyd9Sm+GSbTkPtryzL0NZ4lVhhlx1wXChrfUonvfNralpmIoYwicpCJG
aE9UMydn1hvyVXpI9lEH251k+672pXwJB8SBqc8oVgt2yXfg7tUtctelubYkvoU5
8FwNdVrinwLJTfPu8PPbHgmp2jW4/swBHFPktMWuOSXR3cXCopeqM1jckUxWTa4F
uUaX5Pw4EpZMEs3O8R6vveXARzBh92LK4n4xlTbxu05v5s8WjHwvR96DOrEgDqiD
dZ+xqWJYExlqM7+sTDMwhJ5mxxn1lT0oYcItmfR3LXLzs9RRb+qjDytzdUzH/NOl
/5eXm9qj2MDy8fEHO5yeIYhLv8tL3r4uRFkJ0vnbTY2tpDNh4bJ+zJX4LFQc/7km
ktPiJC5aeSxEJKWqaelk8H0lcudGrmwic7sRnVfQbPVb10W71Pw2TdGJd4kqU3W7
1vcTVzOWv3Mq6BuJWOgRXW/lxIPb9nyhBx2nMI2qmdlBguDAddMkofjW8ZdCYwuB
ye2yMZjLNOG4twlVtQgTW4ExafIG4mOgll/QwjY51K7GNtioucW9qA+DAc4czr61
mgxYD03l0mdk+MDoDUB7GPpaa0UbVh5C1P/jMvuS1dGqFm5XnoKQKWewyaTcky77
yDP1wqb4q/YAoq8VXWNkJaPOStMBLxCAVyYzSVR8hi6zl2vGkRuyR67yF0fvlVN2
Ln3H77bF91NXBCk9M5Hz2U5OClr+Zj+Wz6JQa4WwFBkCmW0AqpLjvrGCJ2ptX5YR
0KkcYF9EERm1v1srTT24aLE8CzpFRr1f/WgfAI5bDuwvMt3fEovPXeMPwQ1hnZ95
uQ07tHpnk98Kx/IM8eP1Zd9AZl9FGLaxUkU7IBjP+CJ+qVgschwnSXfS5UaCzttz
QeI7EdyDK6q0mFLum9dBQwPsxL4cjcVtz/5PtjkpUTa47HWtVrGdVN8++roSG4gS
Of3OSKoGqUTAtCkFQHUcZ4+Z2g05Ds3R/fQ/T0vYKMXwYjz3Y36XYunihSRRoHP8
X+cppUpsoVlEW78RRGBvFGefnJc0ZH6QIeS7oVcihna9/c6HRT/462CeEU0JI2Q4
Z/mf64UsWX7qluANl+Kss2uzvwn1uoKEnjevqbgCHm3dLbeoEndF+MfRfnO2lmKx
Cgjp3/eFXpFUKGKmTsdqR5SHfnAYaAktYcoT7VJWqMzYoFQ9VX9ywGlGdSJRXrF/
GB2sRU222BwJBoKDpStdc0DBttStG3SjmfTZmXfMDMI42sIpXdSW+6ddTmCT1HCJ
aT4ACrGeHpl8vkWYZmvEOm8ZRGkNdkWiEiCN6zW9AT8EaS/A8noYZWKsV3ZIzYbk
zBKImqbSZQq5WWNMF20fFPWoB8RrJPP9xp4k4NV2TOpuxLronZoeVCERtH/2IM94
GAVp3Bu3WgTGU2/20SsSYioiieReZk9NnXlHgUVTKuwBdBii1QG+CMD9+QC9heeK
d0kqXTNTisjaOm6sql5Ws2PYNRfgrEPrbQDjoW5YdYXAYGUYfak2IdyfruriSG93
thvoq7VGBZsUqbf8Gdi5JarQpMkoSd+GVIlJ4h1kCL2nDiMJGnN7/IE9cor9pysM
ModwcPdrqBxk6lcF9nxbtCcpW0ps0be3uKPwyzak2fLpy6R+8tAjl+USjQ0hmb3p
Jz4GgMP04Gl5MEUYWupErZWb1l4ZTCJlHZ42mniQIy9MGBgD8YG/JOBmu6tAB+Av
NkNpvPJs93AFKivLsw8UZwP9vFoeaXVOm30L+m1NkYvp8WPlvxJmi4Rli9GR2Ioq
ZzECS8ZUI8uskzSzib6oMIo28TWSbrf06vMWf9PR5F6sXg0TjpanHnGn7og4fVwO
NFoch56EhQT7e2rD7oR9I9809SSxedUQQPEJD41GB+Xp1QVISJCCWr3vGYi6BxuU
s/2kuHUPj7NWgz4UMwKZ2Fjz3mq6Svwn0UA2GUtNrqG4K4glShMm6zq/Af5OPe0G
09csN2InEj0dDHkECWtx0nK0af+H9afY0rwKheXyEH+bzatoTYuw+ssLupFHdF/Q
K5CjSBFOA8REi9YV1etzbkIzbWyF3xA03SvYM0LoWuqrSgFN3Eexn9PgUAxDdaVX
E87aEm94mOwoa1i6EN5jrmtfQlt72quZhzuOmKX/+Tu8uk+uHc/Fn0rHpZo3s6/1
D+2alqpsQBPnfCW43fDApQADNRDv4Setp991HpPXVd58Nj4wKu+Sv/9wE3iCU29W
ZZVlspRjzxUCmNb2lQRAJNqZ6cbZmXdX5afRqJi1aR2PghqoVMbR1Ouozwa2tK4+
AEZ/tIfzjy03s0iRWoH2sX29tdwiKtaQudWzzpCZu70Jo5vFUqMHae0AODmatxp/
asUBx4pZ/swYoW+tauaxYSf4guAdNK2ELkC4DM6z7s5j9l14k6jpmoxjKIJ5+x5t
fT8PcowKFBYkDY5YJmUmOH5Q68m3Nkor3CsjYMOZ5S1KDtmwO+8U09mmXCSUFD5E
5V51Ik4ssRc6P3i9Zhzed2hbcBz9Q+qgCuBjT4ZgRXNJM6eVEEW0mi0Z4ygf5bp/
yXV1VrL+9zpVAQtLmnPo0eSKgC4P0XGVqjv/iS4CbUlAGamv6IzKajL5KQLRb/87
bO+l/nx0RKiTRSM7V9iMdmXR0dl/ZVZLxs1tjxRlAe025meoda91K/2cGkp7AKV8
2d2Ln2S6WTNXrBuRDuREGlEYhMPF06ORGdEAJIK2/Fe9KMmUWM/uMO15Tcm/z57u
36oYnNQTkhOgJ9q2UuL4nXFYk2OGSXljkoG3oFiFjdxQldUGJu5BAR5boUtliiOA
iwX7NnmvWb8y+LJqOZ8L4gq0n2rmthH5vCooRYv/b4JC4jy776PI9aCw7mRJ89mC
/xDaWO5NxYIGmORNAu6DANLuIOT9UfkO27h6jZ1RAHqu3sv/0AXMUeGSRgWJux8b
6sn/xGechaVStQVVmKCLTKfCn73XZG6RpykBgbzRrRVBwhAK9FcjNcwnhpe+C15M
LKBJgmNuFV2IHDY1wfpwtZSk1h5Z7JRNIyiuztg9khiwV5AU1lh8VYHC7+FjaPvb
GFKr+/p13KPxiAfJeQDnDZ7MH8SRsKS6+ju0H9qYEEhie1WlIhD55XfXvjv61EPR
/QsLMiVWy32kjgI1fKntIx8qYO297KO09kZQq+0l6eIHyqjX8iWHLKlhOUOZYF+e
EMfPd1ScFLtp3vvqMA3BhhWHBxcUiFniFP9irrobufWa4KP8SDy+3I8BG6feTGC8
W3N1ot4dtQDdV76WqVjdWhReoeTZd40ka6xYkSFHirvqq4U5EJp9SYwA3GX52/XW
2nKoUUBi8KgO95hREPonuJeTB2wBCMcRsU4/bqHeGsSQuey8ltxCBYKT67BOnQ6x
nfjNou3PgKX0XCtDfode2RdtyceRecKe9vpSC4bZvBCPg2RtykeJhv6w+qRincG/
OVHQRtb+PRZpkb2Rmy03KU6UsoW8zktt9Kv5S+IwgDmRUw76RXiIcCy2Rno+/HUK
AnqqdNFZrTvNlq6pz92UcEIFxSJ6Xw33z1KUJ+WuaQPdPbaACuGIheMixCiOKiDG
vFsvfEQ5hVIcmwzxjl3XRHzjXYItvGNULXX7/uqeOD81x0Ycuu2g+TzXF9byDVue
FOx7DonCBjfhuOfH5GLa/d6EqDQe3P+CqdfklynaL5oLVzqlSoAZMOLmCqhmz58M
mCfg6NN/Ra8ldIeUsB+2hTCRHqDO3sEGrHlZnMos4QlIsUBalVRHe8Xry8ZpAsoH
b300a0W7GX3g/Er8yJOJc0L7G+GU2K/hpijZuXEJ/dJwAWgqcmWLT81uEvPeiBn7
wVQDmKHoa0YVkQq1iUd+85JjIUWEN+DeHf4imJIKhpwCwxFQDsQv/lvAO1jiZauy
uFXTgBUnrSQrBzgi+dKNginvfcuoGQora7oojwYbWadZQX4OD8ybUFc2JgcP926O
Rge9jyGxpX7zkAigU3u/t5qyUVNI9var50AQQRHEVmpXL1up4xK+LwF2CZBheiRN
i8EYV35Vf0UQDdgtHgTgVt5DwNLnAE765dMxK1e6ckjwIEE6XP45q7Jtd6K8/ofw
HSoVcgJQ5oSPFDkFByA8VuxOIHuATIqLZXJllJVEDeCkt3NvtajC86RaBhxSJS3l
QNrySildR4zeRoNEFGvFLhXLM0Kvuf2xDwiBnmukyhKZQhmfoVapon9JsddSk+dQ
IwHykjV85/REl0wD+UrUOWUNAbhql3XuZqWKVsHuDAtCqbne8fa2u7FeIkqGDB5h
v/bMgFP52Zb/3JZVL+RexPAjd2WhCQDrThuBJyWyDCjAAgKVlKC3l+QLF/Iqy0bY
d0M9qzgwTCngJe0UEkc8nd0qj3ZQqzqmxfNWt8dAArPH3g/DIoMupJd9WadevGw3
Wrle8bQ6qVqijOCaVcxsp65MuvWUUDNSsC1FMYTyv4PkPa75xupGvu6uqDOmFRUB
b2gPiVS5/4MIhMZ7UGOMsCKMsKzqybJMEvaMHxtmYJA/ueIBrP6mS63wJ7Uzum40
N+9T9O763yr5mc/p3gqtnIXEJdsD2wDUqj/Qvjw6o/OD2eAIVXlvSZJiZ7CwYeRv
Zke6bSXVzJGxy2Eg4oNk52zquVgLybSK+BPnr0HmO/Udwztwcph2NIYh6dXSk1rm
2x94u5v9PUVBdJCNWztPyXzTSLYczPDQD9rs+HX7xgX6FrZL5j0BLqIO+wqFeemJ
0RPfBguLq1UndE40Y3HyFCd8gLOJj1k4+Vhc8KG/k3Xgm7SYWXRGhdDhvQ2ulXvd
+fogtXf5noFLCNhThTZnJzxkobTtlhp72PTqdgC0nC2Qli0+SJbrsAMeWSJJgw1I
viqam3s3TY3FDaoX8cR5E/afLlSZZn+xzolPt3RQFfv8vL7AMDuRblTSzvIhVatQ
QDvH6mtM9OTJiItaVQyjqEuQew5jM4zUckYYYlFVB463e2KnMBYw5igPGjF1Pavk
up3IOxNlLEsasYxefgg6CGAOvaYqGrya7hx/iMm4JYuZX7+Oqt9qwJlpV804OeW8
/LXxDBsPJ+mr39+Tt6T1QAqH9+EgNWoScCwaa2uohp6PQMcS7TABwRu9BlDoB46b
iGTXVZB0ZkKPgJsqwn4XCth1tDtcXfanUD2idc7ZZdnPf0dFUbn2IeJLo79TIkYU
Sxbkc8HW9TmCxFFh+/V/QTecAW9ofJCDhKXXnQErmlnDQn21x9YWWmpjFoBx/zIS
PjKk4qPJLfgqhpetg/LvKfCMiznHcA2m7eJ1x/5hGR49t8NzMiEdV4rUTWuI4FMP
7lUQ0rYIVxoVP7S5ovI5iOVnQaxC3A/qGbCDdX+nSLYKRifEpLz+sP9vqczDWBT1
fP0U7TyTFb7tAyJRgT/G1Q1c9MhbqGx6LE4aeT12KrLgdkxAemBuoB7SSKl+Tdmt
i/i8SuQWo9KZRID5pkyie2reoTh83H7AHlkXThUIcJvKC6t8rAM8vVfj5g9QuENe
ZjuOri7C2NV9rUwBNCUlf4J1dxCnAIVOokjAzXfWCm89TT4sUXWNMZoOlLQpIOqX
6UJwFVvOvE2aEtKaQjoNkAnRlboWtPARLaQo+YpMemJKi4CQPwXpERIB8pc6qldq
7Hx+DFBhVMy3fLtYsjfmV9txxetkae0ZARfTp4GhD3LB0PFKNN/uFN4vPR4w9RqA
RWivo/eAlKU7t4IYODIK1lt4WHeuoUc56cOCl4l7pWhSUXSxusrIG8WknDgRcLB6
MX7S25adZxQHDfuU2Pvsjs/6osqvVQ9K6+rAAQvOoWqkZqjligHHruGeX4iy/c1F
VxWJfDUBY8QoUoPlcXYTixSh0RrO2gbcDS8RaqTOKRLUux09K42k8HH5UY5veU2T
x8p/jmHYZxkm79mroWbtSU8PS9YbLsgBA/RY1XrMV16vJrBv4ZvRKNMVqyCsQfUy
za5r7Q6ATKcpr4vcMnUp2q2uIV3EsKQlJxw9CQKm/bk3d+HPZZWbNXLhNbIJe7S1
9w1ot/MEFZ6J8vYF4JC9/FgYEy28l99r2C2SnnQn8c+bq9HTMcjkOjrboGuOHr1i
pACV7C1++/Ey/rO+Jv63nuOeJ8llZudOH8OLleEXC/DlX/IlNKNn9xX6GCPMBgpA
8AMzhDDK/X3zmQSu+gcgpl9Wj1owwJ0Bfc9AO6X3Uo+0O1UrKRqrqFybZFmPN3sp
DTVjC3kSNq/bpw4UrGm3HGCFQY9bfIPW47dCdbMXhYf1qfhJfI2BBMEi6BgPzXBy
m+A7W/xFeJZIKaxUfvmeLWtp5y5kPLu6LB2rDz+WOpBqHJ5EMl8W5r4/I5GYMz9T
QEKl6lbiNURa/J1wFv3OvSYrPkuP1nx7B+iNdxOxA8h3YmPFytapNAXO6AfBl2ct
t+Z2ngGRbvOvJHp0jVQKc2GohPneBAnXTXBrIcreJO6r/ZsDbkfazQmZLPk1AXLx
NBqAFyPT+T/RULYUmPLjLSoYxuQECHEi7M5WFywroSf5wUPgPmyBVR/c++/d4ajY
PsNFw4L0LfbcdPDXuaHyFU9pw+/OwXMqjoi9Rqm795LYPcaXCHsPMqYLcMmTv5gE
148qEpsTYy59xouSpi+X9SSsKFfgYHe/1kDeCASY8B0WoTs8+zoY5FqFHelcp7Ye
7CdRRYXpoEL810oq6y7oI4Gkiymh27VQW1GgbUUwvhD2EJKuF3av8ojbOQrqT7S9
lAjpUlMPp2L+6MG8DOTAOOtr1kaIgnivB/TvFqRjspWEmdrxB/lu3v1qKC6oCV4R
AC0tQ2p2ZidoScj4yZIAtvRzSkCjcrfYOKzaKmI3IP9m8P3xdRnT7L3X7w9fYHGE
5MMbwzpBDNub/lMK7u+rXFZXA4REdhan5QIvT3O9z7ZD1A1+pyDONONOgWtvVkvU
Hu2pt21moujdqJ1MQMGul7gsJyyQBRMYCOwuFoc7GsiRTJXfU/PqfeSj4Sk02kBY
ImsJeUQmP42BElZtsN4T08F9Q9vwlQmxX8gaHhS22UTG5PN9/cJPoWmElLYHk1p/
lyeIKrJVEQIKfR+Y3q1RMY2rjpZiB+zLJBpAHYeiSBVY1cEKRzCVVxnup/a00hls
iqeuDdGg1cBYGeXhfm/kx3tc3AcQysA4lqIMnP3UtaFSkL1GwyEK7VCLNu6/5COb
lf+UXFr5VZp8x2jUPlkQoPHn8kKmO5FBOVjIGtuwXeGHGdsoEQtUiPZ44Sx57JUk
O61LJnVqptn4KxcsImsyHG9F+DQ8pntRllXqxKHMODfsNbFpKuV9AQ5JCPn51uX6
ixx6kOAozAFA1kHU/0N8jKLlMm/IzaUmXhMMTtGcfQAzT1aILFM6pLCPjXS6towV
gMkqSajGjrQ9Gqt5qgv4EPTEFJXxr6NrU0xqaEvwFbI+uxnx+4Rswn+VfXBtmYgA
0Nj12W1C/XCllOIqIzmziPP3cXyrDzyjZPUYbnTtk5sD/PnncCORyYFjCRzftSfO
+nw6r9VeMP7q/F42ATAZwWZsGiCeG/38h9PbnF5E1DX0UNQTrouu5ggykL+2Jb9/
iZPnif0ybXGJ5+0qCCB0UpW3cVkRRfcBNkrI0H4MnzPAUC6UsEHm9TMwBhRiLxjb
qoIUXRALias6N5CngKw0ZFyZHrTtDCJfmg+eI/swGazcDU3PgX1ixiD6qAZN5Axg
fTqeg6ex8QZrThEKo2MjtL5p1/2ER1LE8XXR0hWuKF+YSr2MlwqzfN7S7SZj25hr
r5I1BNROmQ61uU8NoNjS9NhOob44ZJ3agc3SP6JJFI5bqF4W+KRXh1M72XaTYjyl
ACb8Mi36NL0ZSA36aiNeJyEElZpb0I/sIqAnhDwE8NU065djaIuEuE74UIMsfdfm
+WlUHdjNsiGRNB1EvnnK41D/Dfa3vz069fy+wgXmrtM3PYbnUVhGbFxZVBCljsTF
KI6JuwoMGOZOW5N2jxTUAWFzmshHstUbjDkhuNshUXUh09naxw+eE3nJqRDm7+Pb
zwAb8E5VQvyXDMMFZfzsbUI1UPwZKU+EXR0k+hRYp26gJd5no+uNczvuqWVTSEPJ
QpoNdS2Dpw1hPVBvLHEoNS6nQlLdmCaP4W504nmK/jnFDbpyYT7BFp5pyWjX41qj
SHFcP61a44K9b+HEJqoBAYm7aMA619N6YfLO69Mp2PLd6CSSHAtQaUg7JPTulSec
lPolSzKjWoRvSi1LQkASLCDuhCBa7FqIzTvu3eQtxy1PVXOsFjugHT8NtzKn0nsw
RxoHGzIxQHsDsvpJRMZz0qWBiCIajR8rqSTgbo8cPlpgyGJVfGz2Usezv2JjDlcQ
L1ZdI+AvJl+2MxcD8XVK7/IC4cX0p4/fBeRH+0WRWDC9O95GXJ+KVQFEYwkXrP5/
M8rr2JvmApdfYakmrVeHxLEcgaQM36LkMXu6nNj+FAhFoI7hE+QVuWWbpBtg+cD+
zqnc3IlQvhp1aX05fJj/f+G8ARLSsy3KEaWvnSlndxa8xV1UHPUyydgHhRPLeSkq
JTuWDbZ7Dwb73h8wkfdq1H5JAa4strnHACDwykkaKL4fQxvsXZqD85a76mJ4TUkE
Cct5/DNunPhCgVASB/NrrK6XOxqKdjwJPvwJkGBwNiKUKWqKRef244fk3eEnXOui
/gXnRAMiZf5QYjsMu30DwwgQG0ZuzPXfdja+gn6Dt8LogDWqQttcm576Iva18G7P
+OIfCS0N5BGDSHXcEtXPqOHPM1iNNZzWTf8yZOcmUCdBleQVZO/hRg8rOic2HvdS
dEha47jtk6Za8P7IDm5bufr3VCYJFabh3a4gyVE9A8YToWA4oKDbYG3iAaWVXvl6
d/vuitTM/O8UDOEk/SKjMRCu+wR4x3ojuUkFHJfU1Jn0XmkBBbXqG8yC32lCjJOJ
oiNQDuZ3iCvb02TbKfitLPuggqNrk1mRRc9do6ad1aoC2jiouhfP5/p1Ftycqzr4
2rIpsoAD3cxDgJtsdeDhZWzYx3dXsb5cim7D84yRhjEeyIwpZHpXOkVKsxw1zivS
n6hFZtoZkcj5BsXYe33Z9BeDiQUUgd19Cwgrlz00wAZtUxjNifRjHmbyFKW4J5OA
7lwHzyMjvMJEMDxgPl46COiwQlzrl8TpFVdK3Dvyjqpp2b6Di9arkC3x08RR+AX7
VXAV2lOjkqHJIcJX2Q+9q0ZOzTlTRi6yLQzHbiHmwi4SJjZJ2qPtwTezN7GJZizZ
iN9KswNYw/XQ+fkW6KxPzI5NmAmpXu/yesViWGeZ7zuZc6yv8Bp+QXybKKvRxdNl
hveyJx8V+aMAwjFgoOGoGtr1SpriZrhM6DM1H2Bj3JbQnb1AW589vll8kpJ4Dczd
WJZFq0YCZ9JbLU4vbq3LocvZConki8+xUJe9KHvCCv28359jdqkITT0LGYIRlC8A
Q+mzXUm0in8lPoeRK8hdNoVcRlBxS/dVnNDwimMv8fnvZQJ1sNeCAYemdRCR2me5
7r9NDmoaQKKU3cFbFXshSg04jXX0qEazw9ZgoDrfP/Eh3sPgLB+Kjj9IK3ImJPVe
0UwNafGyIyEQkg3HNOuEqQH12VHUHvv7XtUe3f5c4xQT6OhoF2m4hTiaarqAZIG2
P4uu5TnEDGJZE8QnPtNMn19/3jtl/TFBSgCnsjnPEkn7XZtkIKDZ5xS4CIbPWhx9
xqN7nwfyl3HX7Jrg9kqf1559XpAd75B6LcpQfFNbUu+tX+MAERZdBg3I9swAfrbM
dL4lPD/KOKQm+Guf1UkIBqyiCMvT9GaoisIhBA+LYnAj0nN5PFcZKRRVjkjEsZgo
iKt4OqXHwmGkgAgx3W91r5rV5bNenj1fxBM9l5NCD/0M6oLbHV5vznFGp9KYCXt6
NPIAwirH6zva9FoYNNh4J53euGzMl+pC6rx9sAGaONko2aiT4E4nyN1Qp9+yXrvi
TLlwWOHvliQBUIgPovF+Q3JTAyD5qsVEtaZZh7kPzi2W1fXfBG9bs7Wt4AzP4Xz4
VEQHKam6vXdo799mXiBXGZ+2oZ3hpzc0D25qGcIKRH+bGlG/vnnOQl8s8K1zD/1S
rdIlwE3BrNm8bLkwSZn+4KNLecOtCg8LLqdXUPn6huBgxlkeZBfSN/W8xyq+586l
+Ifg5lJG0oQ7/HVa9/WgoRMzgML7sRDnm7zen9PN1JWd3Ldome88o7Mzwexw4+Ho
a4GDKroJn3p0Dhyv20NSWPRbbjuNR8PW0IqluQaHnyFqp1Nt/UxByIndAUglBb/c
nNJiEg6xojk6wMz+LThveG9ebVilKuQ79shZhkL1BzowEn2ub3ctQ3wc/gTd+yag
YG5kZNJ2nisbtbfpyKCaZYORh9j/cWQejmUM3PlJfHlWdSIqpWUxFFapUoIGWYEQ
5OlOMPX2aacUAwKGa3XgzEuzXSNnYuvwuLc4uBqlx+jyNRv14v+iX7owThMzzOGd
gyZfuTDbPDgMi3g/8NgpmOFSQ/W9WmHkRXtx76sbZuLU/1KUCWuqptK/e/KGATRw
E48BrbwQhY+QZtvfuwxcJiKfjgALhYBM3QMoDWgahs1IEBQe/VC1rHUL+1xG9ymV
nK5XepuoyiJpUlguC2s7xWd2Ykil7QlmiBZWNDtkd/r8eApxNWLiSUYlJR6/KwDH
SfVjv+kTXXWRWIur2APGFK799ry4FQUuy1/k7+mWCLj11JkB4x4M5vKb/zRuaKAL
Xzh2vgOCichQzXbG66hunMvUktaqNX7+OIdppX0fCQgATSnJHRa3yUMt+owT8L8/
MPM9JqHKS8DRk1SEMEjEgM4HDEv/KT3SJcEdEm+vJ0Z0AW3CTB5ReSerLDaZwrkD
KUTjkDxXdU27ynCgQOP3wp6ORrHUBMWNriutDlc/fALiiyVcAjzuxxPRoiRQB0uz
TPLiT4sKAOeWo1loWBr3wBZBS3kzZ0r4dxan21ZsDuMUlRchhE20FtY9Yc80t3o3
ljy33wCB4OXUIJtTltaAualRX9qyoiToO903MY9RRswdGKBMdXD/6ST6EpdWpQCc
Jg8T9YNVDZx6v1WnLANsFdFZSm45Q0ZXAKYspEEQJNUv42AtO6IioVUxh0I/KrEo
h85NSWsxeDM0dTW24+8eVvx2YSGvAmVWdM/PYlmIo2QRzsry05Gc/Gr8qIUHQAUn
iA253Eksl0Auu1d3r6eT8mIwzYgRn/BjgU2kLZg9iodB/fFe794/xQk/7eN5fyn3
nan4LIbM3bvU+Nh5bcYs6uab+xNmvkaWsOBrYiPALfq9vzok7GLobTD1PnE6OaT1
LATY5sMNAgJGWpf2gk7+EHBKfpsD0J8ag7IRltj+QigdW40nRq0YUomel+tvzhtT
ej8UDrIJv2WYyaujz+4Zgfu1jO8MJJxIzB6RNIgxK5ZGwQ0iftP27sE6Pjuck1Go
VUkfzdRKjRpvuLluGhwEbW9TgAjvRW7FiYSiakf0aMMxqQ7xvnQIWjHluwW7b3Ee
X7D6Or+A2s+7inAHFrWGLWat+Uf/fefouwlpBCGfvHjuuy94yC3TOiI+yPSq+OI/
+Ox+tcNJjH0Zt4YlwAZRYVvdCRkObYWPaFsFeQKttLK3Ap8BKqoRyD8RVAPeWIHm
nKcCogx+f8bzEuEsoqjPn3UAuWpM1D+4vFYPqN6sNGDCFxk/PRo45zecnZIy+uoJ
4ut8om1nFpfL/dkF8CsRlzSkV1qqEuXIxM2SSkx+rGkQGN4a+GiMcmNJ9xP/FFLM
fKrX0nX9gUepTPgKYiWUJXBCWqQG5d73yck6OncM6Fiiqdgj7Ir6SGmdCOAaGxyC
qW+ROU748on5o3PfhP1MU9RqyfZUvXzM3KWhTy/o+VTv88fMf3beqoNHd/WplxVw
j8IWBfl+g7T07h+dg5RejwD7vhp1cL283QTWUcqSvTfTtSpFygHAqSDv8+ILhaGT
tjW6fX38wZwQQsmv6jpGIqw/aYnb9bdT8kdDDHyzARnH6nOAwM2EtVawr+xAF4XZ
Ld2Hs5i/K4wOiHjoy5Pg03N5CBmNc76QhPTFjMcOaYIY7dsHjcn6onxKmT42ibtj
F3TFp/8ypSCWLVAB9D+ncbMjCIXs4AVRWDPcXGcAQN9c3p4q14hdQm7chjuNrhwX
i2ambx5xQ9BxGB8PoflrmUyznNJQsNmF+7GC8RUdZ8TWZmeafG7CcysXywb25YSh
vU4wKFQHGRw8I8BUdCxP+CbAAq7oXFXYgYBwqADVrWpsrIiDbdo2VxubzyrL8qZu
io41DjtELaoAeQiMmQyF2L5HoSKPaA9MyOfr23t7YfZrz18RfvUcsUBbG49c5514
JtemKyMT8xHj3uwRpTzel3hP1xaqZz9cx0d206V2efYeaeua5MY89fNHsE5bYidJ
Anm7yTW63Jwx+440oKyDx4CGS3Cb7uWQ4j5FHF8qVHOiWnZ2w03GeGHhTBR/PBOI
INweRC3zrpt0OM7HLjG7wYWzL4/OdBoTskYeD5y6iVUl5teik+IZ1TPELm3rnfcS
A/Hae3Ddug2AE3RAQRc7JkhzDw7hQMvOug5052rYWB5AJzjVYK8FmQvPOKnvzmZK
H6zqh7jj2G2lHcou4wNKRDtJUfiMTHr7PJ7yirH5LlMLd9Sgc2WI2vU8tWowed2j
l62aLFYeQkflhoF5j6pi0MK3YUE2XlSQtxO3G5OamIHutGKIbVfmlgzCVAXWd6h3
R8VLkrqcUahDOJTjQaBNEz5VCa5lRRn+VsYMfg8f+LKkUPect47UYhEwgF1ldPO1
IxRUvINm3AXKCF2RGa6mmfI2beR/f+zkS5HcehIgoHE76qohMqpT6eweRcV5xhrl
IFBvvywrK9+K44NKdJWW4Q/NXcponJdxo2sxwg0VD+wDx2AQ7IwuINrBjs2xcLlw
p1uc/Hfda6ZgqtqNfpisaUBFJ1Xlu+C4SUSkFEsVozx7N6VCVD2k9oCakWDk4/LP
9QsH5mXQLON6hq8lyrQtcJRE9pF8EvA8M8IOeSXhVDnLJ02MY+GXhrMezAx/Verq
+Di7btVD76t1sp/ZB2XUrtYwN/C99+STlYrpgzT1+TJzPKC3T7ZoZ6bZFe0Q7e7s
H7+L2/6vJboaGDJnIjRddbodWDhqS00jjtij1M+fQaW+H/81ILt/jQfMEzplQmRT
S6nLpjAWkLBUiSuArTJZvK2FhWF/lp/RY/gzJ7MbWN/6gqJZnVaPI2LrzWcSprQT
gX7WytxrZt68CdZM9H7VNXKtLbBr8UTC0KlmVeJKZTwrqOwoHyzKH6yasJslGsv5
PkIkJgbJO5ZArHWpyTRCiS9jF/uoWW/f9t1z6rCXhcHYxScbINdUWdw1MW1M6RBu
bLHHb9gJJg/3qbZIdvAB/J1xdDEaUPeJjPAgBaZBGbtSLGTygg5dz4GYmXeyuB+s
9JfitI9UzDmA7SCqnJQT9NMi5xf8PNm6taUWfqyAP+39qRwaUndaLNIrJ90NitJ/
0sxzwzbBghcVU/DVqObXHAWXDWaK7EKMT4pf8JMAqZBAHlcoO2KavI0bfPXIy2AU
opwg52AbDQqcTXzGLFj933QvTKx9uESJDV1XOnHmyzbrHtMMmqrriaVk6TJx0hxZ
J+o1iYwi0/fOvEJ2Wynx6PzHO9cVjbiO6mrNDKcAPF71BxoW0rOgkA63xmqXBf3h
L1ua1jHHBijjBbWRYm3XXIQ7e9x3pblD1/7lLPMOMLWRabcmtS+zCRzJjCcpSd1V
rz4ZtbpsnhTd9DmX/zmuM1tPtM3qPSB9wsBMyHBD9mtawTXi8rDczvySGsLj2LVJ
+79LOJsUTFYcbKsz8HkgRJtWm4hi7e0f6Xlz17aZAMqsT9XM0GWw1JT2zFhRKq5W
WExuhatNQLPbtI2YS0kvt7qAAm8Vb2Hdgn4iL5KHJgXrInIKmr2TxUd6P2pdwt12
zY/s3hDYi7QCL/LW3D3YGfaWFEJtvUYtD1J50+h0TBUl0ZqiicEhyk6swlLztZWv
HbZIUkcZI6zTOW1XK9PPh7mg3uiNk+IAuo+FjpbWN6VcDFi8zah8uzXO033xJHAi
o3B5UtRSQ6xj29V3Ab9UzdoYcxG7E6XIxeoi/H1dMN800bO68lGC7M+mNWqYYCmi
Hpjo8Tk7gzlbzhIr/g0FvhUsFOkJ+p236EKvh4TOoMB/FykDmJKUCekXV+5wC2Iw
s+5ckICJgKrti2G85WUoLkhVdSxtLwELcpXx8ERr5t+CKqjkwn38gCe9DU9hdBdU
3MQ1/FZ65jOH2n2zO2o8YXmlBC2rgcpm7iJCsH1RmJXMpZXYHq0kUsVaWC039n5y
HtozZOP/oLjE3qx3kaow3KVAnJW4krzGHWHr4O8U7V7/sfryl/fsCf3G0gAMpUww
FaDZgGCi+mtgo737ktd5QKZJPUFDqcJP7K2Z457rL6NpiOMXpX0q8rH4Iz8GNNV0
TDPUfLjB6GZrhFkdGIY2u33uz7dILGeW6JaWykW2qz6OVE57QflvBmgdb1ma0axw
h4ASNLWp/GQPwDxV1Dr48pPQJ1jbR8zv16NXgnxsVE/jLU3yIlhUjzA/UE3CogAC
puJ9SBzpsXkM2mTleTRdDPRtfD4Vfd6kBFBLdslgVOq6e7yclpUVxfbW0AsBMkth
ttH1FHZogZRFuAHsyleYenARnQzN6v2NpjFaJKr7S47egw1pacPSxH0i8S42Ceog
Vz/zYfADAmMI3upeRVCumRjVGKG5BTCNFo4Xq33MWayac5oo1/c3DKmtGk79Oem4
7FABxLTn2PXN3MQWsl5FtsRplFTltT7tNoe8QOm5/k/e5IwCsAIe36vP+1aF38QV
4LHJzcVdkPrdFkupbnGw0eMHuuiHU+NZfxC0Fxls8XuhGM3Wtc1r3hzIQBMoJNye
OVeOVfLq4/41ZhKhx//crnvjvtfW8K9x0whdm8ak6fu0zTIEraRokOCDmWhCe4VA
h4B5qJLmGS2EBcqG9ZcK3mdCoOKsKoJvEVHE5dNg7ywdVp/7A2LqwG5330BTijdA
M3mBYcXBanifa+emZRtTA6BwIuZEh76tGwp7aQT4Yx7nyUrUp7hYeyU1gYFs2Fku
4Bb4zdtbWpGv8KU6VtAs48X4bkt2Jn4Z5ZYm6xuQWYaADz3wisUeGjuyAhr1aejm
PwtvwtQoOkt6mzS0WylqHhd4Mf10mcTtpuNjux9TRbggsRh2JLx0CMyR6rf+/Acb
qf/faJHhjOBcsr+pONScSsOAfHOZh6vS4WFIMLz7m38h27yPF6+cYwH0lglNhUWG
+J0i2B2iJdWNOKXw4Swl6QetGibUkmRvPK5DYq3zw90dq1wxEVo014RbsdtjQaGb
k4BWce9/28w7Qnd+k0sjkPd1ZUZMT1ppYLW4DlVW0uFa88dEt6HPtjdjcObrqNR2
sLQJ2nFCrUundQMS+XlqgkuwIkgTFnqtOUiIJtiTX19DqmXnoQbVIaqpEE3hcOJU
Kn81D/PUylNeEEgBEaY/kCVx8haLpKyG8t4DZIPKT3RJig9GTS5Oywvl57dLMTxp
2pZULvnc53ZKP9s/CngYcYIPI/03TC0ga95tmrcKIIKltUxJV+/ihmAhIZN2Qnv0
DbvKa/SLS5rVTLTTB9RYQ/u5LmpcPDM1jc91eLJq4sFZrKzi0MK79xyp4OaRRI0a
KJAOlL1QCNrPqnkfOAQeWEHrVv7OmUGiTW6XHsJ/0z8PPlwFe0mX5OBaxLFNvSvi
2vt/luNxOTkmsItfZ/fERccVILXAqdnj1s9s7k5ra1EE5JE3SDr+WkXvUklu2eYB
Ct/T3+xKIjNQGgbl5n4ZV64nVLlHfIrrvFPh52HzYphhvTMx06l5fSquDYuQwryZ
lk8oBYEs9UfLFlQ3NUZ6g21rpgAplUnYXPMzqNPdM6tNS5XdSV9PjVs88hY9Qt8u
ym4DmglRM7DPLJo058bjNKUquYhsf/DDJtYq6HG3TMyLhXbWbf+h0YDE70s8rVOu
/hSx2p3sR4z0pDv6bQLVgdHdBzoOqj3wTP+e/0wUM5iJLRSO/1/L6crKBXpUUC50
8hmEMx/+7NW0pywdhK4ol51q+S6pxodny8c4WoTSJ21wfyRckUuiIuYPV/Qui4qt
MAtEfZgqYGi8fIE6l/a0L4olWXcHx6MqnQW25enITj5TvNwKGJqCoDSR8FuQR63q
kuC/wojL73kGGQujnQrzfnxEm0cIB8ewmESmyvecjG8foxU6YEkkV9HM21FImM+9
Eo2jQEU2n0dYE+VTcuGNopcXqiNb+tmLesG3xYJi9taaIIbfDiUP2qu5hzu71l/L
+97+4yk2oeVMROfPXokHVnt3RktCidmla9zq76Fnfs8G8zHougGNXLFGirwQooo/
FIpic+J4raOqVobaUe9dKEaeiII2CN9pJyjZDHI6Z7/KzTE99I2WZvtF1aRihEaG
vc5QI57M+7cvanYBy5pf0pFop4Fy/II7wxVDwhHnCtlSmJeqpQVjejPlqT1dr3Nf
0F1XBIL57tGZE91LULlC9p+AXyAvsoGQHv5esuPW/ib9+FlnvyhpVGwHQDXwyq2F
6IvvBu7jhXY4ed+j5mr8XIzdVXAhheOskuChAnwlAS2ZpW66nwblJ3UCZ1U3W7ny
wOwkr40Ib+Iory5gcdpE94JYv5bl4GwLZkpCL4ZwoPDgTvwb5K+XIiXtPlQqLu6k
2J5xZafg9GlLFDtax1dwbLncai8wbC3DnHyKRF4f9T9u2J5U0vz89QErlmud9aAZ
n2OgkGkYBPqPGgv19mROBQJuIOo9CKHIriplW+GewgJWSuXW5zaF4tulDD1UtmCe
ROiD4SDAsrvFuIZGsYcLKEI0wiIX3wv5tVVXAJ8oC1NBAROAyNHl5yZTYBrwKDdH
5cZxXU3CcFtcFLv69uZWncVEW8AQBmnsFnEA7+SL/sQjMXoOD9t3HoufN9Lz+sbx
bwxHx1cRN7tLvh0XTBldz93f2t8oeaFnMgQeZpOF9ow8lhX9PQYNvhFZLAChOu6S
CsXVpmMO9xOlAEvVuxndp0eCwrgDgChRoCmfRupTsSTUWaXTbOn5OIECFftSIMjZ
/faGmtxpwU1CIv42T1LQDCwi1iI8y8HWeBT1X3K1nu+jcih4gj52HazUzm0KOrgh
ywqA/e0sUc+u121hYLWSmLLtyDKWKhQ8VWgHSGhuK2ZBcGz5vf8xpq05sxrFDdwO
cc5bh2Ii6cBRFSde/Q41WYbvc9uFart49Q83CgdJHoKL9fOuEp6rASPEVymCm0Qb
hqJmJ7hKyeAHS1mZeEfpFQSezJPXFIQjOqzLcfx8ebPoeqiFsTjhbLLyCAS6vlqp
IZ92/XCcrOWT/bOjRgna/zbgiwYWByo+Jbq4ZidFZZ2t5VF7dmJ9gIwr8+fPuw/8
jiLyefRSZZo7oNMtAqT6h+1JKTpP9z4SVb5ThIcSXs0EVg5K7+yFGga4/3RCuZRd
xfdW7KQJu2jy3NFLuBti9XQuSeN18A57my2AjwgMK2xz8H9aEIAdbX+Yf30InBAE
r5C0TWQMu/pUT5TAPE/0GMqr5iQsAokWgtiQdtyKMWz511ZwzeerYqFj618mpQMF
z/JS4Br3sbUuzgot1GjbzwYGeAaS9jbnbAn5iBKuBZbcGwOgrSQz9+2OsJHrOKjF
MzGdvz2h1hUFU+briQXPWbuyOicllhACHOt6/Z6C3e65R1B3rJkWs6BYe2/CwpV9
RJMlA62i18WMJ1jpNWlnrKR55BRAToP5Bk6Fj6JWDDyrTqm2tzcMHViKJyj4La4x
sWxbLNXr2Lee+ZlGld+ptD3A5zXFT6jUxMPmsK6sNFyrQrw5lr+nqzjhboJNQwCw
TqZAsVsXSx6jCAziyPjTR4wyjpjll6qftH1gqoVhDZ7n+6foRO7sVgN0xqDdSXyi
VKGAdVnDKZ7zANYRtbLE94FyQ2TpnIs9cqWaua2r35S7sICjoFRNMvYAuWsphVQW
9c4egnJ6p5aLqjF6D6uruzmFHqo9LU0zm+TFb0HcMm4nmM2RB2EeykTvOAU48KDP
6RQv1BAr4DUY6VtEVoqmnrjkw9xsCdX+xp++g/ZvSAEQ4jbhZ2KupbTzDlshmc8O
RRL01XGt7qBZeladFxHHkjt0LzslxKKzAtiJmMrWisjzxuzOkTapZquC1SUqed5u
XFmO4aYPC/E01bx1TyBALcgKMkK194bZyurQ/gpxphzXnxCin6AKkl781/jlog5D
1ZhfnQhLE1vJUsLcixbxYSaqs1rGEhpWRoxVirVZgsI+LtfIom/Od0+Bt7aGJmeJ
t3VMo9lX1fZ5pJ5+BktBZIxC1qyeYVOQZdfrZHSFmBqONO1fEieEMN+gvobSKnrp
uDrwJmPO9DD7JEPlY20jUyr4brfivhpTejpWeAJz8nlXM6NgpaTriEKtyQD+XXNL
W2LcmRPYSG9xVLneJOJvXDrtg4H6QS0H42DAmuVp7GHaqUoPurDWIn3VYYoelBFN
rUFSU5GDxzQMfyCYZuTiy/5459nfgv2B3zKmRuBKKEa8Zfl0eS7n+7UeFwRvz6nm
iTfJ//XsMyYp52xIfsBIGlK0tLhp40OLRZAnjY+qg0TX2OX50sa0Id7y+SKnpS2S
jvNhJ41dfXPf6YrO/6AfHenpAhab6zwu/YOFjwAG1HyY27Mt+R1YdBBvj+issxoy
QGGDi0jjygmBRRFxePnbxVQNSUq6EFr5RkKwBw/XPVHUEjk2lsLztoQpA22pFwr1
2uqHhWymUyAKjW6OLjru5FfMFLqcVyaHYYY4VSQD80k6ZWSI5BuyyqOK3Qpk1gNn
YpW130JLIyDZr1JOsO//zRcpgI324bDVhN22B9kT7ED9E+LD76i1S0ix3DPnVi3D
GZ0SUkqSr8LKGlvjHWmbqaLl5YUyB8ktys2r6fwSSUeWvUSOAO4U/5yqavkmoMFx
tHIbHElyDWSaA2+ecI1ka/NmhobPGju3zAvHDXJQ6Xk5AM0hxnyiaBXt2KqJe9Ti
EVNX6j/W6RDx6pFPzrYT0hxMVgI9eZlfKsfpkVMWDBqyJE1VXNJ/jS1LwhYEZoiA
r3RVlpAbu5qLlnK+BGseSmXVILZA1F/JWLRESghFf33ocXxG/dn0+tid7bUQZtJ+
UELy+nHKpmY6/FriMSPnqbWRpYEyJYupiRF49oFptVSLs2AsbMATjmKVtEALYDgn
BOIU8CI1MZYnR6LiMUPYKNFn6p9Wv16fLsH+P+jGZDR9G33wdjFn1ED5Bexvg9Uq
Dq9/o4M9xU+lZpAPwWKKGNiZ2cwvNfwZGYiqAtEQPiqvYv/bfit8D8SH+Wg3/Qsf
T44Psgwxu0xjUzq+DhOGg7DNOVJnbHnHQq22Oyny4Quv81w9UIMvbnBoqgM3HcA7
duOt1D4PnGJnXmXqlfqqHVLDK0EKRYA+DX8a0JzF1H8te7/SCtVjAe18w5hHBvw0
1LTo2pdb4kqehhKxgYaQjy4Fy233MIlLFYE7gMKKPjEMlaSFDO4JdfmLfbEKh9uv
xgBHLx1sEEvUShaI8EeI3Y/Eqgx3exN0LmMOPVVw7LZJjN+HlFY2V561Ekp+X8p1
vBR5STQY7xPGaLaTCbpXgHRonwAk7N+FNZJshtA52izLmwKK0aSDSfX5Ghf8VpPr
QZrMhDn4f2mRobs5CdMH66Nx6eor/6/VVTYxRRMEUAxz4HZjwhI6CQMuqSvS35rg
PUEEB6VuFohdYlroR9o6l4XkUNZVqkXMkp651euGgwvT4wo9p9Us0rbuUaiFRqx3
nehtrUlYpE8vWHILhB8+dvb4E2d3R72XS0CCXW1Qdcv4s1X7duBsla6rbn1HsCkw
oElXgc8c3POCrX47AFeWs3hM3Q+XNNBqi9Rta2UIgO62gkNAdN9wjPoix1EOzx6o
X6qF2eyXjtuOVoY1fjdAYGBqgDmz15jYDAedJts5nEmiJ4iLd3cLWe/8BUqTSpi1
zCcLrwmSLeUH9bbCep6yPxtouPso9eWMJ/ybGZpOgHEQccv64kePq/imnt/R1by3
WJtsRv1haszM805tGREu9cFmEyJyb+735lutBdghfWokpOQohLg6o9wzMiaJhnDM
n3+3OqXb39ljwTfuFRGuDQUQRd2X7pVQy5k+DjhhCQ9xGFRJ/YZHxOac2j41rMQM
35J3rPOBimWNeCjuUvUUwMuwokWUq1LZEoYtjfXBDWht4nUlaKAu7FmiQy9kul1n
wK55fULsXU+ZrBmJABwsPl4m5J/0faTgKX0nNXrwpfY9Rbw9Q8BlvE+5lnV1oHsr
AQG79CNoM91k2O4H7eJ2zpk1QLmEv1EEv1vS5Q228Yu5+ih2q/xUVEOQQ1yN1KCo
pmd1wbDFaEqhesnkFQXhFb7J1j6g3zzaJQR7aTqmFSgfGtgrhPnL22ELK/yR7OyW
dnaECxCOemxTlUkwcdnUPSoIEVQH4pJR19dxx03+lyxZ84LUdnT1SUNSX/QoWkpM
WYAJV6H1hY1pMyxBKekfmzgPX2IErlWrEHVNMCbLoPE4BkixsEqAJHcFRPD5x6hc
e5eQCVF5zubb6CJOqMGL848O/SQ+U8mGbXhCfOfTo5A2KhQpnl3uBll8YAykmRKQ
hSNgdgjcaxRNrjZSDFrecb//HkQtP8oXfrYq53v1vaVinaSFjtLIiD628VbMgDvb
Ti/Sc54LFgffMtrZ34HcZT8QSx2BJqc356S1vV30TDVyAzh4hspsHmXtfuKP23xt
AV0SrUpn40KSZCO+xOa03x7hwXqgKYdKOvRdSm0JNrywqIeQn0iZh3mx7UO69CI3
Bk6ed+xbM2HCJ4WyuHkf80JvRd+XV0dko798Y/4a5ta9zlEyUO/pZ6cijqYZLQpH
Wg6sp4S47JG3Q7WBqG1Q0wrwsqoVPjfXMQSOJ/YT+ZAfL5QdtDOKaGeRWcp8ZYUc
cNbjdixCP5o11Gma2yNTcvS1oU0SxvvKV7LBJbO2P32HU8KKlm2aIA9Inh3TLHZW
X89sAy0El6gF56ECMXLLBGubXTyXSE3aQXUrr8xHaP2EGT2xi6odX71uMYGT9tYc
RXHPiiYUadlMZNcuxGWf69Jyw+ZV2Njv2iHNFkatz9Sh4tflxpk6IAndqHh0e2xu
W1SkrhHGVPaKWyyxKA/MaACr7G0dx55yKSmKEUZrl5XBXzjx82stkKdxHYB9U47W
wNSQ4LK9Dq78oM9IJ/VQLZVQ8uPJszFGF1Ek38Rxwqo5cjdomWn19wCsc9ENtZB8
mlNkEIn7RkYvVFIgzDpfXAYl5Y4JaOxbmfQXHeODWVUNq7yHL1bcdN+saLuMxdWP
huLlJz7dNG3DR8t1LBFeRRLc0xlmigLR7UyZJn9J3vmMk6dZuMkEPUyWWN+nDwbC
4nGM2lzZgM6MAyynJrCQlCjdLd2a4OE7mRvLCfWZHrKVIAvtrQUA8JyeH5lWArCi
qF0zCaeETjseNTq5uG74TO5JYeURC289pX9buSQl3qcgEBtEy3UOecGrruzkcE+N
qvgQ++7Olp3GXeG0ZbBudSoNF0M2dcesGviWmiykxy2s26OwEIM01oBWyt4b7yYM
tyACFtZw99lPZSW3SlvU9WYuLTRxfQL5hhBGVx8I0UFxpAjKhQhMbp5p0nNV5M2G
s2hLgIRtnyl9GgHPK+0rtzFeIUrtzzUTTOvdGwPKYe1xYHQ5MH/SbzvCFkeyiot9
07Yq0GGYVgGUFytRfGdbej4mPkM5Y8TXEzkKt/ggaoRug1hnEAG0giadse9KIrp4
F7v16fVmuXsrdA6a0rArIlUEfMgaRMJk22s6zrcNKAQWNjcS1ueY0dpJeZSTL/1S
IquO9kpPQLbjs9MyFTC+S/de++HoSIuCpXVJKLVQIi3dy06CXfjX4VJ12QpgXFbu
Zg3QOQZgYJ/X634D8oBNv7fZUQldZflbQVV9wywMUSeZicojg5+c8WQS9pyyiPwX
dXQqChz8xnjGnD8rKyvGZMGo6VwJnbQVsgUm497qnIv3ATuEneekIHQnkCeKI2I7
S7bpTnA+zVBo/z3niLfLjRubYI6S+tjpCwBcB7hVpoCzsBhEqeIkx3N2CCsOQCjF
7ea5p+viBPf7Luuv0tO5mRtykpHl7j+4HV9OP+tHs4LJ2DdflcwyC8nCl7hyfL7L
H4UJdDgcq/WNlyW1yEZFKAtHcAmgVUfFDDCj+N9VTnh7YkcflypAoJw4hpJ3vUyO
i6TnAlsWlUJFU9zlAtd025iDIZr2s1P8OZD9+gE5jgm5LQ3epFchWBXeouFjLOVE
U0rjr5RCA++D5Eo+KhvH9foO8mtuCa9h+3cjs6Q/VlbdPWMfNnJL0dubFArq0MBc
Q5oQ1HRVDfSmnDkpGXZsEuG7m/vqsZDKMd2FBbF7KBzvj66yZsUC03O7nbh/QdWv
eTLGt0GKFG0LWJ9LY3FwJCWKibEunqi5SjyV08n8LXRV/vxYIxaAcIqnm7fvhnOn
lBjFk9T9xf3TfwhRn9NUwcWnEREemfg9udE9KdZOuUnMnvxNJjVkFHRAcoL2mk0s
EGM7asc/ptg4w7I2HfuxtVE8qGj7miBnwmpkg0q7AtNAotuLYiTqt4WBTSJCKRFU
h05qp1Kdiw0Lrf+xX6BzaNPjFvXkf0ZuP0DR1tBLC85lkwK/8NNfFYaTuwo5BWD6
fuQiZQ864z5tEjORY+pMZEurRICqjlZzmp/Cj6zZMa0tctjFS8NpGhG8kq9rhnod
1d4vykApGGWiLb9mU5ND0DF4Gr6YujzdokwDLHfDD9hF72juD+ovSS5o3ZTYJzJJ
APOu+uMa0A9S9TbZQhV1nlIEjzBxjuOznAzKgYiyc/8zq5c1QwWypWUmTUYJR9pW
vH3AGXVOT/OxaN8FylgmGwt90TQIBTACClk4ovj1BoNeMbnOQNJsB39glPX8qAhI
OprkOzD40+p7gZTQkYHEtMJq2WN2f2e5259QxDx0Y+Eo4Nkw7SDdRn4rfs6uevz1
DHbAulUiXUDX0P3HtQEdKOx4wMjYClLFBVae/63comKF+hnIctFba5dnQXKseFzg
yls04cI/s4us0p9vZvKwFNMUPXnGOOCndJb/WBVhJ8y97jULpTDVrxC1iZ6uiKEO
hqt4Y0uF5QQ9ISUsX+/TdNQKCw9C5OE/6YXIrDVsupzd6zAgm/AOilz1gDpJyqP8
aZgqtOJYM0LCa7jhfB/oIF41iTWxe9pJo1zERzHUa++DxGdXwJIxD2NJFyzIarXs
hcyGG+HW/Ip0ti/+AbX8FoxYF11V23mkdVdQueeCKaWA0ehbk5D1UsqKax2+ishP
z6K41FoAql6CyYrkNL2ja4O2e1LbRzaZc+KEPzBanh0y2VqdAN+Z3QeDISI9yu/1
oL1JoYXB+uPfe7aApOyyIGxXeJA+NQ8RZuzvmoOjKlzqbG6GRKjvI548GF8nJ/6l
DWVazR7qzruWUKNqyK9lYtd8x0i3GI9fJF+jA1Q2nyjs+1ZxWYUi5BZTeBZYAwtE
pvVh9kUE+0mpK9gqs+0haRFlbbRQXWwLp+NpTX2eYXMi3hAdgsxPSEjskzJrDHBv
gUuKAKoVO+zuRr7NzVW3vw0hRtIjRMnVeQeRVQSOpljfoDndh4uxlON8bHRYXM1a
6mzcJOQekNMF9NNkhvHOeUTjYl9q7PgFi6YLjs2ftZ+BqCOTuBAIpE3yqp01gKt3
Fb1VYQjTMqXvShNa1qRtmB2QF34Ahg1v7hSsCoc/fiev6L/qSD4CvdmB1g6yLWMA
LCv1FPnw0FJ9zqtK9UvZNsc2lK30IxAUHGp2WeuYQfLUF6Dzqs5Pau2GU3G5N2tA
vrH4Oh0jamfz1NzXltkVMhB0ShSUCGy9bNO1b4YLmTjevbsfJ6K5Kj/EeIFN5v8T
7EFTQ5hhKYm/ZSfv4d87/oXsYCIDvFk8jH0YjXXcV/06BGniJfb1rN4R5k0SzwFP
S9A9KFpU3+zNjBlXy78ZkszJtuJiJJfdPjH5ntySdJgUa1D4arFXlZHsfolJFN5l
mVaf9kwVzUtfvEVTmTdofFMdE6yZ5Sz6jDwZwE6moAg4KG3xsy3SYk+IcXnFkrlL
P6CPJ8m+pfnIzRxyJe7UQfXo/1WTp1fbz+T3QuCaeWR+n3Pw57odVj/pomrCOa/s
sbu8oIWQRI/9IJ5mlS0BuNdtkRBruujOTs77IZp6HGHjhxR270SPN07QXd+be0Vo
k79oYpSJT/Z0pIh6lx50uvuJNKJY1HnuIwHvRTBEU8Cy7Cj1rDRTzYi36UuV8ScZ
7F9InOZQzyX76702/PZ71Pjy2RYixthYB8SyhTYBC/H8o0JFI/67ouEii0aLtMPw
39nawkjkw0YKKKAuHrgK6NHa9XqfRccZDsjS9I+faGdTsIo8P9ESCrylEWRT9eyC
eZKovlCwWvScebQTUxbpkGmR13s5+wCNcR3s+T1nesiTySggS6WulEYckX8yd8C2
Kj4ApRTIalrHuTcUgJOp/Qctl2PbMI5Sjoa38nz5aPlqlnYmoXwHQGm/Z71jXSBK
tHjLf9xTFoW4wEkS+aPAWi1rh58lP7XBmDmIrwV18F6L94BkX1MXyGE1Zh29ZjmZ
97xbwWyH0W/I/T8TNNYZ7/NTnZ+UpOWZx14D24IH9LUumWBesXrDdjcM3Ljcy+rm
eNHnJmmnBAUXePr2ghqNy4PUEH3IqQ4cYkoUOmoQnRzUSIuyr6O5ussBkTzzy04g
g6wkNkEjEoNRVzLAUpmyjBB/sDbY8rlOi0iZoFnhbocvSyPRhFsUiNnjAR420HJH
k/zXd8zFursVZ8uNLnTzJUzDkdWthpvIeXxMQZDRtYZEUMDtxcsbtP76gu225FVB
QDQQWIz8eQ1qtdROwY6EqiUnaFO//XQiZx1G1n+pSiIbBzlJF0fsRCR/vbcZk5T0
Qr17Hc6ZULJaQNdft2KBZtpUzfL4eoPumhSNMdBrzZW1/gp39mvUDSZUUtycfDol
g2vZ8oRIl8EjwoYxR/7boB6mmDABAo1zsJz34sdz/AAWaJMHSglpfzIWCccIeqtZ
MopfXPtqlyCHo8w5Yr9zj1IVSiLcoU6WexoKgVTKv9DjYNsVH9jd5/8rvqMajzwa
tHwRlIq1iFH243krRbn8j7vWP7JbDYG5/f5TDAPpgBonxtrG6MX2DuPiYPxTSPgu
yodEdRR04nLf01Ry1RLENsnhnq0nJDNYGhGaUKxteZ1IAyQBspir/1Y3K4hsgHop
hlt1Z7evTxDr6lehPWVAktHmXxY7SiIYJ7pwW2yCUY+bqFlP//8l11EEmTbPPOqV
kvxIf6U4sGUdiO3lTiAQKTyWIFOr3yugAvmHEVfndkNSruSRYP3NYvcBg/+YOhtq
/zJ7cvcDGlCASYeGxvy5jf6LROjEhka5hfeP167hqjSbW21eVvO1OOVC51mTDz5x
QMggqPPFj/7f44HXy9uyDopOwQ5U2xHz6pyqBmXmnC9rB/OUoVsgvkWbv5oLV4Yy
wAwgzy67DyEti8E/8rsva9DYbxqUakD9URTMjLTEJlrWWSFBgD+feEWkm/+y5GBi
jBFU68JZxuxpWojtxdQc1sIvXsptz2Ox5xdNmlfkQBaCHsVLkL0tH3bSNVSa6N2I
sMIXMBoUVXDonyQbRqEn+qck45YZmUbTC7R1d3mgieUrFFBEdKkDxfUhZ3feAyyX
cKQ8oYWYc82l8PTyWretyZeBTwwVgDXqotZRjDmmSWtCuXnCPPMzb9c57gzNm8KF
cqCDyJiKJ0gowcCGZ4v8gp4c+otD1RfhI18vOSK86YAtUqyQ/bctlwf0TVJGrtWk
aKc9w1jLCIWBbPvLoExmJRUWDyQhZIjGIA3FaTsjFxteZp2PrvoR6gcOWWWeyieT
7wbMtWgIYHhQo3CTxYHQsCanxbZbiNJieHnbckr9EDqKGPGw6ocDkTTfQZjy1doQ
BrDfuo6yBt+Az/gNb6jlpl/UUebcjDenT3t9D0iam//rgKeItFTqEruGktqkzQye
qWaEyKXNWnAv7ps3TCc+KvTSEIj/Ei+oA5m6p4qalb0tu2WB5D90E0JxPLsE9mqT
uZQUmm34UMXV4KQ/fElmjhNZB2kPV38/O6HbI38l2rwqTT+QGY0+L7gc84yW74h3
7d/4rBep3Ei2QbRZ/osB524S9iQ6z6wmJJn/1CDGhjzvyHBnVRacYJbLyrs7nHrA
xpXcUCWUldn3XofRWW8tvqlj8tjICECfHrLxhSFWnGtz6GmoOZ/3+JJpwo0msA6E
rcuVE9UN3wOqIjLbYTRqmk5kfR1qAv83v94prPrkWARb49+af9pRsEDPgX/R4kN5
UWi1juQBDThPTNNQ523SNuk5TsZRZakViMFyrxkixf4aeyPFrVcEnwpJ19tjCAtR
wqE8UPt2SA8aXzkWq44vhgY4E+LTKfuA07y+LkEQTUQ+K/qH7l7SDgA1dmMzOpQy
P4EmpH+90qEmn+aFEeg2rd5zZz5OKIVyUdFuiG2d9CW2B6h8KvdfxSiJJEpQx67h
jwIVl8qQfNKVvbUeoDudSzYWprSI6q0rIBZUJnbVeuIOzhFTBlSx6upQ4C6REH0c
amD/5zb3MY2s3yTrGnyK9r7dtyU384sWFWYqU8LIB05pCUdrkDTcCcqlHlHUG2t0
jBA2IwgVKbtR85pIs+rn7cDbTYo0OeFR8srfzxNJUW8B0BFHCoUxU/QGcLugkc3V
FPWbMToeUjTWiKzu/5OfMUNEnNxl5LoHtLSPgJ8eyOCqvHf3W3Mt6HAfGe96ujJr
q17RQiwks+O6EE9vogjpBQ0MODs3u4CQfDxXb6NlktQvP/8Qfh4AdoogPIGY1oJs
CAnarzsCBR53bZMICQiGNyJFrfeUH3CPDLvIvw3AogO8iVxUoB8v5/jXCiHzvySe
MOZrPe4dbGEpAoeQflg3qtBBPgFbgeFzdl/STi8YLrFWL0aAYdQLzgZTprPvrW0K
RLbjHB9SG1C6FSOUHpTqV/0ewnmR1tIUQEiWXk87F+UNuvNG2r1PsZZIzWaCx80T
nabIMrKe/1Y8ovoL59e9WCG/3BVKqmOrEgVBW+ZXEmvsZYFW7JqQlvlyH/y7+66s
npyWvtGgm6ROyxdMQNVy/fmhH6GykMESvaAPaJDbLgqYEPeFG4y4GywhyLEVckTM
nXml2xPSb3VxtqUlHAksnfVt5Vj2CGYo5JDfmwMv/Tx+JD84ETEOb5c/ZHAyQ3AI
rF14H3D1knks+efsBwC+0b6j4isN+Es6ruqEvI7dfa0RvMfYu2em75zVA69YQXlG
JRaGvP24zf+kA/nLWl7ObMJZCgQlLSd2aZBD9TrrrjyypX54CUhndPLLWaJB6wxr
a/UWo/XKDxOP4izFj/Ib/8dNhB+vH0WTr146UbPkAirbFXOY+8dPVcgJbsXF32RC
UwBTZcdmfi3D1V56a+GHEjovRJtHitKCNqzsqz3btd73BhbrTFfdl2ZaPKj/FoIM
Iaa43Xg4qr9W4rMYIL76WL9qPJxRh1gHFlk9U64TExt1MtoJ7+D6lxJh57GbcWuU
keBI+UDurwlpPXwAWPBeLxlYof7T19hy48qeyHjxgoJBzOsVlCikpeykubPq2Dwi
+IokfIqwvfvilihefm8a42pdagewmNUn5hxTfkCz20J6KPHfYaS1s2YlebnYcuI9
ziAkS4SOlTBkSouc1ROSHwf43cLd8l0X/z4Xi6exvbyjzd4egD4uvxBJBoz0gmVw
U8UWAJG8fYJmKwbdtoaMLw8RMqYlOjXiuiPIgJU6Fte060iDdm4vuzj8ohPLWgIF
pvQG97bMm88lNs5hA9giuNFzsIwvJQDDzjNVIxQtPSWW6MzBVmff3Vu8vYnkr3o9
S3lIf9/dm2mS0H709wK4VlkXUPXvMo58JrRe9TfeEybOAZ933BUVntCF2hWgd/TY
UL29zN0GEHQ79Uznv1HRjMGW9Mp4bTnQrfMXhLDHyny4UzEHiUyFHJGKmR+hissv
za9bAfDiu1jhUMO+IBqXCGnP+yAST7nEqxnayN/7TqM717lfK58SuSA3vV5ZZdNX
x8ofBLOrV7H9SDoOI8YR7gSLBIBSXrSb54UTtqSgDFnkSzyeUFmTj/azltiFodKU
mpa23Yuci+VvYK0SktHyfDJSNh/o+Vvh0bzU+zOUw8Qx9hjXksm/KdBMLhoCauYG
wVZM0GK0ueK7Sja01w8v0iPPb530MJTWJBFA2t/CbpH4e4otNMG8SYfBDhXK18K4
5nwFd6ADvdbOVS5Cu696vKNG3pUol42zWXLOj9A3bFgUdUVbmk/CCXiKL67LZuVm
7H4+jN7JcCstc+1U09l2RW5tbIPMZuCy8JFu9earse1mV3aqZUPKsXK3ZRVr24qL
dV84b1mlc3PrglCd/HOgFp1AmsVaKoR/B/sCicgNUP9eVNTzT4DBNIuJfGse6KnW
E7fCAeIssKr3lMPoMRa83ZVpE3cehD5tQGquYjZdpTWRz9EA2NUNgKKpv9mwS26c
FunrddTlJWlVBTnWoGJ+7RzhYl5uFDrxGz+6F3y7bqDQVQV/pbVYLccnLJci6mbt
L90PuzLBnuzynDB0al8ZzbwFy77z7gZ9eOPh1KX/DjHL+h4G92PUPsZT+tuTs74l
GHNP5zEBA8pFtCTajGDdjWnFqH4bBTaUXFauGwkoJLtLuq21XwB29gIIi5FNIZLs
Krty2qCNfuLrVO3XP6XgD0rOnjpaT9oupybqZ+EYGIi4qZ++28geH2lbkRdrpMQ8
y/hTTWVoUGPd9ufrdn/L9QtoMyHkt7w62h+cYqvqAsbWhgac/HPevyde2Aghztre
RcszbwxzGdkUcHkoXzXglPJX7w+wjhAolKTIMO8Rc7OgcfCqSMV3Eg3blPkwBgtC
Wps9MvIOUxPsNo+kT8vlHRWqPz+59sQacF5wpKkeA1OYsaUKh2l2z/Fz/DWv1n/G
9e4vGEvr/5kXjkP81UDSq5Q9npLKaKZheBFLfyfo8BdXuWLGphjx4EuBw6w3uqBL
UVncFg2zhdJ1CMW11tXuwZsHnJSn+gbwn43xb0BNGHUCpR4y2sYV4lk1biwFHCWo
YFe2+RXb9I8ZNTNEXNJDaFUWUK0cFaL+DFCfqq1Tno27sMBOiakN/y2SdcBVsV/q
oul8j+caJD8kllrq+UfFgIMh9TJyNhD2Kv5v1+0ThevexoA6pefud5ktrb/Ik/ew
MuB0vn1ncGXzbIlfkkrak6CKZ58qfNJWL+ZtL21lTfhUyXcc79Du0PYWE4KQFWHm
HI4IqbhxVOksU/l+Xg4NWDOcE+zBil63hmCK7Sl2EQhOTXGBpz7Cr01JZOu+6+Nl
fidUyZ0saadKXSeagshmTMga7/5XryewVLb+FITRYSLRHLUKLJ/5j6n/kdJoU58y
VphIx73AsIfLWFI5HkNMz3lJELzxZBNE6GYmuRszhpFtTIiHcbIzc2KZ4uw6v5jE
dpqyH1MdOoNiKhPMjZSXn8D0jO1PKGSnlBdfv4dBI7BkadFX93fIOxCY3aeWiUGN
pJVQEYSY6UPIZD3cmqCgGy1a5f4nzG5MUV9EHjRf6cNXA0U/u8TIh8CbUB7lviZA
p8NRDJCzaxS5zoS07laC9WHqRaCb/vYS+LB3JQgMLyYeLsjozatW2HrxmfSG66As
w7pYaLEtKH7BA4Ejqe65FGJvbsVKvP/PA3zcJgnL2MuVrTF3/56A48zxssn52lSD
I4E5B9RHUORDz1m3HG8n3DkPlWomZnEkg5eE1a/gQ4bTz3VUy9gkQwZ5VsFSU0MX
GFZdinVUQfyYEDlGiCbw/bX0mF1kfgeNemV+Q/x6tkv7sbHbRWyQQzAZ+qWMtMFV
jsMWslgPvkuGBTdICPIzsgBNM7AgLlh6stCVH/SfpbL/6vY6Hwq9uYqZ50hzUPfu
NwZy9yDWoVBNmxfDdnOPP8ub6grMJhIQNx1bCZQCiWfdvUyLsGV04nxbD9eg4Ih9
Djxn/ihr29ZpmgFQQ1AAUdEWiFF04OVLbewWgwCuET7Wow1b8W/oDqIdfTRrJ5FH
8H+Gzy7tZcRvYnWMuEnUGwaaY8o4Y3YpRImSlp6Vjm6GrS3o+X+ntZQAoCtllc70
rNfSh1xSd0G8ez77J4RJ1C2BRTsN04j+pLclV2/iG1pqPuN4ek7nzUVCQRRgwhaM
/jQFa0du0RSX2iWg3mA3/Vx70f6XwzBsu8HDmSG/j3y9kzqpiwzr0ltbnEHlR5UX
WRnSgx/l7Wm4k3WNVIHL5DM2MKuNvcHLBzXV0HIno7rwJ6NcnCt2I/wSWy63Z80t
AEVTrzzMjejxRdvlA3xwbOYCV4+NO6l0BLhiasrgjYFj9WPrU58ProIseGmOAVNs
t44BlHEEo0akmuMGLqA+aYLRbDG1YjyqdK3RgFyWpk6dAm4jlKqcOl4tCkV7Dsoo
q5PaVFr8SpATsRjcb4X7rKrAjmc2yz0mdJ/qPGqx9GOLrvlJX9+rQjYCd50EcFDV
XNTEhb9cWH5IX5MqlCnM8M2pMfpZl3oGi2Xgu6lG1vcmD/D9hWlQRZ1uWsXGO1C/
2adrhnBDBpTidooTsOhob8bdedEn93ZeHUa6hhiKYfwKtWqEJDXO7upk7UPjHcz2
luctDxSIlbl9Ms6I5XJFexM3W+TKEoPxHiqJKZgpafzpmSwyufExlhJdLOQm6Bx1
WAmc8ehyf7TPmQMCSEARtx87OkWCCJbckH7JnSmzXlNL33V1R+I0XcDwtXwHk1c6
RBE4TNTa3mHN9BKptvQ/nS7jBK1cy0eGTVyPGe9QISCNs/cYbTF5CAsRLHGb8fhE
sNeBQXDc00fgQm1V4sRsl06DHR1oWoQjAAGiXlN3Eop50NSZmSwrBXWhD3Mi+hkh
HIgSg671BowcyglNaqIDrxTXM2MY2zvEzrPmzNt+kTwuxeDmMbupkalzSvLiOcfR
s+TDnEAzMZ7b2qBy9OfExQJU4P99hYT6nyZuZ6kSTSfWM9aSMWQdENK2A+qsD4Vl
IJa5UhDgKaBQonZMe0IKFh2e8/rmQkAEtcuUe33IKQhq3WQj5FUg0jVaBvv1QhXM
r5QCzALvtAB1STSyJh0qSpunl4wmTC4X8ufNBAElOyqfrTn3vQSRhinL9D6wElGQ
vtypwzxymXM1OZTsTVjy5FMbmjW/FdaCRwNfn1Q1GET4oyqrrtmleaj8Zn2Ssc3A
tI5bibsOQGIUAaHYhuc2DeznCkyxNNdnZhSGov4HLQ/UMBzvis5Pivaf4exHXC9/
xAxP11ESI+cV6H+aXP9eL0AoBB7UpRbs3a6+jdLCDXA39HgU1xhXEsjWyT/qNDoj
a+DRCu++Tl6N9TlBO6p/qPmug4feCLOmZqwOmfbY6zlkM5UfThtySMAy7ZSUY3Jw
oimvfZqbN1zhCNgrZnjhkxkUIoUjCchZ9xd12/wHzdJqsjp+wB2/FcFKMOCWhzEg
UkCPLhvWUWdm9t2EWsFA0gtnPb7iu+fDMifLmfHEXc3vKYmfAJWWgmB/3XbEo8gZ
/QqE9/vweFTHVQ1AbkaFpF2cpu70szVamUbFWx0dPsKU/41tInCbh5X9wmj/ROKr
x/0nQo60O4xYKHFMvPJtZa4CnZWXPhp6Xus5JqigAdUgTdYe+O3dJBiZ4Dok8H4+
IVDSIHo24Vr1D2/Zk7DyzdA0m/A517DpYDrMEykom376OAELMcdf9F/ah4biT+h2
LPsLVdKFczC1LJfa2Nj4/pIeo2YgaVFYoJQAJzDMQqeZSLHhDcuqrThNQ9vjlhxe
MXoPXFh0SYLq0+67PqEdPjMG0+3lFm8PqQ3b3v0dVSNJ3p8A+G2GDbojdfT4PS2d
sggMs4knaoShkgHByRIeW4lVFCA3YihLbQepZUohShC2uRjDzBG80n70K/rpTjku
uWPOpTVzEb8CyK9W4Yf4U31pV8BrcaLVmEUEn+9becLCOGLVNjNb6u/kSBs18vuG
2Aj7cJEKklDzWPsz1DT2yKAJWPR1TFj42cNelwFNh0CVQ4e6wzi7Ta2lCFWdLWtw
CtarkoKDGpiB8tG7Tr6nu6kga6G3NOO76thfhTo4wND6elfp2pqc1VS3eoHexyEQ
AOTAmsiKZBRWE8dzmeljaoHoelkNdTVLaLiubE5pg5cJroFc3cRAJHtXh7T/rYRg
cY4n2DZbnQCRzoz8ta0uefkM8onJCi/MmicHCk/WZDBaA5fC+dzGDTUl4Jh93Yda
aIdOOxpCwKcD45YH0wI+pJL+0ThtCt518vx7GrH5n/3W0X94G1d/ufWKKgV0+faS
BNMdhOc9P75raGOBTKtU2EUa6yIMu20yshQJjKwiceGdTzn79L5XaHrKo13kWSjV
241p4PBLvxOB9znpbbNPliHlx12DMvd3szfKPKEejUXf10J1MfuSrvMDtnynZpDm
rerhhbpu/9i9CbMSD3nTVdozDkS8fOxGxWTXY1VQFcDAZYPVhvYf25vo30OVfnKN
owPWjdtujYI1xgsfb0n75Q0VJ+xEvz2dVtLoe0khbhVqc+w2eXmrA/bP3PMstiLC
4QcSvboMVqV46vt9OLBW/7u2vvg86jNBjg5D0bF3fCotnQ07PXv1ADy/FMBrGRVb
1EBHj1kZNAcQqM0LDmnOcy+sUhaZ4cWtt9JI+oARGcBQbZlnKeLxgPWYkSOOlk35
cWXduUp5dIn6twFom7iHH5hTvBTxKPENN8SvXwrANqEpwWRF1s000jV0Mmbkoya9
L+9ppgV+obTVxhlHoJcpLK96JS/WhdxYkgs1y0Vtt8boHdnAAUmPwY0cL4ohdI68
ZM5r+/JD4TKlxK6ufz3c95BeDMvJq5Hq40r9GtJC7qP6toNRdZTf4yfaO0ycRGCv
3kgR3mRwpSHRVIxanA2mJZaqHSvPlVG/F3UQXetUxOO8Mfx91x4zPDYg69aWrRRn
qMAMQN5S4hGEVrImov/IgNzWr8tZfEIVv2Crt+yPs14aaB+/SnJLZW1HLzpFx76P
TNl6Bz7577+CbcBC67u1YYBeQNplD+y4eYPSv98n71gjUKTCkrSFCgdVHNC7K1VZ
3M5p3S+8EYpvrRQQIex+9hJkuCanD3iIuVNJ4k5yAqWQ+U6gLvxIl3af+TMJCclW
feSGEnttDjbEuInbU5w2SyXcmnn2r0OktwloxM/4j8VoDidVWtNPxx2kgVHUBVSl
PSFSYXP08SMCS81ghvwjFOx7YRuAyE6rf+oNpu6qKpQbmpoYXxxjb5dwtMRhl8JD
wnmAR97EgEuip1fOOYLajbo3xs//ebNiIWpztrYnc6uHbyQ/LiI1pJOMXk7GRQYq
PmsghvHdiqzIW1JKyQLfoYxqxIfLHOj7lQOv5HPFTByKZ7iAZAcRs7R9B0T7xNAB
ULlviN+kxuslketCzAyVCT5tBstaCECfVVM4/IUnGrZuYvzL3W29CE+0Ri7hqMts
oKhyc7KsOnHbdwSZnVM/sahl7DKcSklHs8gRBLbytX+uCjAcKPslCVni5pPbm3AD
aFO1HiS+/ttrH1cd2aBRnJ6aLgdaxy/xJYH4hKmIkGlyiwam5PVK+4crUqR+odhK
YqAxRGy1clOBRZ2+aN5uY9IJqfqyITPvoyQ3vcgFfBwgM8fagU39OjjxmrC92Qkc
rFjg6hhm3insxFH7kjO1zV5P2ie+6aYA9draaqxN4F349H8Scz+YbExb+v7zxggf
WA1TwDakx0vLZ/X3sSzHVMVjbLLP6hMtDvAzXNe4/cR/lWpJ6K7Ip1/qHfyL4zbV
r1ygqoBv2Ae2MeJR1wpMGV64Q8YcO6njXPWybPwiOfM3Td206OvOQ5aL/CkpOXx/
K2lZ4qYu/z0mS5SvoZCT16iYPyJrJRycHy//6KUG18hveg/1l/IXqI0/dE2hYVJR
rUGdOUD24ZOEPdbDwfZA6W2sL8sv+KrzUaQ1vWyKf7lNefjzqUJtLnHgQvbJW9Tm
uNcBy2dxhwhq0pMHRgNxtiMer4aK5JEqEnD7rn2RK9yOif9g6RdKDQQv+g63g/7s
uG1CRZrArsmDU3JblyYklBCCMQwrS6gUmjKyl34P3zeKOdvsF40yzmb19c8dLSSB
HAtSgKMfcdliwfIqWmW5L4/O1L2+4jIvaRjBF+FdIY8tlp+5lOFo3WQmWr8AXZA/
OP5RBUoIMkaZze1/PKaDmgX3bUlrKujIED8hESSq6QbynHj7Ws8fXIFWONXt4eDG
TwHkaIkzlSgF6KBWx1fDc/8hpVM725JIwSdfxy5sC1m3q35Z3yKVec1VPSilmA09
k9/IHGutND6U7z8oysukCFgMKjWcomWcUnRBGHxUa5U99+w6QbKT5mFk0mPGmeTZ
Dv2w00R641Y5oADcIEAEUpF38Z/xb+EnAeySi2zOYqwHR/zHMIJb/X2SM+jtD6wR
KXp1MB+AXFglQGyu2TDJ/tHcGUWtsR/aXfilmbs1edidq4VGiW8/mQHB+exSPd7B
1hn3Wyz6FrhJd+IJwMsV8R+YvEgKhn8Q0XstkVZHyv+wTj7d7CmQw3DRwfDxtHNg
Iz8VZSEGIjmOwp1m/scLBA1bKCNm4pD9XX0s8e2I34gtkzaG6NGuDXecwExNONoN
SCQcFJuWAESPxVf6ixOKRXUK1ujetMOqIHQxDOUt9kpPX1fjOCRvQzBpw/kJSDl6
8YpyNbLLvFdzn6rp4O8Zd1LTHLw6iTmaY8MJZ/c7bLTesGy+lVB1UHbjmkWbMN5Y
ORLo4QBAjqfcG79hchnGJCatgqNTck10I4x6szziSXbXEv7k4cZBVoncSeFz+/cb
oTkkP2VscGR8gBBUJBmB6jGFqhVxqgF+a+ZIdPo8rNGGfe56Uwx7HEI6QEqROQqR
lQTgL/LNB2ChWKNQehe4dE7nviSHBrDZokmJObA7ggH680PLaMJrBfCpOnBy0gPA
kRwJgBa4Lrm0QloNnhVfQ3UIdOSe0fVTi1MJ++UlDgH0LnZSipz42Kx0jt/nIi45
WXa8tbXCuCwhU7571POupfHfTXC54qjNl0BgCDU5agJSFDegNnrV1lTDFM/fXhwn
BR3IsPKx+IVhYVWSnfmlIRfdBlU0M9PB3kjvMw1dg+DaHe6kp3fm8BVExbjPMHGe
geWY+JeNOcN1FpZM/PUc5XCQXRuagrLGPcfQcwGIaINeRA3ujKMXXhdy5IdVKfeS
+ZQL/VuY7TqFYBq9NBlGkhp/j+uWzt6yd/0SnSWYnkpikUElH8W64pf/Y0Yrdy1c
aMneX/leI2HqZJTCMS+eda8f7X7mlCNDzfA5sK7ZujPHSlfmuFWLSr3q9aTK0hLO
VQCgnKiyI+1WiZixCXW11M/iWpmINSRRqq7FNBCkrMKySWu7+yCr3ibIhU8R1j0e
JXukzTpcxXaE1S9/yAUiAXeBjBS4XGK7PS0kU/d1nwuQDrL40oVS54NvqEsw93sj
xN9a96BzN3AuzmI8NUuVDOkCoZ97SNJszHOh02Mb42fIGDd7dJKEG0giPZ52vXXK
M1Bh0qHHALhmQFZdOn/lgppKuhXlT0kuJSHbn8a3kPdDqoPkmRWNa+bA0/IFP1dp
IA8BPneUihPqcDXlbdDwFi5bkVqiySfX194/kIAq2tyU6B3wNJwhscdRne1ta8k+
ww6/6gOjRgtKcetifaJQRo6q77dcDS8Wtt9bZtHK7Qund8gXlT3VVU8aYReky1dg
pIKHZoyIGGfx1ypYthuepwdaFcbp8meDociERnxYV1aFHvYxWCIVMjVWxgBRzhtl
S4D1/zBq8pWJ0Lj1X1A5v1WQ+zwEFU1noxF1We0FZg4kZlm0B6gTGjvu+4DVQzZ3
3UQoQtMyTSl3r06Z1cwMBT/vkrAqEhCDMDLqW1gyZWmYjAGswt+SngzdvjXFuuU2
FQ4HN04rdSl2z1ruIXIIXRjG8hR31fu04NueiGO13RRlpcWIaqM7iDS+x+zAnUlv
4E0NGyhqYy76GJGBpSBSSBm2Mzv18LnXfqk4v1t6nGETHC9C/02ABtq005ylYjuR
+6+a1fy3szcv2OEb2bRaiBxH8TSmtO2ZM0l9XTC3MjrQ6cmALVbLISQ65IrGmvLv
vXgRtD5cM+HpBc3JCvt7VuCsKaGoiqPxXEYdNJVgj7x4B4VTJNjY95QGaippk95E
2vN2NWY0478t7WT4B5jMUs00ZXlAonoTgkrPkFppfzB69VNY8GUSRcN6F+8pa+aG
t4QoZjvZYXZq7VydGSmkBJcpSJkBEiwHmLPh64L0dzmJQ1Cghg5Zgtc6ouXv8D7H
niTZ0IHJeP0/jIcvLy+t3B1X1eI1o4ZvPdrgnMvadAAx+UzjTkl5nvrBm4JEZzh3
M55fDyPdne32gwfEMm5gfH0iYEEtCUlbeZATMTrns5B+kuTZNuJu34QVouR7bxcZ
03ga3Ygwbm77UKIpiPr2OT8SABkISb4rciMnpAI4SM/n7vf1I1og1BG2hgJVmbHG
+hI2OrtJuztBAbgYbxLF5q+Vn+RC11gAE8aOx/mZiJwKvgHeqLwCrQB4KWq7kCVC
DrM61e/Fmj+TIXdYWYKBpyQvnbNB2RmBFtdJHh6Vf//DmhZDNAXkFe0ccBEwZ7qm
FIpjPJtNGt1X9eYAZsJ+OsoYrgeggN6yVv3a08VOmP0TYXyhWMn17olpJejdfeCU
+GMYxwUdpJdADGBKqE6zypjJHHoVObdcaGTt5nrpJ/2NfP4QFjENvyng8pGMfCdz
9u8VHQ/EZIaq72GwFS+lhEAt4NJKRHdeYH88zK4kA2HCBLGqstVo29xUkJOIfFo8
LQb9bnCQzSfKL/SGJ2Xo9bWH/7+1TeLnrBoGtQyU0+QuYPXhR3kgVKyBQCuvea7G
cGKddjfdIXGYH6Vz5zb7hzQZRbu8XwyFWjhqL3DCXLfOjN3uZ+r5369lZDKr32q8
1DxwSRAMDWhOG5OgYsIZYXYK6qmrsRby+LIUb/1SDxCT8VMaFipQQMDGb8Fq8GbM
Hp1Rkw93xxRRK4giUGGrDhbbKjMN9/2mXu47n3KEGPjlMIgAlNJoGMWA0N8dL9qr
9A5EQaftSHsS6frZd1+RprnQyzMqkuIYJ1t0Dhng7gDAcI6uxzF3OzHnWmHKLM7i
09UN55cudMX57tlsJogg8goFhJoKkPjI2Kfm4V9mH1ALPiB33rKgpmMXtQRlm8z5
JtUcE6wMgrHHf2suxy/ASsenfzieH/+y9550TITNFHE3+JAGKVdiYpYBOKL1Be81
UnbtuWts/BR8P5a/9XtKw4FnnG5ycPBxciabzdF5nSdaXtZxg3IlcOoi3cTxqPcv
ueZz1QJ+Kgw7LIp5h+fLYEUWu9kfvBdJgeSAOWehj1l/AggtiOh1fS3Pf85HmTY7
6S9R11mtth6pY0dhe/llcQiitOw/dvyoAJaJWsdpqpAjBR92x1N2DZ+3cHnXwtnx
Kcc3ViJzo4DhPGAOgnq/NHLmjLzUCo3/oFqq8IkaKdSJgEK+HPtVNW6WKEV1840Q
awK32gt7Y/q63CMjb65JSCDuXt5Rxz72AKAQXO4+ayp/W4mygwzpuuEc7e9FOBaS
HyQ5MWxCmNMHpOT/t4YrZFR/f3kRoGZrgWros0GkpXMzab9InK+/+KmjGj3QdWqM
OK76t3kvBZWndYkUMABcfT4e8eS9Srt1M1VAGZ6Bh8SeOKndzqRjDd1w/+G/oKgS
uOauRGw5UWp5gxp0sQqxsNjmK8ZuDPFCk/vuvgOsgroHx0eRI+/to3OfxgIcmig3
PhZPdSmqccgyG24zVzd0IXVPbgHM8PUY7juPE3SJKan/l2nOWILJSiQAHg6lEHTI
AmDdWPmlsoFDBmbPRk8o96ptXTFCN8ooTPEYUrMJY8dfTfHmvggGOwOufM3ue1ww
Nmm0Zc/1w/HlEBHDQe21mPq850LYmjkTvJeqAybzffWwCSfZ4fKgiQk9LlOh0xfT
DF2dS1P4Sd4IedejPtEGzVYYQl9hy36som8c5bcbtUbsjR8JZSLBboxzJEqH4vbl
ESkb5ju+Daxg9ttkYj6gYYOO6eVGQ1HoZ9yNw+8Mf8TUIfFP2j+IPH7OF7n+NfXZ
FOrj0ctZIG2IV7LAr5G9BlQ6MRMFBQLUC6FO0GhZow8ChAUAoR1uTmgg7vgrnFff
HyyzVANNPc5+Z0CtFTQCmCPgPsVyC9ubflBUdTMeBWqlOTWnztglbSUkqt2Lz+DD
mtVWf/7qzw+BWBljyxijsmYBhftd0W27gqjn6JiXqBCKGWGWoT8aB6lgBE49TC4+
BeDZLuv3dbhFwfVHLmYNPUQkL6swHIgHoL0p+Rsj6ANT3VcGg4PRa7BLL189Cw7j
8bUQpDj4a6PkrncpnV2YjpP5auzPPew3r+DpIjGVAuG51rfpRruXXgiXAG1gnMfU
INSoXe0A7wvkv/EMg5V6jlivMNXXlZcJFxSUbTPaOcvGyv7jaHbGK71dUeFEJw3m
xNw0wORyWSiRNKfaDtC5QNkU1bT5ZZK8ULtpJTwQcP6bkwznuMPOQ8tyw8Ydk7j6
a/9FqTLVx1ik95BF52nBDNBlEit9o/vv/n0vSR/lYULdBdRj6RgTGO03Fl/3mW95
yJvBMuM1b+QKl2dT0qaKGUGGnTguNLNBV7nBINESIM3xyFiPGBHj1kGQf6E/MNQP
6/9AGM04nbNV5SnkC24jQupWiKgahrx1tZ1Wn0V+YL7/t4wrhjmfGfE7cxDCZs+Y
DVjxWAU5AYcxR1SySwNR6Nbubg/BV/53B3rSl02jhUzj+8zdyfMV0pScN9xb4/gE
Asw/UGcc5jNt66poLwcZuumG18TJEXtDsCuQiixM2H3LABCYaLEs1rfv+vlQZkDa
VAiHBQoKJLdAV16jbzGklrRIMIzdsGC9kea99+0NsPSoE8QUBq1MzM4RIt0/sJJQ
AYAEyYEWQCRRy+EOCLuj+vw/5iLu/St59cAzYcnUf591m0TqKx8yfviioDb0KFSS
Rxqd7lf/6vqq99fgnelGJvcI2ztD7RftEVErMVVZ8TAyou6jJ75Sm7K7VC4F6s6h
3xpb53DNRd6ZGA9bqm3x8JSAdjb+SBY2mnw44z3d6MyTHUZGWiUDTnj9jgpjrwvj
rPCutBoXEAydeQrfrCE/48N9w+g10KVmkeEUygu6phEAngDCz7akImvfutm37ryG
DVGjJDKNDqH/Wdsdhcv7rKPs0BBYE1ElnEDrGo+nw6p/YrEB8uCy7jGGL3eYhBf4
pMDrdlXUjBAmUHLkp0eomFyeuOtUXp0AdRf8bGHN4BCeagA95MfXVFh9vW9LcdAN
Tn4Cp1+mtdFaJ+Jr2Ei0P/ikYlVOhoGQJ0XS5PJ5CSNkNleKRY5P0igc0agLWTbf
Du0fmV0t2PponIru0fJRzSi4rH49OKOB9OC2VO/5oPFDS5ewnYvBrLYIzeIkaRn8
BW8sQmlimr2TibUj955iRCWrFlTTiV9wtR5JE5HL44v7zlgNlkxsqTskr5g7ytpE
LQQOJ6tyzKn8kACME2rfLk+ZCurD6qYpP7aRnwMWbxNNWhkspqqtRbUGJCFyAWAo
q2I40BAxuP2tQqx8QT6fWV8MoZEUjsk14y2l8sIe7fiS95n2azzEgUJ6Y2kaeuMl
NixlDkRZgTUAyvzukxPVjJFgPfo9SOxXcQT7gMlWKIaPBYvAnnOllSdDwlmDSU1d
jp/rNyAuh/WCSbi/IoGkPSms3w1E2OgNjdguZ9DeG/FhVDY2qvKuevnd/a+8L7Ix
hatyEFh+cZsJgYOPP54sEjIe7BSYaNPzG8UUQWTiSwPz3BK2mPwlPwbLbvmLPJip
HlGhIlUvcYi7Ht7zbHfRP5T+wQbJj0u/rinByu6Sss0tTbTXfGNo3UZxa/6vZRKT
QauYAYP467bRomFkYzcXpMHXaw5HARTsTfjUqHGIx62Tpyc/pdUXR52AMWGt0smY
qeh6UD6HtkBNr8xcoDd92uMgq9sCqvc2L7jj46X9P6WIIlMr9fb4tW7zLGSKVG9a
KO30yhhyJqLwo55Udcs5dhto8ORGu76TWNqWXw4YodfzNktqbd50ZPNn8hCW68vW
fWW3ujgsB21tXul0nj0iic8GeuK0yen/Z2/cZmBZe6BLLJJ+klwnxUXP8mnPRknS
AmHihMrBqxN78mxHZLJdPO2UHVjykDxCRZygg4a7cmbX0VIJoVrSl0rY/2r3DhpC
Ea+97BfFzDHrvC4SA7mc+rANP+PMHZHyS4gLt8+h1TobliDqY4/1tfHCGak9TYoz
Hw/l6zAMxyIJNgpjN+8g5HhkS2+REY9uBAUtDWZx4QlYPkJgX/RG2w9OhNvImQ5W
bdzqqXXJFzuAN+JozqLa8szZqAXAW9jP3cHCJ4PVq05tV4VpEFSKi3XKfPfqBwrk
Rm65q9p2+cKvhgCQ+PFMbNaQkfHg9wRwl1pgGkYx//Hi3mp5ySnD+lICjgCPqoM5
33U4OyuMRbd6bSROXZVyHol7us1VvRJt4vPcnuIv9zQqwERaoyAnkU0BGD3SPu/G
7jOQnbLXI4oetJmwWzM2XcmWun5g/yRO2MiwbmbfGgcbfZwFIzPIT1S6X6GhJNBr
ONmezVzQMGqh6pvWOEBOPAymMvWxDbCvDkPHoOKszuQC5V4ycbg+Nqjd0h4kX43d
QiPDMAOI8kAlRSZbPI2x3Ci/UVY+wQkSiv/fUkg6UKrbT+ixul16aNOoUQ2MOOk4
RxX+cxaXzVKjGAaYkELhBCl4m3gGPsTyzTsYY1ZVK7rQGU0cZyTqRG43glbniCQt
AXws+F/VrGxTQPOTyePpeKQHbBY7uJ6LnQtjYCuG5OQEhuUZCs6FUFjqAfwiCqWV
7WSvJfeEDqu/B91TEWVDtPd1PmoBbFK2+TJNkffyyjaaMl/lOTOuIZZe08T3B0Jc
VhzLeQnhzyGE0h54jLW67AQpN7JkU4V2hU5cY45ekITmFffxCn2JNzQX0lIbDtrc
/cbucY23Q6C5s7x9Fon1OncbKlHPT41DQJ510UFJ76bZ/yiOH5cxOQBkRb9nk71X
S+R9j45489PO9gBBBpYvd7uw63FhI5c7KVJ3NJokdyRWoglyLZSTcGCjuux6W7gf
xMTwZnaoJ4AIhL6aCNyRCZHsf6OFp2HkY7L1oFzCjEyj4lTT5xJOpWQAMi253fzQ
9KoizPRzIVae0Q8nf0xKkl5i9aKYrJICH9pKG6SfPtrLNZxPDdelmhxXRv5I3WuT
aMbXuGGMrg0IruM6xrnEkcC1UuToqcyG4Dw8IRANsPsOgBu2cscXvVeBYf2ek9hq
3xCRbsfIirxEHoG3xvkwDiGj7qpx7LAePIv5FZlyu1tOorVfC72ATMow3XhfsQzx
tngCz7JqFbQI+rUijDWnfobUTwlYrZmr+1GZum/SaFp8DsRo5YF6YWREVRkijs4F
e6Sto05KkGzhm76VRlMNOLiGfl1GK3tf3VJ9c2gXhEQ7+fCxYy5ecTm9e1qCosTH
ViBG5h60lNkhaiHw1N/k3hVCR8kVS1MxRgn4EWzcFzhvc9FkMaKBGYjx23TK63LL
t9+3o15RmTdI9l50oipNRYK8dDhNchOMo5+r0eloQVfqW7KiWyV+cykLUnbGRHwS
ltUawEq4qBKtdUXruUnnZJk5gqHuRr1ViUR+pg3NXB14nctJmWDDdCC0M4QsZTGb
9bIXJ9I4WJGVPYQAoFBGCDB6LfACqPy0Aext88hK6DvCa84dcZy6hninu4o/cu0E
G946aON53iOua0M55yXeoiv4xmJl7jJR+K+jfUFDf5CayA6NBldaE3fgj/NhK6RA
jDIhWmRzbkvHJ9eO92+uG6p+GFs3EN7Ny+PsQzfMhHRCjFjsjDjDmXyRIUauVBh/
pU2+ur28vA7U9DwcNhZVPsgM9a3FqkWZkd3Jas9lAVYVDflClSEMYSI/fe19nrNv
VjNvwNNZ0ID5d2EMfN2bW7a/TNEW+US3BJLbRs3UTNZ+tInotVC8+U3hbKlXtl58
0eDfju/wwfdWK9rKy0Uz7fUajuEs51QTQ6/r9FCmLYkfE3QHLY/AU61auZsGbC/o
Fc3bc3il+qJc6E89aX9xKpLK4GS/b8BMdSag18RXLNNTNCHXJFVMP5DmZX3Xy9xW
zepiE3TGPNRhoTwD97Cwkl90hlcPLiuuzleQj7FCLnqp/oZ2G6MyAxLaVtuV1RTk
D5lmHnz3QoaTlHIx9c0BgcOADTxvIWDV22DHCRUDYmp5QRPiM2GioLlEwNAnfAFx
rDV0BsJPh6NkGTJ7/ljP/5d9dZI2GanfZJaWOXDBEwRyMhS3d5JFQ7PSkj4iMKvF
oN7qL46r6Nfrkg5X9FOQveRxu8IECiazlat3I5olKfwB4wdi+d5IQQ8sDaNendxx
pDSMWGo+B/B+LDiAQLUuQ35z+kvEHcHwPx2fAWkYPaQpaL5L1FSdsw71RhQN/Yqp
+wpGuTpKeL6BubTBOHdr2DhesPXqzmytza1yGjEW3N+xhHoleEDscJ2vJysVqpWF
7YYluHsZJjrAUIZxcgm2hOxke8bUcOCQ4x/j8KRSQigeITHjD4dJ8DwUkHvK7ipa
bkJ5aZ9oD7puiQrgZqk0UwA223b3EMvH5+BY4sUf5Diqx8RrgNaRg2AkKmwCHrq+
L2aFIXtXXikAA4tSu+eTSpw5muW8CEg7L7YoEKQK5TZhK2sXY179L3DQ0l6HwKt/
qDCrB7acr4FQYoAAhZ0jBH/8Mlg98robhxvAkYHy2sd713mp9Dl/2mxguM+XJBsl
jYWPtNWxYFPA/xAxwUH/8Y+ajZy+OMA6Pq+heYreV2smhhw2KSk+bGUyPEwEQFKK
+4xEdlnesRRICBMOWTl39gRuEewTcJMTu2SijlJj5vgAuZblO/Yub7cQX9Eqgrwy
4diEk/VPfp+ZCS1LtomgSll1rJdmbPAoU54+P9V79xTH71blgYE6csF5RjL0oCmr
YuM03wC16WFze6PX1i0e3ENMippi54fjOM0wfNTsCn5wh3Kl/ubSQDGlqWK3P7z4
Xw3UF2pkdNZYWmeTVkHqZK+voCPmxDix7/LRTEqs73A61FN8iuCHPWSjVdMbmQXO
aBh5gk7tmaeswh1Nlw7OnrKRu2iu4RiiKukxlWjq2eEEtCxXyVvOCGdHP2XK1MIN
gA9z+kyOMqr++8Wk1EEISdrIxiRLNQh+WegG5c2tLJqjGw//3rw+ZWg8s1nWS+5I
p5d9raAZZGclfcVG/FWm7zpiUyNQcDLWrQtcbVZxonx/jsQ+DZBuiXy2nqNQd18r
UidpFKXVE3QzDV/h2WNVMp6sKQ7SEG2lqwe7Z8mDBsov9x37VXjW+XRRGMtknlH0
jBLQM9Fz1vjeDTD6LbqpAiekemZXTR5a9QEOD7nqgQ14WJ9Kxt3VJQiyeen+kkim
0FawaapDJTzoYMXFBifyDVSN7ilOpzrvAxlyzR8N7s3tmupD30LDTayyG+osP8mw
G2yO6K+51fqrSek/Y+qjNUnTVMsBFYgdpEOslqqj6FAMwMRJmMp5WSJun8ukhnR0
IaREJodhM9wlcnrQxE6Q9zEL023dlIUS3dsJ+764qwSsp6Gz41n+qADaOpXYbBlJ
0nsxJxCzIdI2NcksGTnD2Mcc+ssVuwZXzX36AN8cT7Sl6sTfB3YcmRJTz+NgB6M+
Ye0tfAh+loLHGSuBbYUK8W0/dciH0lJ3W8+BczAMijczbHScxsMQ52eluvPfEO8V
nZGobJeArZ/Vs2jUSpsZJkWVteUKTBaIGVN2yUD6fofg3LJieNyf0ZMb0euAMret
AM0R4x+fhUqVKLpvcZP4rbljafuF2/7YGP5szv8vTcep2C8A9CTqnpIAVFWipbCF
RKvhZz9D2JPPGawEIvkuNdGvxCFTSNh4pQrAjJapND3y9HnHdNPIBYTd/P9BFutT
7d/2YC+Y9xtbyWUp+LLJ0OI7JxNp6H97r0JsKm5f4v2xV69KOYjFjCm6kOp1xkrm
cYO+D0wiLpC/4D2FQcXVANug6frhmq/Innd1vLcAq9g8SRNrTQJgbLP6TZ7i99gm
WG1OiIpJHFRMN/QIUyr96/Af0XM8V7xceF1QDJJuzutycvG+36C4NjWDBRA9Dbtk
Zq7gS2BaJxeUXTcfSR6LAIAhIne+T8AI4iGCtGu+kFL9JPHfXZFYllgFkS2ieeJe
aIfMxPgKaVsCFtQlRtq9Vhflj4AJYbFpmtFqxHhJ+qXh06GTi8L+ZQwjPTWm34Kq
rGZZdfGjwyjQ+UH6UmfQ7dHcILK3xnVSpcuClmuKIhWXRE8h6tjMkYkmPKGQocz2
o+WAu0rk+e9RBiN05ho0oEwjQUWas2NFBOR0SYtkQq85nhEJ59tcgX88MEdyPDPZ
Gw9mAQ/Pn383uIxiS8CMHGDg+CA1NG97KTVPgY03XlxgfW4sZahoIqTwtHzIc6Gm
595Dr3/PVZJ1P3GfVrM7HiyKmWgeBv8KvZyMYgcqA/ZExqaR2u6ZDCVZdp+KHrXm
/IDfZBaiDKx2kMPUIvuij3v3wgPGoGPF3Nekpiwi92ud1JByfP+g15rtSJBMne4u
r3N4nbgM9ERETTldCwp24nRcA6rp+AclkCEvjOoBl/1t/4lnnop6Koe80k9rl+K/
u1wX+mXuI8oyP0HxloyEBojV7syyfH6TVmrmn0pn73ouwvo7PleoFvEOBK7mRVEc
KVBc+guwK0Y1e4/iTZl0d1M5XsWWmD4HxQP7/qfiZBfQ11fbf28ya6G43jE/BAjX
GLcsRyCOZqmQw/iiwu90W0zY39vCwkjo0e9Oag8DuSPqKvBhmSa3nezNTlyNFNK1
lVx3iqJXsEoJSaG7pishcmE0S9Q4N2iZzMJ+OYL3zASFcvU/sPMuRDS1Yij5c/t+
A6xAmeyEeqjaJpJQBG6RwPD6If5+wGfIRUh9eHSf/ppCXFTjowVyLA5TCR7tVFWc
61/dM0oY+bjmNlzSUk3jAeNi0+Y5Qc5lDVLlcBGigQ8yWwKO7KQTk35MvuRhnZaJ
XKwIUMECmshvmVz5Z3ckpGjumZkoprQyK8ErndMfiIYOmrKYnbbXqgk635Lk9Wjr
8LKylPOLX/s0aXVOyshktR0hZ2zUtFwr85dmCkGs3P4HO8yDDMA5ICWCc7Ok4EjA
R9gYKAwtQkeDZm3CNdcH/JtNecTPo68AkLDB+WPf0PkPegd0+VOaGz7BfQEoCJce
pk/YZ9gpwZLQfLNr79ByznRjPE+Jr0ZV3Z0kl9UwdBXQh61FrYUl2gDRgCo1bkmy
VGoPN48OZyN0MUqng1LMW0wpAyzhfIft60G/8G+weCZRs038Ka7uhokhpC24YJnR
sPj9UJ+kBab8vI8brZ/mcmqbLEsR7s6oAKeTbKOmtlf2o9UCoKy0kj66jWD8fnFJ
yaOisRIIy0sYQWNQCudOplO8/ZsmEjmFNWQ5G7jscMvd3pVzHOvweMDV/1BFblCG
bOm4dsIyp5M9ABTUm/VxYeduFI4TIfNs+OUTTdqc2s5/I1vgM6vnLEkPoYxkU9Pb
pXfFvhfZediwU9s9ko+PnBpAoaLgTh9dfCeh+oVYJgnyMfhoyXpcKIg3vDgkuRt4
8Xjmfh5gAGYgonJ3AN1bADaew72mY2q+FhzA9SzUmGFOhuFjhsP4YFHUvtqnW49b
1G6Tow7MJ0lvXMD5rTUw2idqBsW5AxfpMG82Oq5YqHLCDlQechm2tkBwhtYKDt0l
0Ggh2T/bSVzc9I+HPsCaRc8qyxe7z+vi+BPVKqMmiMpNPhvEVRytt6oGRAdBdflN
ZR4GaiOjMPP/IuJn/vFOOYsfdvVHl1UHQRfRIjYfeZA3MnJ6/HsZNppIeDBpQsTe
D2DaV2n0vMIJxpB2TyD8sCyYtRf9AC1s+65MJXvn49JqNWz54XNjGxhxphwIAURY
zQ2ecf5hNujbDQNCCDuOq9rGgE0BxZdQekEv3MsLUivC3zZvobbg9wq6kGHx+xS8
8dSwFVGKBnZ/1S2Wie6X+hxqcUhj5kYeOsU5GipZBX4WnpOlFj/LWy234EMqUzQS
Q6kj0qggWCemQtpXNWv8o/WlIiVn0SIHuKZoGDuccx63Wg0IPaH9gF7ps3O4N6M1
K3eBG2x9UstvYwJGBEm+o1U/6oAt4G87GdI081ifcKtjWTa+GeLG55h23J1pvxV1
ytEW2HKD42grkdL9jpYAyPTfcyr2hESyhNTS7OwGzOkqPXqQhyWFKefaE2QUwK+2
NS7UPFHmX4OqAfz0BNMiNT8O9ddy+bSQuwIUuswf00qqrLTyDxLmaLNOp1vNAUv7
XuLBSAjhXC4pThCZw5dXEKTAFXJ1XSqrRchuOuFSV0PRBmlpAfeAdJ9AxeME1a+8
IYvJFjiF1JVlbbIShAiPdhNv/037ZZ2o1QT8hzBOj69zItR9UmlM9S80sGPWnQJn
KijEc2TC4EDq5l2j8Fup9bJvC/ExJVyitrXyW4McOrZhV1o5xMWmZpWY0EuFF34V
ITDuH/p0TCG29bbkegmIF/LjMlB9MSJImUCnEz3HPvGRhac0BZ7FSCdpzgBaMWQk
KzP5PcORSkDg8y9UXJNuNvJbhbXMxXcFBnp22IGpdxC54hQ2LlhgQtgANseT87Jn
zFpzXsCx8PDeZO8Pp3hD7aF8tA/B1WPcGk2wR+39ap1tolky5qn/DVQfRMuXAtbg
1EQId8XXQOZESP8RbuBbsbiXo6leuCCJ2PdhtMVfJ475/NnYS6YxBeudNcjZClXB
x5rWYbg4kcaqg7d+6I7kLMh9puziIPK+du2h2AXaGY/0+zFHmQ0T4PayaABQSTDz
1zWdNrIO0FO6bg7x2TWx/ePBVDVRDVvSF0ZT1o9zDYIh0sM7vkmoUSYH4nO4cBEY
ZtzmqaIETpaEMam+W5HkB6t/xWqNuYDu8YHPzJXgrNb+WjZi+QwR83z6Hpj7gIBu
GbClhKpmxMZJ2btoI7K0IUyCMSx2kNOzsEHPVrHThFKEL+Fkc8LoajljeTjqRjmR
cqs9DF08usu5mRuJRjx5oqGsSweFO2w/xi8n0/7Wq6iMfJRDruArKa0QsJYpXBCJ
4foUcNnarpqwHDD+dqws1K0Undfe76oOdBdcSKtLgWfPWY2H2sV5k2bLu5EY0/qY
gY0wq5dQbe8lh6XCKw53sK7oMtbH/UdH9d74B2u90NtmoGZ49JnJzYkVlUAA5CPH
zkEn5PfmWN33gmR+I1ftzHRGznuUlWHlMT51+zpoiIuoZz00D9uATrEgBWD62g7n
G3LAHd+/AQI6VAIiMsNGGX8+m1OkBjl22pK22CsQmYWoCTionMUMixMlLnwxWvII
wc50FF/v7O/fSiMnnLYJfxtCKmeXO3WGIizwu4IixBqkdwh3Zm7Nd6Qb1rPfAUzC
mp6sB+T1KtcIdun6c3hkMOrA6m3sEHvrjsakRnb7uUzkVdzrVVxMQH2WkJCGbm4E
5KTeL1NEmWdWrccxkJ1DNk3NOvX28pQ3NaftdGnxgfa8OAXT3zQk/XaKEPKZ32qW
AYdkLW3ZDwLEpyXQaLFWbxrCsvo0t3FuUL2vXBrmpinranPNSYwuKTK11KhDn6PP
bsKIlMx9R8JZsZkocMBlTcK8GilHwbRImFt2eL3j+cYevY/WCLOToB2jgyk82IlI
rvZcIsOlkg0zr5n7uvdkZ/n5ZBAXtxDKyJDlwjUGI+5yPs+SyuMzlaeFxS0H1bem
FJwNwiooKK/TCANNDGniK918a9MkUjHlXDxQoxfmN6OzV7wTH+5pYKXziWg89qAg
ca6DqIIIGOLpVWIgSJzfEVIN1s51jIscbrUBbMzQFBjfKFrx9ZCTvJhrFTJCvMd1
ZPFzGKa7XtrW9Rd7YsZVC8XNyBmkUUjMFsu0ZJL9LJ+R7PgM1cSCBrwDxPScPaY7
ikXi5w8Wx3+KU2tDXr41C4qQPa68c6NP/O1m6trhuLapFTleZ6uT3EHtdSeo5o9k
n7Tf6vGob9ke76L/ffoRItG/bz1o7l18iW5hErJ10fPRrT+zjDZ9CGCoHGp7YI87
xaTQcFTaNa0VEOh6O9dMZtvgDoBhkTBujMArtiYVnsetdKuSL7sVcIMi6t6Rjp9p
BG3FZBKb05QGFYCfysmciV7FnuWACJTeObuYM+qlxUNt2s4a/5y3XzYXhgunlhu8
31iy1xcg5XgNQnLEI9GQ5plVFWxKl8xg/8U672TyXODQGxi81s37N0p3DNVntssk
mxvCxmvFMj9dRdxkJcbyAfC6Kx77ihciu2MNsMQRyytxIsvUoM5A7NU5KNPvpAaE
RiDqe/MDY7+QMCVXxwF9+xiWHLEjgT0Sv9F+huECHjUfJEdtBTzSzLopj16djgEQ
LdPGq9PoZBc5LpXp/xwWv2OweOdi62W5MaJw/01Py2HqK7vu9izxV+0d/A6urlES
2SpQtC5xK6hhuPibarmnNr/43MXdxqa3JOTlTGM/hukZpWynkOMh4PYRzS+v3919
Cj53NfOTxSEG7d+WDRuVOTDUs+dNXXpcD742x9n8jf25sMGu8QJ6V0jUn9VcRDMz
Z9LNzo+hsbA+XNhK8Z0hA8YqH89iO52/jVyZeivxEpndRhr+gfmLeu8vHKbIPxsO
3ochidpTGqTQXEVfeYVWkY8+Q9XWT8bIWasdqjUBwWTvo9y3/0Tg+2In1hXATkVW
VcOOaa0oqAKonNqmRR1rgc4sCVxc17T0Z7OtZ2dOoMQDvw0JfXQaXeM2vAhRbsN/
24sBsrDWzC2zLpUv0H/cnD9V80M9mf+DQvzyJBKFXdTyKkA8VtJd6IzuhR6VYh+l
TbuSxDLgnmDBuTLylCodRvZYGwGpy8PubDD6aLrt+5B5kLJh18Qk+zf4O/HGjx+F
IW/H/TEVzqJLfrmicWAtrQrSxIcvy1LsIIYnbcUN0iTpnqHrvpLzLZ6ZrNpwRx0w
TOCoiUGpsBCXXYU+QAIO7+RNY8TChRosljdbxSX058XMOLXgr5YG8wVDg9c/uTpP
7Sxp/4v4zG+4h346mPzsc/kGwsOOfZkbK06PTQ2Oz2WkPnbsWqPy4SJuj3TOwkrn
/IGRWZk1wfoKn8fsPkATZLAcxIDqcj6O1eFjeNBp6MPg9LniYubUJYLz8Xt3WpvO
leNKQ51Y6Ue1P+pYRpSkSQIIZCWy4GguLrJWMMfs0qoZ8R4U4IHfX46jxSg4KU2B
CX7LGpOLvknZCs/mNd3MoI/2I1/rhLFIcSRiETBcM+TrmAMkEdJRvDqqJO1zLQpF
S/XB3v1DXWx4FkLI2VYUH30ILGtwQWOEJa89ISW41QMsb6vMWt0DDCFQ+pskwEc4
mX8QX9Qs2trZnGiOv3sO6AdWWmIzajuZKJ0dkILOapX+I3AJ1hawNKiPKJ0K9mBh
w4E4vsAXNMPlBeYdQHgEtcQm4XRAswmiIeUTOa1vVMl8K/7pcyCk4uu4Wm0+mdcT
/RpGDOYB+v4R2mgNZP26Zhs3PVWnTk1bZ1v/S/FEjCDZjbJ6OLJo7J9juzwYdIIt
vzr2ScdRegc45LenDD5rstJxlYJiwNJ8jtIVrTp+NqPt1jx/oG/Gs/sxBOQW/mQO
S3H2eidyxn6yZbnKTf86mxBnIMOMLFr7c/nnxjyIOEnvehMLnu6QEocwIRWD83f+
kcIAtKBhvRkj47cn+uIpVPvB2iUXmddyn2cgaoZ5yWpbSHNqKYeOgfhjPZ+8Btsy
0qJV8dyutfQBAUE/36jv7YcfYk82ZI9gE/OeDzml3pJpAI41HqX1E1/OTeFcotnQ
Xx+627qF9hNH0rxTe1RNVSrFq/UYIfyfdzKNM0XtIi2uew1Szcq+pjWJJWHSCru/
1gDLvkZ6N9HODI/PYJUAsJYBRQWH045mDS4yPpR9NJZJKeW/We5v8uVxbeARrkUE
QB03apkhEntIoq798u5gQnLCkcbyqNEfRnuUoxIUMXe+OGUyAUyBzBoh5aJHxtW7
o14DsyHJ3Ng6s1YEQsXnlmEauPBnT6zQH0rpZScbw5FdTd4Q8RKfhvk28QwYLzxJ
NwQeeysvsg5qd4xkCVueE9NGmeR40TxLVz0GyV8Lxmev72VQTGWJlneLQ09zja7o
FwiHg2QUqopgAn2Dm7xtQ6JjXIYUenJhPTowq8Wlicfjeyj6bQ5oClnKBLkvLZ2Y
rBnO+ajAWPHrgJwlaHolYPf5+PY9igXgTDctvNPsJLALxvOnwidrzkfG4Ffae6ql
p4yG1A3R0wtIAAxaj0ZRyiaKlRfdLFLLbbdZNVU8kg+yohVIqmXieGHqRdOwAdpn
c6J4/4STl958gDzSVBLeDYwWyh3CS+9SwiZH1VVP+3F4o5a797mgLLny9mhfVssG
yO1c+zcMQTNKEmdk6hP4qxCJH4TLWOSN+YdS/ko60qlZTrqzZb5BhGLcADKy/gww
b7F/rdlRB0SIj6XlZeMrnBGVTfWItEFtgsGntedH16DJk/8jnvgE/DgCfpmvvkbK
Tp3JW6DlYRlv3uQB/GCP7auHX2Yk5a0O6Di+bmQiBzxyuCJ597PrYa0y+SezPOI5
1J6tA+C1c+RViC0reIEZz9VYGBs43x7IR9CzrqDjFsh+JQaKJx47bUM3fVlD2D9v
PcrSVIbDAvVJM2wuLjKMJEAT88Ixk5x+kG38V4LUCW/VLtGjpEW9Xqaye18M1EDQ
kw5a/xhNSlJneFWnXezN6wghhHxv20FUL9UvpJV3RQX5hAxQxTUVJd6aj3UA85wF
yHiCh6ID1pnIzQeWnvlWa2NyEoDPLauDVXtd3wrjjrLlRKi7kV2AE4zs85s0Tuz+
R8aJKdnItARKKCx8kRD4yrDf0krGHLvCpMevAGmcBf9nvZQ6/1b0qatD6POdEOcr
uEEOSX0a5r2ceHHSg6a40bRDsrEL2RkQTrucbKTUf28jGAt7e2u9KbfuOUZ8BmjO
x/SCM8Qua8HyWTPl6CIo1HiBS5boE7WkI99MY7sdXsxXVsgVs9SODxtDxy24z+3r
+WxeEZpZSyaUjw56C6ql5SVbQvg+eVHhdbYW7lWZ5ApmO9Bp6Sbla1uuxsmJi6Ns
8p3awRBIhhKDNvUuX/i6/7zKBRohiFI9/9FdNblaGau92LkPNTN3GmMi8xNq96AV
5Z4tQv3tT5F0QT6i7FfNjN1Gli3MD8wcK5KYN7zboXAbzHAY6aB84EjFnMd3C8UR
/28XqoP1h8BcF4PfJmxs7vY3SUuVBUHPo+8pbkwt286z11M7vDI7/B9eSnKCeH97
lFRfaLe4v+ocdc/imXfZGKhuUKxPagdXQ4AZif42W4KySmrBUaE0zzvKgaFxfHfI
K40J1yw7A1i8x2ziYSgmI0FDh+tzUcz7zKf4qLN0jHqXMpkkmgInlfCW4QbuaXjU
3JK5I8GM3wyMxTaHBRqEsKjjI8GEnZhQeww+9JRRPan6eFr88CDM8YAduGYUOIsH
6733OpxfP8T83UQpR/cct4QCoieMAbp5a3BNWbtFe6KPdo3KHXAXV5PB/bA+/vVH
ZQXjFabWx0Hd+f/ni3nDf6ngV6NhAJU9bm2ajCYPnE3xRnHurR1uIPMz4B1KF9+M
KBl8OUqE2dWGGi+5AlxqvxJu01m9/KnQ7+smGeSMW6FQfcCfn7og8Bg5TDPS7YOt
65m/cVYz6LlTj0uUNyu2LNL0Q7ncI2wKE0TYBXPlLxlFjkTorIIhzTnhEPNJtIWi
v6PFIzeoX6UILdPrCZg7AghQ91F0JM+3ju5S4PCR5qmSLiUIZuw4gyCDdKzJ/sgb
uOQ/2O8d+MaaoV0dOJV3/dmjTXcBo6CSHRIQwEiKwMBmIhCvly/3hvJ8DzpA+rFm
yuIGQaZg4jfj4GrkbuVA6hymEYUUCJODaN/xfPzFZsEP1Tw0Qw0dMhiRbq/Z6dig
c25xvGJlrRyI+f2HdSa++iySGAZGlGb1bkxOlKC2Ivpz/sKo3WP6j+ceR4QfMhPJ
+LRXT2Jc+kAbygMZ+lHEMepHExrF4RJevO6KR2BCRRsYhGTUUIIAfOmhFDQ6Z9VE
pJMvFsPXWXCPj3iwiBwnLobHLBP/54iwi1Bl4/zZtJqS57OjStX5zEsUYTI+0EuR
2fan8jsfPpYXWnQyOUyH/s1WQwfOc70YXyTxQNrDu1NOtkgs8C/MvkrpR8z1GcyM
D6p7Eq2p7GIho6zkvY86DH0Kl8p2LQQTMXSLDOCQm1UCHhy/Q9JD9cSB7PzRcA76
W1W6TubTgw8wE4zFU2NLiJ1qRQyRz/C6u8d5tRE+MWt6n1kpR6uXpL4/vxYHZCHK
qkYacwzf0uILBooYyZ897so16XG2zQUG0Qi1Tl9m99mpIRA4jIEtFaiWA2F9eKeS
2Vh7PVgsoeAuOrIYZ0RJ56GuNLOkOL+nHFNQQO2L+PhkYnRv2So/UcHxH+1l//EO
hnyrWnGfe6Y3OvdRTr7D2yu3V+4qqQhhtW7cgayFmhT66CP+59M3EIUQxK2Fm0kC
xpUQdmE4BLLUL1D8y8oQLmApisx4ScQzIHn6stCd3Um/Oz83oT8B53/kcnjvbkQI
jpO/33HG/L7u5HQRx3Lhxmbg2ugeJFlSnh3jMrQTS5AhHrYmfu+sutSTK7CmLBWD
XqB8NSA25NtJO8TEKIevQ27s9PNHHPaiMRxPjc3uHr4KvSNdVuXCnc/KGJUVtKRm
Puw5onJf1Dh+F6+zXXdRjGKp6bFbVvh38vbEuQSRX6Y58S5GUFUvZSxgTO/kK1Hj
q7ZqkocBdbgH35JiOm67x2JBxV0g42aNqN/vLapQQum7O4Un3gKwPzx1fp9Z9pbR
TdsrKAv7YJtWSzRq2EuHuZf59YDYMtXv8hMxDn/2HXubIaDWTm0uRdkCzqNqz+Ez
CVssYiezN8Yj5zJA0kpg03dLmAp3OWOjHnX299lqQgmWvNSIa93HSGxw0Qs1QUi8
VRPmjK+/NWQEKcRoECezrtWOy533xVnt3d7FYAm7hLE6NNUY8DCeWB0ktD3UCqbe
5ugQNOWcQD/MvEArXlK74zqjJ1YSWursGO+xg9hbfxPZ3zRadDTB/4SJk69orChB
7VstHXS/U3nNWEL9fBOFkZAVsD+Twe1oJPEnWTk2k1g7z72j+7iha0FqQmU2gS0B
8mis1zW7J8ofSd9niSonFwnV4ZS6E+GuqsaXsG7JW323y9HAd8SXlzySJW7e+Xvt
estx6NA8+e2eUk3DIupBlASWg5kPJmdRhu7ybTanfP7s6ATW7JUVt+xUVcxoHPe9
/2BAFWWI4hvOCOU7iTcsVQ98V5VChT5a//RPxfbmbpOne0PbegVmWAzUsxYRABpw
E6xnPcYUNpmYaT7DnE6ZJmfHUQ0mxm1AQkfl3hu5flqyhRR7jCP0wOy3RnGmsHK6
P0d25AJHXpAD4Z6bcOdpxFJ8vsBCyDhtBNPcBaPmnqclBf8UrKybCusm8sszy856
EY7RWQKlkry+9sUOk0Tb5zjYuV6TSgbvQkVn9Lu7pj9J3LivoK8+8EOWCTYcFSC+
Q/LzsLPhVWSXAoRCnJyL4pgMay+tzDPGq/MguaPsLq5RiCpvqUUANUOdzwIuWncd
afFxXC+dAxn1tlZLwOywJrx7t82a8V5c601fOV0FXkUAp9ag2p4rWoHB5BwCRfFY
WqTQR5loJMbGw0nExgWc4Mq3kY39vITjYncclOBBgYBFYiAR/+Pn5QNNJQiouhcI
OjfCm53zeFVS99JSRy017Uj5DahZo/FKCif/TsA4Fmf/2SFlgGNehXjDNjRfLgwF
nStO16Zff4DRJ7SFmUahsiIEqMeMVe5YWw01xKquX9ZTR0tyJt4jiFvvLoAudl/e
rHMudbOOOS5sXEmgWWJ4Klfl6ajK84wE2P1p5CDywjIzYAasRqfM4+vtT44RJaHb
qYoh7V9TJA2vXNZSvBQg+Y+UZtNhczch6+1/dD8C+ulZYTXLz1WLhMGGQAWYXz/n
KPghz0JvNZfTg/7nj+pfdvl0HgmIIWPBYJnZQex1JaOYyWRGRZ5eF1eKQGA8Gplr
LGSlMLT/EbGd1hs/TdNodRU+5zOy/08u9cVQ/nni6nyc/SC5ykPa7z86nLGD6jhx
oWFcITwUgnV75V+noEJnl3CqtAhb9yTs62qXdIsFbufrRJN412eclI6yB/8AzxK3
MyKqIaFvGIEV0Tr6U8XNjM+p9+nOM/9ER2VvfTtSS7cH4URi4YLESRIyWhOnuVlW
GWPIhupeLOD30q1lU2zWyrGhRIz/hZZRw2fZTo8tD9fgQ7hmpLUaZn+JohqcyJlX
B/u3P4zyusTLyHBtuy8nB8VkCwNawnoKICQqc1JRvG6poNbcjTwL+87Xfmxot3Gv
WinYoVnpWSkU0VRSPn+ROqPJa8P5exLShkWtQH5l7ccBjXPyF69jsaLvECSQo3Wr
A9umqfNInxyVHUr8h8PCP1SeL+CWp86Stt/kXZTaCmRmSNW0eijAoxUf5FWp9Xvw
hXJgfovjwgk3ydRlzSuDHJlKc4fGnw5T7gmKg+KAJXlpyNXYn2Z3wGQFFQqEZw6m
9oO1hxYJD8pzQNl2+7Ia7+jyToEdJPpGOw9656c5u55OOZTEF/QrB/6cjGy8AdE+
4J7Xo+BgCG6DTpqn4CxqqyQkNEtOUokHnJwtsw86YA7WFAHXBiSQ5BJi/0HgjyCy
garoweXVDaOVeyKvUMfRp9blsDqczAZazZ9/figpFMZKZgpa2JvqLeP9m7C97+pN
ewfrV4vTYZVWQQRQJkJOJAFZtJDZjxc6ueGL964gW1YyNxIHEfY6i08mwMMD/2VD
6+FKCkUddinWUIy5eDQ3OF+Pu6J0shFzeT7MP7J/oDYbpZZQ4eikeAKvbE5x5434
HjKIT/Wt0kr1Tg0GWEJRovbgdGMZfc/r5LEayepromjunyf0i9dZcsjo6JrSUQNi
OxrVaT+p5F8GL91f3CBJev/9ZFsDYJff6trzTta2SCCTvZhawzREHnobcixOgK+T
E5d5yHcm5atIVxKQrYlT2Z8rAjVYfBvbK1T8qb00T1U/2V6h0Zne/lQDKMKCgKzL
laNvPHNzU2NYKmU9U17YFfR/qgh7njxxWDobWuWB6o6l4CMxL5aXbbDBpeTNo1tC
E1jloxRBZr4eThxRL5GDUNQT+XXOXVXNa9uH2tFQbVY/F/h1C0tCTuek7CqzBeRr
m8Qy8mppU1ho2AD/zyZkZgfcQr+hLhl6tVPhC2Zn7ZGHoncwq0CQIbCzLaDabLJT
RhRqO9xUzqsMdd9dIUrgEpIk/6/U4JkWrD9iwkXAVn2cHD/XQ4aRXONp5ISKMyGe
kTL0n5SGdmpaBrimBFI+Z5tBmKNfbB7iP2Rg7mTP3owJkE7fn7ID8jrLa7sUa1mB
Kvc/krwuvttdJXREwGOQt35gbA9SuS6q7y0KbiawJl419n7e6QYJUrX0Bi1tzWRO
jvbB7tLYfRlU/yh7YNe+hSr7B7nWn6gOVX/fRcfl+fREORZpm+Q7Q2ImMizB4xBb
riueu8Mj1VDfu4MPZsA/cKWH8iKeEA+FrdykkZsg2+FIw/20b3BvZzaN7OHeBzdv
p9VwMF1ehFEedHLmxLY2NAjvSnG2wuVUVUF5uKhu+HcoPdQE26i0+vFCNUBPiRIQ
mxxKZnTNQCCKElBLASyKnbweG/BeZl5P75d6XAjQkfygKZY5Edeav/G0ruiF6MTU
ZGvkswTbGz+hVHkesH+HlHshfQc5YCBhQoCgQgoYdSNC5MFYuVwbNWvl7s4QBbVM
0DUXf3KiVKsTmJ0IL2x/wyfCtF9K5MfwdmUoJApDF5SCGL0xQmkrTWgVQYkS8DPg
ojF8PONH5FwMB5qlEouUXRwtYGTv1t0FUmLDymnXCIQjxskHPuL6btGpBIL0gbte
uaPRemqAp2fchxY+Y0WSqOY64qBHLDX8B7q0tVdyS02pHaBc2z7fogQvUFJtkKm+
q7lOe39R0DvexkcGTN3CrFJxRwt8njHKvuY51LBKBPqbUNYGy8Ky0CSdW1mbyrff
t6MgDgSLAfQslb/3ZR+ap04s7akNrCfX176XhwgwDL+oW0V4FSmaIr8gIvX7521k
87IA/fRTNq52DFLBdOx+xmciUL4xSXVN2KHXCH/UiWzW6ReBpTZkW1yYhRU/6XQc
M6gET7HYH0UyC/Ml07PKDfK/+MEKJuOHth7u4xCA8LBZBdm+IYkAHVYKiQ9U1Sz3
wtpQO1K3zgr/txOI1sI/lKNhdIhu5+rd0Fs99KZAwwV6yWJaUC5aHWJ0wymnmHAX
X41maYrHf9DTVifsZk18KOTB9A1Gimae0BiOuscgwNhBvFv+IZGWYRpgjwA1nctR
1Mo7ygD3SIDrudXPDx41W8hCR/8hFkdoVqd1NDwV7c7YQSWukohzGUH3tJE/GOQy
/LyX1+j0uEGV9mD+CsaVYEZcc7QOvK/9NwfE2CQ92h91011M3pJ0FU9aRYVXZp4E
Us+RHXib27K8AFaMX7YwSxddSbrCMrsOlO3kZ9OJUgl+AzG6pnQyTuXR217rRg29
zm/HpVZdH4I84wTdnYZt2r4iipAGxqqfyMxNN9ODxR29/thAubK9TlUxWK776SyG
Dyh2zxboPETAhhokoTsEda2aJG8Oyiinapm+wNs9Ct1LxQeay4wArRZqsIgAF0LS
9HUqRGkz80h4V+uSBwNU+mD9AfKZW6z2xAsR17nGyXEIe/OxbR4/SWNDhATZyCF9
JWW9AhdMBFlnDTm3wRMt8f/EInso9mQJVXFlClOvFB00SiCsgbjolVPPNu21Jhwa
/Ggtfmale0oQFyjC95Xv9bgKVFj4bXukRyBV42AQYZBH8UPB6xzfkJIMXAD+teaP
6Bwocd8RJ8n1RpZhjJA9D2VhOl7LQpwTOsx7M7cRPaSh01xMOCevuWZxteRjuyau
rmHclYUCrBhJ3iVcSiS67s65JR+5K97YUZYfJIi6wOAY7+0G9KH1OdMGs2t8rhl6
SCT9ABg7k0DBVOD6a4oVQoqN2y0oGx3QMBI9IGWH66KB+nC3TpJsakwZwHpOrfQF
MMRu7WlBHMh8aIj/bYmobvnii+CV8pT9/LZoZR47QWo45d1Wbz/6GdRugNZc04jt
/7M8J8X3Dgw7q9hODwDbve1pJBZ/MTlL9gvXdqv48LbE1arj1MO2HtUEmocssYt4
H54U1O/hCvdNIFUZgQ79UmVxmM2FYVrOCj9FZZ3UzQcByVvF9kiJupMLCmv9CY06
s+YkSTG7SfWayBwLoIb/Bem189ApPIb7eVEuLJdOzsY8+5xi0EpxPVDlD8+PrllT
Slc5rbRMj1K7VevLY0hYE4UrZGqXu2Lm1NslFmkkdxUcYrOmZl2q60nw+Q79lBnt
vdHPlNfZeB2irCmRRARRc8gMFC4aLu/ibjh/2VNbBv0nKW4GGbaSsWlRAO5R7xCu
GiQoj9H2RyxTuk1KJOe/1ooRihua4YBMFp1oY/7DRDUzfo9Ron4xX77HJNMzRTVE
v0jgR87wfJk4Dtpu0U+BRPazbowRfUki8obt5Nth3rJYIMZuHhwWr7t/W2E2zl7O
2Wy7VxFYh6/kZICRf0c8hW1UiGxcHMDox5isqVOh7JZxDJM5qhdt7KJ4+odzh4Mz
kFP8nljrystzTu2DNXOZ0a0QwWYJ/2lG+BlMJ/VxI8QgpHTkGbtY9SfEm3NtrJ/A
JbQrWOUEaiBZdo6UEDSoCuIvq1u7kEUlg9SZQ7IIoBeiIhgVo6sYP3nwCV2ILi4Z
+89dBPCwiYGxulaGgTxMMmWYPnIbZdXFPJZ3SgksiFG6uy0lPAxVIV5h6k5ZUEzx
2WnsM0xtl740kvy4n1U/JyclsrbnPxbIgvLxg9tlcrBI0aPBbJwReucz5YFhC0EG
ZfHM/mIgEw/2MHiYwVEhv1SP0B7CCgsc6LVVZyUQH9S15yFdqkk4Jtao+m1y3uFC
2r+YEqHsBy028vyCrJcstS0tCSWfVRpIKfDcYXpl0uWYbHzlXcWAYcoUir9IxFqK
DlV2l4Q7KacOqCwUUIYeKmCulpaXeUcr6lWJOUBFt34j8r+Blhs2HkGxZMTqAWj8
lFnawYlMBccb54LL3ScrjM/8+/lX+TqWg4D+tdvSZv76pHHNgN+n08+0FN0qPLEv
gXVdVryNoqLVLtBqSc4RLdKMG/ERtXoKzqPi1g9U9mxQi6tBVBkit1zv0WgfNOtP
NPMMy5ThwBo4yqoXr0XqVZyulaJhUAGcoytYpFFp9GZtUY39zloklJ0JX9+kwlsd
Nyozbbn6f9Z9uAMwyoa6kFjq9NfqR4le0vNs6SL+hn1J2ZT8bZpvEuuWcwsvb2V+
h6ocsnI08mg+UKr/k1KuSD+t4WTKIjOQngfCRVOHS0jb5pcNMsHuVWb1bxIPWuG4
JNcseZyA5wA7IduZbGcN5mo4wdzObY66eGog4SeBW1TlcSo+hdYc2TdYoJMgrq8y
/UmAAz3HJVV9WPn71Sf81n8eIkTDRBcgCDsZ0znlBLThbWB8nDm9TRmHhhIkinkY
XEeUzMTvADPAc46ZNWu4Q8Emr67pz1RbvrV13vJoDRhp0uMGLGS1qVbV6A09YDew
2RfjakzN6jM9fnkC0PBacYev+G0BkVGiCAjZNe+jYfc+xEDG3jBV5NizulDyiPbV
OLeB3CCeZSNrpUUChDifX/0rxoYU3Nyg+mDBtChb4HwrgRd005fcAG+VeSGAYUC9
JK8mnIVInGG/t7MP+xBgandZO1fmn5AkOTpLCdiJo4WOB8tsh4wfrC2YqiuLtm5W
UQENkzNzQpk4lkRA5ZBfaxnh1+uMMRQgnM3tX3jXJjMZD30cvm3JVEKsiX4fFL1M
CIWe09kQfHBC0CuWV89dBGlkeat72el+96GISnsyVWCiwX4tYNzKgaW8HfaHxhGL
EFiP84v3r/tlyZdMnAc4TrawFFRwCL7+yPn3ncVuhIdeOVt7IbfLCjG4FfbwwBoT
j600qj4pfJ7vG0iLOOwUGtJOJEVL9MlQ43QLvq0AhlrkTc8fF89lAaEoX/zoaoKG
Tz97dDJnyK6UUG+MouFt++iacXVtv2/30pVAVtBjH7Bi9ZwYNPPaB7gbsd+CuQus
NpebWRQC3eGtP3Vof2SO/9XM33N2pBIIoWbWYz6cZ+tEYtg/6kPUlRZNMgMoDVHd
6Pq6vGgCrZMGrO8Oi0baP331/8ZpxNnQx3Rq62FvsOFgqAHFgHeZelhNP537Gyrb
cfaOx5hLrelCaldNPruA8Ys7kePl+ckIYqsveuyAumnW2tlp69co9gIGacEvtPQU
/HTvt9mvfMpKJjOae736qRm1o9bFp7rmMHwpS8tUlZ3kIPFjgPe/qrR0ZLfSsWul
mtEfKZBaExzdLuS+FittmmIIIi5ikkXOUlJq/cilEdLiAQKzqreVJCphZQzkvaJH
68bH4sYKlsSFVcCYxks/FN3Xms7nh5crJS7IwfLtOf4Cb+OA4XC23CxKFJgDTNjf
T9xxe4xvnNgWoQPP0pegxfYtmm7decP81hR5T6Pqz4/baxoW1ZDsZZv8+e52/HFR
WxsT5rR7sfJcgZkX7UHF3mCo8jQoCXaJ4JPjRa8XnqzWbhldzj0hmTT7a1SZ+Sxx
BIglo++seoHgC5a/h5KYKLXW4C+BF+g7a1sR0bk3uhcQCo4sCf58utuWgkeNLScK
NcBxcIXaUlL6uZqCaFOM+nzCEtdb8CAe/MAB1eWsBckgUE4YsXoGPBWsC2eFnsKs
2z34ijouMKRQU7MKj8lmlvITljcO5MZCTct5itsfRfaAU2xbdjzKdpleO0fAopCP
7p11LZKU0gsq7Y3GHpGlJLClzbjEll1QRIznhWv2Dk77vC8iyCilYH6sZ571CB9X
5DJxfMvQjnIacu8KTyZFeQ+W+tw7xSsy415ERBXGEcJKjQlJfN1HPfXAerbwVm5I
DkN8Z61+BaYQg1Yn0SfTGfI+snB7gXhwkL3C/oZJnzcbtERhqz9uKP418ezg1wVA
njVe0KncZAoWQf6Tv8g8Dh9Yjy6AL7cYXRaUFe/civzE/Nq70zJh/YEIilfp2SlM
HH9aTCvespX4gHwGi756I+61/I/YXP+2Nv/yUsHsJ4HiVWCAsIiteVlU5CQf5a7X
Kk0agsMjEGJxEGcRPqBN5u5Qm41ufLmvgBdm+FSU3HPkiltvJ/A8V5YpkYjkL1fb
cUau+zVz3KTEDVnKtMy2ju/SPE/DRsqGnubJd/H8cCWEvMBRG3cxWpgpL66VnApP
Ak5xPo4cxHwvnSQIHHLVJ5HZoQ3SyCmVO++nO990R3K/bT9M1tqc/9E2GQKIV7zA
eIS6lq6k4ccJ3yb08CKaV/jJ8LrE8Vp846yXiW0VJVCQjNfImjMnn4lMXQZaWNKm
jIMqBN6z9FqBl6Q+rio58gX6/a0Yxq3XkowNEQQ9cUM/40Q8lUHcnnca81HJsGbK
O+jFrrLWT+O4KSspA+MD97feLjmHaZ1l3aXXys4xnTKbo9unVM8SgaOzArEyo7z3
6EMKKeCM9vCv6XoSGLKbIA256PGkIeIc8zwz8LOiOGdd4rNjIDVqWm1+FNdmMKOj
WP8CCjpdY2CbKJ5imFR40VLy6gAmSWglvEYtqcp5lwjB3qT8T5HDjNr5yguvEpPg
zYoiH8eTIClAMWUh5GGvQq1O4VXNyxIgBQoAZ+4e+7c9vK304PliYerJewIOP3MW
uFKBdgHYgdzFe19Kl91ddaOl7ZUULtLYqMoVWKgBqUG+cngjqt1/pamTB75MVwd3
VSGeU6a+JrJme8K218v3FzZxeH93fVfl8R53QH445YVxVrNSIuXiN5nnjKwretyA
h3+S9hekL63Zup7pD0ijewq1jBMpyQ/lnV2ET+Efrv1cPxDA3Km+QUW+NEHnItzk
IDN0ZJ9oJyXu+XtfvRgUYYwMAoL60M167rexLGaJathojZQjFIto1y+JEu9aj9hL
CuBfL7McDLXXyXKYzlT6uk8sZLkHmij5YSWd5ol15UiLdjoaLMIoZ2Grkaegswvw
/MK6njM2tbmbgd5FkOHEKhRpuJg7RskPPi6gWTLhVjUY/rWdCByOKa4oO6A+B0JN
FgTU31O7TvdL8rL91F3QlVUq7YHCRwlZzkRHK2Hu07LkUYE5skejnxA3KXH1Zymu
ks3WMkp2sWFRb8oEfnaBw+gcBMO6BgdMc6vWWtg91/NV01gqgaSfnWzU+h+RdT7F
BdwNxFA7GlDKvOXTBEG4rFNqLclXHyoswacwfyPySnzGgtujsMs+O260It5MUj0M
kVrjdtEtLEUtzWBo6PonbYzn2TgIahbJ13z6jwzHV0KuqnkxTJ9mnHC2YFDjqrik
DHc3busAZll7zcswMlqhbQpybjuCBG73ttdjk/nWXB09CQNWob7VtfSC3O8vB1Ph
gu3RhwH9D3CwmeJf2mlzXMDGz2YBG12n6jGEdmIAQoFo/yRuuf5mnd55uUo/Wa56
dDf8rmFSAZCOOGdfhnQVSAD09HCUYTqysaHHQ9DKuaZLgQMyBx0YnT6enkLE5ILP
WMn0rds5Caqw/jRHoRak8o0i9C9kK7QU3VmHAaPCqssOc7k2koFflnkuJTS5pyyh
3g4VD1pO/VuiNj+oIGaZcwkcCnHCJflYKicUvCgh96BBBv7/nxJ3jM7xAWJIV0UT
yKxas9lq1ZjUvBAWalhbM3MK61PXqu3R/HNVjwWz0oriFlsOkvhzmRUgpIDulTOE
tfz0tUtj5xNy/ydSbD2WlwOfK4qcko0iGrHHnOWcfBm0Ty+1Ib31dTQkjdgae6pS
jaIaYuPqMY3HTTdzVblUAzIgTrrdC3ZnA3OeVG9h5w4fFZIDr6TxuW65kdHxo0yI
tjya7EheNk3Zcwv0Ue6rNnhr1PMHqbOYR0JLJOjgGWlbg6alsexaUyg3vgPTVgoZ
X6x+aWnuzY2PR7MLatqVSdza7x5cpeQxLDdFAsF1vBRrw0ZbVjHWE0SYH26Z3J0K
CsC4e+VDXPjjQsBNeeGkkShF10ch+lcpE1ILgRyQu7ZGexknz2lMTOIF3t9d2UQW
+EJO8zNXViLdFMcBMtnzzkwuwSvZM9aP48/CmBh+qPP8h+oipP1Yi8MIeA52WoTK
gaANgb7N6Acuk2/BPYCTjJ74bv/OIWDds1VgjagwGrGqlroFSl6cW7H8EZhkyKQR
XF7QSLbFEAQpnZenoRuRrKxMBAi3wPSfaoZni+py8s39//WhOtR5a3gIOdjBFS1S
d1uFIbK92/D+T7eVQLKH2Gvk4yGx+uI1V+twitgyUCUBKa4+2ORZpTC59O/6LqYl
deUlp5eo6Dg9XpwYYe2lXQT8XxJHjeuCCYZ6spMVAV28b1IfDeC5hXdpO9pprBFr
TXegiFERtfjuAs5bWz3o6HGtRVUWL4N5pILA4dyF6TkkFOwFZVmI/2b9BSd+QBNc
YJtZYHo6N1Rw2xTY3ZmSbNn0ICPFyoXoTxGwAsdO/RRqFbUYHnJIFBS6U4XDIy8s
SqMkyb+Mqh2NjWIlos9WM+26LAQyOi0/5JBbaagToXFhfCANBTOei/f1LLAlQlD1
m4zRG9UxDaCLA6GbLz+2lMdBYdxAKiDWv5g1HgUUFYK88FS+3pMh/hGOhZX1o3Uj
wDY5eN8mx91tm7HwRmvoSFM8uHURJgNpbNC51R/4Qn6y20res5lLad9XIFeHeWRb
HmJ1V45fdQkcue+WlmOAcFfvRrg9MLjQtSexeGHUIlx7LVTTl1H7Why0TbsuCJ1E
MNVwyx5OAq5B1yMQogA5T/fzISS4o4uAjFHUYoeOK6V0CCeQD+HTewY6+WgiiM+e
xeEEWT8d6hdiNDstmc+9REd0L+dtJmiZW3pQooH5j1sIuiJXWIJKV9Qp0NRBqtth
HykosNNa4FdgtQyFKS501Uzd8yPxRn4/XT6STFXPKXvnHSfjvV1XjyyELJzfB9AO
gyIbgoLBzoeYyUggeJPpBoSPhYPeBsDe0aQ4ozvhUm3/qoLq5eGSE4+Uq2K/X72J
/tuHc4JrC9ha0X1PNEoq8Flx9pHNWJpMQ30iKJAeWMrKtaGJFO6TIxfryukAtgJP
gLBconcpZ1uNi1VHuJjLue6K+uProdEgKitNOp3Bg/d1zDrwbVW+dXd6QXKKG+ew
Td5P7+SF23vRcm2cqzordORkNcRmPmdvZO93RFShqFp4/Nv3mTcYeQd2EEpDw9Ui
jM4K318UUgDfwu22ogFIQFS8nzq0G/c/QEFak1ReHB+tM2MwIC46k4hgQg3xzNBu
4rTlroSsCJPwUKJgKVkg/TAw5ave8Vkme0lEvxQvpfQtIJ2VScT8dQ7ac/TnJzeu
aRp6+p+o2mVIUnzQTkPT2FGo/m1ly+B4BDpEyMaq1XtAYpeTVNpY7sbeGwDZ6iwW
6PVveKmhWayofFJylMi6kj3jbOLgGJ8QJn5zlfr0Kb3MPDnLz62C3pNp1aXH1Mik
n1b1OZmid2DCCxoXYxTJvYok3HfsqZ1KiS5AoBdT4tdma4ZgCHGTTPyXdUmaiYMa
4gcK8DLF6jHEXisZ6tVei4/raii1k7IoGBghjXv4BaUo960IteRvuSiEj0MzZ3U6
5fh0TPn1X2B7dcA1Jk1LKANkoP3hb6V8/MdOzqgt8nwVGEvi5VadS93DkI8PPIae
BwXTDvymxncue7okVodHn05cCe6jy+44dK+SFrH8pYiF71pVGc3Nw7Mfc3+RTC19
tsyAz+LNsMtpPjjlNvKFaKoJ6JuMatLX90xjgoOWOFptSTstTHs6S8/tupjY0LuR
vgMupjuD/Bi7gZ5v3DqwYOJDY454/CdalERwd/oJoC6sFK38RQQpGba+z9uPnbr8
y1KMVNAolHiFo8rCv2WYwEem+3MvDYnR77aDmfjtC8TCHgr++RubzOg/+ryZ80T2
dyvhbKxLTC8kghEjY4sNpwfSN9N+fSkhhIEKNy2J3DcmDuXOa+DwLv9xTilC8wlb
2V52Gs/1n5hQe/DOygqR8tgiNXT9SCEm/GlxgQO3Qyr60na9KltImoaV26EkZeE1
dNrDRqFD0Mq8fwkWtfIx2E2h0FULn/5x54O/klOgcb5TQ41+Fa+wIxqFjEv4u2Jf
24LGGYtxf5K/4oKMVFSgqWccWsV1gluDJJpy0dtpkR9r51gNQEGVjO5r50QczsQM
XXl15vjN716NMV4YcuJHuioT3tAkqYZXpUG5ub0PFQYSMTpDHI3SiWmk+NNkVNP9
Fb0tRBtx+yetEI4Ah/XsdZRcXY96gSfhiAPCe0SpQwWwBZ0cgViIwiZ+r+AcA4ap
C5D54BGxe3M56B1dHkjSooTZLpxvL2tvwm9i/vnOYQ0bXZfscImJRlbiXUS2zPN8
pj+wDdnSFt25XMyiI3MaNDvv6utwpaAHjQjaOgh+GMIFTzCqgF+zSVB9T3/kg9RM
h72CvuNICjrFJHZzelxnDRclSjUy0EPqz1O5ix/7/O7ZndphrD9sy19p8TqkCfKP
PQ/I9vqMH4Dkpzoe0ka3KnKtfx2LLlZIaoRlt5/yP1ZWsXY2OevVmg7HS74zvwjU
0dXuLhf3sAKwpktddaK+KV/v4J7j0N3ZD03Q98NP4x82dwCRlGe/KdcOq2EXMIDN
He4LDmJW4pBk4EQ7cEbEQNIAoUcZ5O5Zp2n01AZhTavQAsAWERQRMZIWwRyH2MV5
wDzBCW78z5HT4hx0iEqcbAkxon3N4UwnowT9g908w0QKbbQl9idbEE044pP4tyLq
ri24fT3kvP1nAxVjjNOhHIU2w5geXLXXqzTui25y+1DCsSevEjmiOUwEU9bc6DMm
4YNNGMqyHIuspcvN2nCkLNy0vFCSvwtMAFuzRh6WdDCB1uWx3ObSYOu+2dFQrT1o
E6Cul0zoYDafWOr7Qz7UTh/B6L5mpHJXaL9qzzUeKXdPbOcyYRZ7KXvaC9qcGYi9
LqZw7rxRvYkru2fsKBU8r15ARuahnwqKv+qjP90sQBmOTm1VWavrtwqEccwQh2de
4eSf5BHWEKWUIgRbhOCHHpeDB2P1d/WrGAWi1CzIwi8MJjYOosa4leQDipIPdH7/
cqYRfj2zkt/0mn+aB+MQaJvyN27QQZ/Imn6DTs0ql9VweRD2lHuOTsRokAkaH4Fb
QZ9g6TCZ5KYFmHmwGi3OHjlC4vueL3qbU/rtJGV6pNDPN/iYFSOXo5Q9PPE7EV8y
gBDYhuf27wsbNg7D3tCp3xrSt5lDXAUqiZP0GlHuV/XlOV9IGILbo8zA5SpueT4s
jP/fKTW5rZa9/bJo7XWqqxaqn4YLLfVuv704dtSUnmwjzlQib4dmhqXCLJGu7T8t
wU1XeXpBAFbQVkrg/XZjMsnryiNBkeHWtm6zRRa1pcJCL+VbyAbVaQvcJpDHLh3Y
FVUES9jDZvLNWMEqbv64wab9p1gbdXThuN/oAfeSJKvKUFbrggM64keTawkVSQ0E
iOTKUKk0WmmNvMExgZIO72B6tRCj+SNu3Kxmm1a/vGnlkUEEvSuM8YyRmGGwttaE
n0Y9pOTVo7PzKackOGkniyoKJMG3olLgIckC4Lt17VMEt4keSiT+OkocN/MS9iCG
0xupvCMYSnSxz8nEiqcgJyPQL6y3IudX5ARtIeFVSY7bF7FpXwDwZyyZkzMT4Tnu
07jiUPIkkdFInGcfPXkg9VtnyYpb/AAuYAATUNsJ3uxtkZjiqBUsdIAAdjnO7+G0
kyMD4OqSAeppz1FrueK+ntnBV/vbaBAWCG4nctoqOG0Ap96gObhaQidnhWQ4OvSV
zMdo68e3kZZ3TiKy4esiqWxVYjnf5FGIJzwIl79PpY1WFqTxSXi5PkVwGsNws9B7
Xuu0WagsMZbqdjYy4t3Am9nhI8D8xy72D44F1iJjd/CiA2oI+qgyVoYHj1BYMKFA
QhSEUeYOrLmVvNKpCFAVd6m8ukO0PtTEE68wbgVAGrlNpR1wl3Y8wYSgVNO+q74b
BZ/Be5nqOqNIpJZ8L1om/W+l4kC/Heew+xLm+OzuPjsVxDHfEy9YosH+3HzlTZny
hFW6kEKKVYnyOEu2aC5pd/Dfckkd4gYLxC7FPDmWOdIFDJj7EOaI/rLB2RVz3MG2
dDi3mNPJ+ykS/YMhHzUuBdUoMaFRqNKY6TmsB+ArUOCUglv4Hbs1dwXTecAv5wkC
uzMMfEDRJme0V9F4Fv8cjyLMn3XxXEawjQ0bLI0W7JqjUqS3M6OxppkAWr44qKcx
G/iSTzx8O3iVN8omWEEUk4w7nzvThlF8EBfic285KdQcQUIpKCCaFPNuGVMgIdts
jc6RsWrS502tjk3cFWgVMG8CMn3KH+eGokAflS1AZMwq1FV1pM16BEc7GYaHnCSF
GtnwGK+zwAv4X0PNP/bVrjJGImCQHK+Ko6uziVWV3xjprcZpUEnNX8DtjgfRhnYo
KIQtoOeDi16M2sS8S02hl584afZYPzldmVHbAqKLRBaMpVS60N4YaaAECcoCAbpi
HIXPzpGd6xr0RQibrld3vZgqqLDqW8Q0eMZ8Vi17V0IwwweIp1QqCeG30IoxIZtQ
vefwL4FHU6x/WYp3zGtxy+Fs9jtoHaHle+85CWP1/xppM+o13tPGB1uHH3ZgSlw+
UBY3QqqQD4SQtjINZmxkqK608aIBqVryxUtlfoyvZ0GzDEfEsogBec/UtD55t2+a
bRVx+GSWF3riSMncJ1BR/uJ3PBXEZ9taIeWhqc0NTnhzP0nUAbDOPEAEj5uSUDjq
YT2NOJNkaUNsb5Dyp62nZ5f+OdZy3QD5PLQde3fimOKpssveLa/cyKidgcwkyDo+
7r6uxFCWylJuBzjzMKHjwS1ZKfO/JqR0tq1coeWoFKppTuCnjUu4cYYkcXIP0ea1
/3SCykiGrcpVywe8A/ZMfiYhfpB2hKNpwtjRh8KA5dIG5RVcB66XwUYGhfz7EaMa
6ADDiEVtOtVqoAEZyYyGG+T4QtnQBSEtH0Jwmv/mgMKjlU/WaAkIhzjfxYaDvCe5
E5JaoFJHlCv6DDvQ4WYK/p1ypIzxtBYM+er5OpNp5qXPH7BGl6uV6+xsTIGDQXYQ
vyygdfKsfKKdfPY38q4hvpVdkNjGDEGS/Cg36Y2qXdGbH+GMx4EXWuFGoM/0DPvV
MgfxjZqrQWPdtuvy9dI3XVb0Fii+MpiIGQMnmYdOKClF7fubXSTO+YnUvE5iCshU
MQC9DQSFjIIzUXF4jXw2NlwdBtt9UEa7zi8DIsgLsrAOKBWiNPirbTV4lq343Bk2
vbvSFVBlBpX1lInND+b4vx/dTnB1r+WwUVFQJ0Uy9yhFFawJPZiV9CtwfpatkhqC
SKNGY9Q2uyuULUk/Rz0+FvgAmqd1httfWdaWEvJKFV44owRifnjLIQy/rdDJJEtw
WSL46KlcRImVUri81JgjiTnFbVIEVxrRPegOfh1D5dY2GsSXbTyZUAExs73It0LW
KyqTZdQkF+aKgrjxt0ynSjUgU4xm3mrVHx/AEEuvQUhLH9gxAdupQXEgh/BaBL+y
87xkVIbgmBS5NOC4VQ9moPqHhbmprMzV6TougqzOu+ViI9m1T6e2amM7nMSd/ewX
I66cmx3YwuZJQYokvhJafV7asf9KDQZZ8gVy/QWAa+Ltj+kew6OSDqhY+ZP6wQEB
yibCSfy3LxJpYqIZ61IGkxR8P7EPSAPK7MR12VUIs0F4t17UrJPaSUKnFPZ/OCFr
fzGOF33hBK5IzwZ9GiTwRNeZ8NUbdlZ4LsJcc9zEEE7jmIQpypDsbFblKyQB7ARr
q36HPmG7BtvOFZIDf8tXRv3/eNOkoWWJd76cVzITzZWSqU6KlCvlF+sjl+CTFspC
3HaIWWcPEd56lgrKVCareUk4fPbBh3+SkVABG8QqdQhcJw7PSlneCi6loiFqP2YB
a6slV2HDjsAbBcbbM8IOBuS8dtv5aLCzzUnHQdXpLfsFNyhYIqBEQFxIrq9dsC5/
psySN2j3M+2S9Z+RpN+RWRI2Yuo+JeqpyahRDv/TWMkcjtEEQhbQOC0W85EVtajI
34OSWg1vqN45zXVWY72vRN6lzUmK4W+Uw4zNVU5xtvA0gzR17bvcKEpy2KYcDbNn
8dGxB1FbkCgUFbZ1bJirnFpCeWC99MeVPzOC4AQzcGafVnXUM3/1NN+uBZ+1LHKq
0rqvYMC07NamVtOba19CcWCW24BUFd5MkZvFTscv1kahlUI5aaFfptHQcCnLznRu
4UrnEly50oW5LiPZ2fd9kI+slubZBUR0jNtlIg0Quk+rLmXEerOnvCYt1EtajdMv
qj7stXNkaELL9zsfou+kdsqMz6a+QGsVmbHxtr+1YQjZiz7LldQhXuGbHiUuqq69
8l0QTjkSx4s9dktpM4TT8HqF6U9tivw+uxvPWV+08FOVO/e5qjr6rYbnVMDwUi/w
zD7jD/Nz8ooe6dctqdS3HlYMrEI5j2qK+DMibFHOnS1W9K7ZeEw9gZHPO4TfE2ta
/PUpWfRU66mX8WpJOQZlVqS7qBuvKDbVWSNTo/V587tsU8+LlD5uO8cBr43BdEO/
7iZq7Yr6+YBo0+aQ/7KlMg/CMjUYHDpn0FK7BIifhLx/rvaEI6FEjJmuOVu4E7N4
ic8UcjnjC2zPqA2TPlZIfZqFaFlZtotdBsGYgOf3jKxekKFqvNsF3EDvH+KYUNax
zRU2QW6rwAJ7l7HxCgnG4KbFItdq9Pc7sxAXrKEwppr8ZELIpOvnY/xc+rwoaGoY
LEIfsqKM8Z7mbK8Ke21zyIJb+0bUDj63HoOjXUrKawbPs6uCZdsQwNfUZmPNxM0z
40x52evuIGd/ImX1QPImU5xVqpClI5YphjNheshYdNYIzQHuEpS2Lo9nyuMN/QQ9
ivLn+eVBF28wzEVAgcLiQSS1Oi/9IQQnhmr9NlOKakejrwt3te0dh8+iO05rBW+c
JUVNI4W5eOi2HNo6NbaHWsAz26Sk3w4nLGTHFgpZm8m/Klp4jxlK2OdFDx7/9W0R
VppozrV0h/tLqHaA0wrarzbxnDsrYELeliAhwWD+EKhoY6+JLNr1hIjrBbnP+Of6
ExiLcsX0erZJ5eksaNL03NGGY4fwkWlBIlD2YSj4S1AlG1LHXSM7i9C8rs0acR22
wpE8v0ovvbeHhstF5pk/EdSCehloIiHzM1IUtNO4Ruor/dSBLFlWk9qyg2rdAZFO
NXSSbUdwa+oQy8AX8af7R2j5yrriSOOAlMP4lc/fwWqjccofbKEzzIC+OQWxSg4h
gCrRwfYxZprPgLL00SLD6uBnVQlx1TgoiLZb8VpsFmXIS/1sr2lA+XQmpFeeRhsn
eBq1janW+4X8EPORSvXN/mf/ltM+9te6hkwxuqKCmZkdlm0QShVgH3vXVoslo/fJ
r5cQlopu0EXdCaSQy9l3K8pBnlu12i1rnrL11MYLzrC3LJUUFafILM/R1L6dNNBe
KKvqibDsJNUfMldFjG1N8G9vtFFkAzDvXJYymISjyXptzCnLDHRV1L9zwjiY+rID
vAbhn/Raggux7ewD4Z5uKlfhWsJo5wkNaoia+kmyFO7cqxuM5H0yVMUtZDCowIy0
gNhm3jdLtHapxZbWSbmO4doWKXAmuk4mZ8G77Zcg2XemYKOtFhxr5qE0IIWIbFWn
eSaIJRmOf4I32b1xN3xo3mMdAe5MD7pLyKtEfCD3pojjSNCn6tDTVRbNY0pFppAX
4EABQVaV65VY07BXJS8ADCITdd4RncGsXomjZ5oPLpa5rp9MVpGY873+IJbqOubo
V9/x4L6VsVyml+e7/oobpRBXZOqjDUL0bLarDrXitU207oGn65KUExiIlY7b4uS8
mWWWK8lkODBqvm9TvM8k16sz8RiYagZo64gUVbRniPO2rylCKjg50SdCkDhg63vC
ojOXt3sd5yNyYaeQCKp1fvIfWyc56sFZPLHHNn1hxYsW8db4Xd23Jfre792B0JKa
132S7uh86byVOr8752tRGAklg8WkxkT7/nqr2Oqu8YDHx27MxFhjy6fB+qwkerz7
LUv9CPfUveMQ7IHH7VjEeJQRg37o/KxTaAUdhAEC8jHde4k2+leglpTpgFUrnXNi
vPw+dqHW7uWT0ITeKtXUNOObbOtV+b7CCytdbgAQmJEUDmo9LOjSXwOTVkTTS4Sm
h2P1Qj+oPjX9P+eGBon+MkV6gIPpRkT6/ZWl8OagJbLaqCsmieMZiUzMPFqyDezf
wgIr+c3JDYYpX5R0MKh6z8HUuPIpFBgo6m0dkq20NamhN/3tL81cnXWIyCK+/7PC
rMyQJn5fiFizosb64luFvSlEdwfOiaIkiXNSWJJKY3PcWMS5UiRtbf1UjwwJf5JS
OKFcwVe88kGYMnB+nZ848pI3K1fxqYTQShWBMHRDOPs0tV/79wfXwk48T49ip3lm
w1q4bsWQaM5cMo2B2VxCN1PEn9T+vDERvIz7Z50oO6htbJML+L6ZaLlr+lqfmxqX
Rhwi6SBKQtcV3M/ffpH4A4MuxLiifkVHgaOhQGdI74Ik7RTXqDBqQ9miezmEKEzH
MfPmlqKJVzqHOOoEpQk+TVIpU3hwxce38MtsdXg6I/z9ro8ZbrP+ncGh7ht6FGjG
S9sHgS1qRQmsn+FgK3gup1xnuHoge411DogB+/ti5kkvc7Gk7vD2K8eKKurU6pH5
F+DifSVIkJDkHyMzJRHXPWrnv/qSrgYtugEjTQBP5ajaQ7ep2O0LsIbO0nQrrvyU
4S4zqB6j1J2ZfIcbGjQt4Li/Z5tpAslSe91YG6AmUgavRDqoh1yoSJESg7z46JWr
pQ81PSgDgIMZd26sJX5ugryIIC4nuU7HaBufZkFGlusM9gxgXEAhBJI78Nvp7zmR
q/mOjND+cvT+Tj+geXGFRP9ITweDw6S0UPVmfxgsix68Htk8D4fb7ZzT8iZZSVFO
n0mznaxgWWE0Zgk65GEV+phGXnZE+6VcJL7Im156NXqAOjAmgk2Xx1iEGvuWMRuz
NpXeayIZfAtVwtgS5EJNBsDhQoOBDBmbPJL6hV2KwLA9+pXPZFgza07fs7HrCHMG
zDZZ5A3TC+X0Vyo7dB47vxDfWIm7Gz+X6mK226Yd0Z2ufhEo+Lf/DKQCtaULrjtB
ztNexD1FkwnSPfwlPQc+keEeqKFJPAUJSN04fRVni0+nx3tE5cNgUNISjuS4JpHo
P8et3LXqodt14VU1geWyOOJp7+ZQbsMngtopNpLrpGfaj5NY1kjWiGJvKwrNA0WG
cHr+n6E6/L5kYQcj6yKGS9V2vzqQsymTs2lhHpZn/ZYie6+gbDSqJ+OpkAjqiG6L
ABVIk2rDaETo0MhcTl2mjcLgypiNUwz59Q8eQl8FBNhFbMTMSQR5JUuYiJEyaXxn
UgMLxVs/L+1p1h9n7c9YW6tHeTp6wArc501V4qI5zT2BC9gwdQzNS0+3P4mEFXKq
pIbe5Zp9T99NzxVbdY6HO5ifO5nIXgNgSgArSlzB/J2eCC8EikqDlDlLWVtSEim7
FiMV8yP0nmH45nFVJLBAxDG53gkZbV2WFPIM3B6fPPb/yp5DRwGDMUE87hdshpYp
uZoEsgvLdsdFazBPxv3/nYzqn3zn/iG63W41Q6sH+yFH71ivWt78yPVntI1QyQAR
1TY+9OkHOCNhuLLBmsq6MrdFj/V8yDGt/41xBy0xuko8Hy9cp1xwl0HV0Kb9l6TI
BZ+CwrzBjtMZM6dCxCBNiHhx+WhF4+VwV5mmyhEUu0Rjmwakqnky5HCJKOUzfqUa
KfEwI36tIDIWFGnwLYuVo7M0lffsscJdSG6hHVl0o74hfK56rgFOEenEWM9naLgd
XTOkEongNIaTgb0ichbpK/cpeL0DgLpoHzFj32wTqMIzhAnfNiU0xMP3a10ncWCS
9o3DjLU7gUqHjQYU6CraQKnOlLD+Ab8t5xtdGHeO1yEtx5dvexcpNTO6c/itYC60
K8P2aJorxfslowuWBrOiAFNZIrhg8z4+uY2+5hzLJ2gpyk6319sTI2vnVuRRRdPh
3B+bVXSY+Hl6G2+gVbDDCyhMvQrqR/U//ziGVY/2etPTsgxbNvDVx0L6sx34z6jl
+j5Stqvfbc2jkFxdNi8vFIf7oRxGazrVims3mEZCHLSFEO6OdcjA8OprbG9UgMPT
T3nMN7g62XnMbxn35OE1jm5yJ9Wi08i5ZjCKfi72vDvtkvzL1iEFPyeGpqX5I5Gp
9+d/eluVx6U0hf4VKAPM85etFjdkcjAYNWdkB66e2YOHETD5Zoo5l6AW7vaG89a5
lERHrQfE/HFmLdALlnxe2BVOBBH8zS8cu6Cwc07uqOGf0uX/C07SpCiPfq76NY/Z
EbYO6qFWHwlKep8UNtVOji1XZ9QSXOm/Y1/9JpEWb1HdlZcvl3ZH0lhH5+JT2Ngm
E8u6V0H6cLtjmEpLSjiquQd2kNYRM3LD25jpF6AnYvnUFMvuWH9AY/kjC9s0a92B
Qwnq0YHTm3bq03n81WRBknqH9uOg8nHOvrxsNzm9gdnMR/OHCzaqgEW+EgbJd9L5
saFwR33QuzPhnfMC7STjXQcexzVZxvI7gwZtTJDasDUcEEuXE4gKAfiATYaEMPWn
jpZ+jjxYv6HCuia1KHr5TfPPioQ8HhdkBERfp9w3b5EUZq0z1P9FTD6Jaj7yZ9LF
fc0RWNSXdmMuJ+Z5z4LMSjw4OkqqMMFUVLvV5inl/iPrtkBQM5FYMcoT3CyXnZIA
87EaJ5mZ5uEWJmGVrR+ACkrTxxUHxw1sUebeS5HYszFe92kNILib8jLOr/hYDsCd
Vwqol1bKGsbj03kn8pGIleFoBCLs1DrSGynta1ffNGap8iAsMajdRfNNkxIOVTpi
eerKpll6bhauZ+LnZqHMf/mHnfOEngEcfMz4+YUmbAg6ZA/rThYQKQ/HeqOXIwEt
f9lbPJc56X38HoxtiVEzIuks/z62H6rJ/D1sd4NQsc4FXQiWVX/a6YeUpAh8Jgzt
hob1sssatFrbhLMg8KVXqA/YMRuwHDsC8P0cXCAvzTQwSVLeqwi/b8P/DjJ92t5U
x0BPgCUfCN3HUCtHq/mXfBFak5GBZ8usSXZWfAi8xFpmepQd60WzG6ycfXgfk/90
XdkJMbxyYnngkiWiFysJzXN+rB/oXIZAArSxfPHv8YTM0W1r9KzHEqIJgiDzO3oN
YAq6QmezmNHH07GcX6AV4XD2fyGpLtLeP91uTSebyx+RVCZqTp9rJYdagC3Aw2lz
aOg/ZbaVXsMSDvZUL1r7XHwrUj1c0reiSiI8IatCrVtU5x1EflzmqAD2jTWyIMcQ
nrjTar4w/tPlqP8VZdUHsJAabFV3gGsYrOz5VIO3BAZgLlI8NE/lmYJORQn9RAga
Ch1vDOcnTTDXRk+coQD8mLmYOqeAiY51M63n3A0l+QY40mM9a81ZpxaYz6fIVlcK
j6G/d8H04IsCrcQ+mQ6sQTtHyMzDCE8CGV/IMuQv5OnHkkncv/hU4ZhTVrvs3Ys/
0sb8dkhCndBGuGVwxaTxy9FmkWGppjOaT4kOf4YFn9fQNhWBhkQp4RlSBSwN7N9q
Vs3S9kVHmSRqcjDfxmEji5arFRRGdc3AbeMClhktKOcsOh3UhCXIlDSIfnxzMIGh
x4bqc8Av6qXmWOHFsHMlqNTLUvi/JzLUr+7AAxUL/vZfncxMoTSalVlDVhmt8rvK
z/+FM1qYoSlU4HNVhcQZpt4SAPK5xkmzez9/iN8oCqvJzcy3qE2ehRCbAdBUwZSA
JF+3Kw2lUZq9Y2ge3pvwhLuYU9X/dwxR7tbcUdvUQkIA509L8KpG7YkfHdEX+iDp
ikjHdk1wXHEfpciq+rEL+fb1MZB36UBEjPkmO/buJ8mroAGpc3PGclGRvytL9cbT
K+Tatq73IkVMFLgf0OeBZaU2h5LQxg5S6Tgv2jzCmisSS47Yhj2ClNLKZIy26Twk
IchV9SI/TcfYfkB9nODbRx36DxUG/zkMgZ+6G8iirO9wkLEYlYJNtBk41a7NU49E
N4ccge3XY9t4F+3btblWWHiDsMSpRLq3IgSbF6yip/qv32iV6VSn6cXYQi2jz+f7
BhgQRnS2agkpWBI1TB/dtRT04wYzPgxBwOOWATQnmV3rE7ev2AHnpsazveJMzHjr
uYh/PlVBFiAx7bz7sOEFwRapAC03+spdr8mpF+NNokOZcdp4L1tvLlpEe1wyr4gk
DG3g18dqZBfH/L+4wohRE/5rPAWx9UMRLMsJVvjXEteTl5izDx/JUBEIkAR5Yz11
sKRi1dyVJsZRTcLZUJ9GVGpPRLwXY2hJ78Y6jBEoisJgqHLBgn409wIpoOIUHvYn
1t3E60yMyJZmpVmbLCREOmq2h8BU6Tf83l2suE4gL4QrWXAMaQwCPQMRLVuGJc7d
DvisFZ4UFubvljmrPgtrgwcvd7wUyyCHUMg2Q1LvDEg9wHAJHVIPof5YOamrBXcn
NloW3+LOVnw7zuIXCxZS8mA1TYXtvdTclz9QaExgd890jVKKAp6DQXyKllmyHAFi
+e/i+3a3C9EmS8ojqg0otBI+vFSWkqdH8ozHdHJFO3Rr8i4VysMfDVWEgB5922Gy
2X9WiRFDaX5v8P4zPvP27vhmm9JDlxK0qYkiAJrM5APjBjWRIqp+XZN3kd5zvu60
EjAUKjZIUFyKOLTDe+P7tSF6o3spfiGQIAWfWz0aMTewyhZar1G8ZZHhHRW2QPL8
ek76/ejVRyP8qeWNER8SOZw/UiHR5gmLlQk7/frX6UaO11XJu4YEU+Jydaw20BXe
n+ZuBqJIM9hv2i+t0WzklstnV8wejxhfnZ+aD9NHWsVWsYS3CATXKW6gbK1Go3mE
lpKWXTE6OLzH4YkYxUG61dKMMJL5v2ytkaF7fgl8Rz7ypj7MjUCKzXvv1pzZ7F0K
ExK3Y0sS6zCpZSbTMl7krY1UBwbrfrcMYlP7GbcbrqA1QFjdaU/af0xm6T8vSDKX
2hHBdqIMvapOPOwJnMmPJrk9sRpCCG1COSjSClpUip+dnJzAm5SpaAIjKGXGUKrl
hUiWJUgHGftLzzA8pDyfTstdFZFuvaM1TlCGX6/GOqeM2P/lLKoD7IHsvh92Awm+
QvoUJLV6kqj7DIOh/jitgwk08Gt7xZE01wsItP+oRCtyGhIc19mpCgsJE3bEg+09
La5rbndDXgFJjCyfAuyAU5IC+cYHPCwqkXK40e0iOMnyWxXNy6fKji4tgQA8xIkh
xiQzyKusA2QqiYoTm7TFGUKnQ025V58hUpstYrQh7WPEGbEWxiDiis05WmZYf0Xh
8IuzNuXbbYlF2lfDaOAhEgHTp0X7g44+ryYATgp9okZpN0LE7p7nf9t6cWS45RRU
HMKCXjqAjCC7ecgozMyEjfWYQL/Pg5P6NDOf90QE8lbfHbDhn/xGn5SgmgE362cW
5aSjmCqxtCzwwJmNj+KRKu2sU3PLp5UToR4DQ3+Q5pxIhSIP9VThprp7HIwgTdXo
nhdpZbCjtdfyvJ4COJlwADE/bRtdWHJ/1gBK4m53U4QpWfPQ9M6Xqg9cqWbB9qro
LThcPvmpiefuIZLfA9Hrr+ElCxXJI4mz0YlPgjv7683KhaAxOKMJ1/Zo/ym+Ygp/
NWRnyS1XxSuvu3ntCf5dW0G1zJ8u49tfLbevYbo4GQu/351eUnrezd3OaI8I7NFn
Yqqvjouf9zhWA+Pb0u8D34hTJ7EGWTFbymLlJXHBHI1pcH+PPW8JTpzm0zwRGhPU
LyIiFzjLD6J+XKKVoZU35ohXlJ732qL2kHmyBH9OHVIdEqmNt2ZqAKpIRMZ8SV4g
JNUSk0NMLRvrjk6DnAwgcN9JgXjxdIQVJt6STVV8cgZjBu0BkwYAom/0Js2LVgEI
C342TdqfiGfPDWERr0ckI2Lt28YVJNq2Ed9qn6rE7+mPxj3WlsBy4dEJXt+XNgVz
Au/MlpOOBfkKDiiabVg5dllnIAKLVePP2rmb5oqVle+lNCP7oBF390q3b1PvJVQG
HphAPk6I7qD/b9mVcIpAwrCt1YSCnGt2R8BxMjHHyRMSVsfpa9o58Zy9o4Nt+WwM
OpbkcDzgpemKF1uzeCdf3kXyRNLnotI627MwbF5keQF/1LBSsC68b0QdpbB+HfGA
m0Tzf/aKiHp/y00zEF9x7XKw2skc25JjldjscayQtlzHxon4WwzDKf5WVQ0URmPx
cLG/dNeaXGuLpj4qeNd7XWcolf9ouot0uAew7RWypqk7aO5UWXYlGMprY6C7Yke2
LjH/ICx5FU65t/l6EaxFbtKYFO5jFwFD1E0awg30OQxp59oPz10Vjd3E55JFscJ3
YFAl9HlxtHCZXrsiObb2hAvOg2K+Ab+aO/z3uvTQ+QAsultSGcfayaXKQQLIsh77
SUbtFAvm1vTYLw4p5fkKLTlewrERPYECfGiyLspTW6gZtk1qfbFvCYqnWkE0rPyD
7hI7/cL3wN6xYxOYDYd1Wav0mccmypl0Vu9yzS1/08otG0SL1e9A9dCrwQmNVpxd
ALCNqNGAAGwUpf+NMxfhzYwxixDD+qASeG7LT3j+7bgvyzOnQQ7Kn4uSF6+D2B6a
4l1hmgcMLwMKogPnMEmURnEAWXvWHGFhgmkNP2TGu55RJVH1sPafbWozLv/dmA/R
gCBniYpwN8qMdn8viuUAVTzg29khvzxtg5ePBTKoBwGm9LqkyGY41tWM11dsbGEA
NOvYSYK+URu7QswLYG48FgdVbvaGLRSmXzWOhXXKEYkAVR1z6srxMb53T14qqgGF
RhorGZiODHEfKN+aqBoeAAXPkXGHfkBZvsEOfPvw7n5K4owMEhIlloAQkGNfXqUo
reDThIjv8tmzr8RQA1RglcmC0Q6PaQYRkIogyp+HkH4Baqua5Ln+f2sl9CNoN+PX
saQBg83qQiRn0wIpzV+va5/hzUyYvgkwtuTy9hGmYWJioLVLCYfD+TQoARhJlQMR
inhhbRQFpxOD7xBjUTup4OxCO9uukrYWNHg8keXKgmoAhC4U+OO5AxowiNPRgfPZ
ozB8gGphlYxZgfQeYjgzugWXtkiPf9TE9PWoXLhfedporDx+6sUDt0gKmpJGcOqm
DW7LkJAMAxjGK6LnLvb55B2vgBHOeIBucFx/SE2OZaJrVcm9vKRfdqWiOFxZQwzo
0DTLi1n2HQzYQUogYprsXktLIduOd6e689a0KjWWiFyacbZw638+mXcbdjU1lruu
Eu77OGYC54YDlSCz/aLkWtz5v4sFkpD8Vb0pjLtaqGiFu8w8UslIkxhHrsw2yzjX
mUxEjp+QuXCzngYgyyJvCoy9uw8qRD+X8ZP37RaN2ZmQOOB7lF0sH8krqGzbKuM1
WHykoHwmUoX4hQhUlJ9d+D6ow4pGyAPkqaNsFgLL0D6t5urld/Qd5PCTzp19ShA2
NX4jmByZ2/AQGNm5j8UQLmDAvxXNOAB0FGk1MK357g1Me8tI/HDz2SeIpF26geSs
6atsxRogszsGie1Sk2FqeeFrb0FC+sYhJ/UJzQJcqbwiqTBRLHY5dKd3GBx26Cz8
6VLm6FCnooYazyI+qdMlHNuU7UeZX/zzOQ92mVvVJu3DXXdkZCKVXvu7WDU/ZM7T
qu2F5EqhJfD3yZyaBTa0vNrDg4VqSIFhvzS6GUOuImILQM/m5FQKV8BtwjWdUvdD
wEnep5v2FY+IRRX1TYkt8lmt/BUw2fmBlSZ3xr9YC8uuZTT9u/urSkP1Hl5hKirc
/0PVhLQqYsY0E/yDatkjV5e+Lgglb/CaN1LG3bl0vs7QVl6pb0Oiwjxb1iTlOl3T
y7IBSlAgfQi2iP1spw3ch1pFU4YzSOKwhnBZQVFplAuWQ2tnwEz37e6WVsidFT/6
s3sdpO3/q+G7Tj35EO3eBCe+zFm2STNNl7v97G2P37Z37vbGQKBgSCuoDKKKn78J
0iBa+CVwzkkCKlLx9y6Mea7UIoATuZbXtil5IgNFXF+6WzvHIIZovQCLyFj0Fu/5
G07vD1RyYAuXpyc3S06SSPG53KZ4mlroTdptaEh8w/6Bu5GMw/6scPXe4X4dPCU4
mHjftnSgXH5KKv+y5RcCxUbRmoZuvcZW+D5cgHg5Np7i9TCERSoKXuh3KFohYAWj
pgJPREX5NATR+OPdtm9DzpX+LUwz2LiinD956syxcSCO9hmn3yJV0OtlHtcrGw/G
lqhxtvUgLdE4YYRD+kX8CuM81sFX7sziyv8FSgOS40LlEMrZRd9Kpm1TBPRCtnJv
fDNgw72ujCZ5tH5MVoyQfccFez6Xdlgu5T+LJvoXYzWncGkp3xClpu3KxbYQgVcG
hi3cvAx5CucwgDNV6hq0siBwD54G8J/ArJ/W7CcEFhhwGkH7wNBSH+vXjfD/K52A
UHvdXfKBICRLZvj9B1veQ9lZOfQ1jZq4lJn2LAixQg/2dLj/TGOZnriSFKdfCcj6
ZFFzb3tLAfZeW0iyxeKcvVs/mNff22JpZZ/FAw6DUt2q8br3VAxnWkc8cU0nN8u9
j0TfhwOT/lV0VN2o+jqCDrXd5MuQVx1Uk0KPnjATMAZGvAzNTE27qsgh3kpdfhe8
WmUVPuH9kzpS3V158I8QUHZHzZ+tJnwjUZGwuYLBf64pVn7UCO4TS8VkUFhgKfzT
ipqB2+4wC2tFeQU4/i6VuWdUZNEOzRjNMkpLxtRD6HaL85PJsRj9/1uPQkrX3kHw
w4/+KtUF0m+2BsYVNhRx45uamhLmsUNpn3iAWwzb2X6MKJUmVRcaYpMZqbCs5RDy
Iqh5VOALglZG7sMoQxyt/SKLHtmbtj1lTqlRZ1nYLkEk0thfQt04wybVyPEBZfBp
rnE70SEvORnHszWMM5c83ww/RcFZ28GZERKM1SLjo8V6ckU69Hza2Bwpnf4eUN3a
zeXh0wlx8+d3uhqostBDPA2spWcQmnW22uypKqgoLwlllO3toy/beCYLYcCYK+gD
XaWWVfEjPLxI5d6FW0uRyMlePNS0KtqMQygNAa6j8IzHBbRf1MVHkz8h4t5HDvYg
O8jqx3W1B73m/JgIg7xlNDcJU/ReGzfdlW+TT5Hba1GDwH8vAyhzDhvWELsX/cTR
pqAqzmymqgQ7REh+TzZbRzH2N5c3+tAeL4Zombm2a6In3M6QLPtkYj25BNMzSWbl
9EcwzaMG0dUYQhp7IkrKJI54Jt0KvIW15LFPE85tSYtiietYd9MP9dUdwszsdEMD
PFcQeSiyPOS3vKl8jYZe2+L29C/7pa3IiMiJFa77MZ6QC7wAWsQlA840iLOokJrC
+RcJB9ajlgIGAVC4cDXegYXOPBGdp3RsdpbWafoXRtdmCfoG1qMNbaqkCz0wlawg
idi+5emxXSUr9L2Ze3PXTZkogF65OqZyEW0M0bmcR0hn6YrcgsR+ie5wKm22bDlX
/CTuB4IptXeWz6pJfj0DOl62gDq11pFFdz7pHJfWAny887cljgA8/vFvCeq1yh2B
BLiwlnIN/gUI6cAFpy2oE12wAa0rNjKm9M5FGkcF9cWvJp1MYyaxasLN5DiLnEYz
eBNrp4djpVpvhs0ofZGTGx9gzli3QLu/TB78IsbVR81H6DZMNYrE6CfhrqHcfHqH
p/X6B0eOXbEY3RYALULyCsGunDbUdg0qopN/GgQ+w8/6tbKTVQetXFolvfk8+yQW
UA7v2uJWDStp6/lTKHUycfenlyQom0pgeZsWmslHm6aejl1sI6EehuftB0UZzQSw
FtKlx+svrAGdjmwIuvAnU4fQ8Ykn5OWilY8Yh96Zu3iWasdz5U67GeHlkGm8nm+Z
e6s/Z02N27JVvDpGy76x6vd4JzQk3M3xjRcIvVyve9lQYJHY7gdChMcXnt+AGjo8
6g3u67Bjjg+JPeqAlQY5Z2wiYpxQwcsDRRc15Acanj2v+vpojGtHkur9PIaIHbQ1
pp/Iazl5CEfBGSl3S6aaYi3rY2DxQ5ZBcI265KkUNAV5+y9t5gVKnqI54XepJBgs
OXPmWsYR4VkV6BcyDHfi8ryUXhz6K7D8C786nf6CLuwUoPywkurDICBQnrLvOPP5
/pgMySwUzIFGwP8hNSwozOtd1TYLdQuDnszHT27Igoalxaz++wMcKp8oDxTKGxim
s6lS8tVas27C552fykvAkIvPqi0MGjbbwz4y5Kl7qztLqckVuLIxZrB+/2w3k86W
vcb/Mn3lFb16kZOzycYJqskFACUZBDJRFArYNGc84mWXNcng7sfWyRvNN6tol74i
1+5i3orbu5sCndFZW1888FtIgpQZQGrIsUsH8YlTH1wajEZux7982LmoYPHqJrO/
ua1MV/TULyxWmV2K81fhhw8b2QtDmktqFDZnnyJrUJpPcHq4EVuZhGoCLAariorq
SkGPGfZHg6ejGlN1NOKYuXIsmvq/aImgpYp2pPqXzcXLrINXaSHaUSseHnzj3tOt
YAZ9T1BVt/A1lPegAo/FHb0L1xrmUmylDpwgKOKP4HkyywVlytWCF9cV8zhf5Gi6
Oxe/K0ekruzepJJolkZCeUMoM3gIJF6ZOGBUY1MvEz2sWwtJkGLILPamFPB+f6vX
z2sknESqh9kFaUqYjGE3gH0eP4j5VJ5UN+9vv2jsZfcGgBbhS7ixRwdN72X5yjVs
8wyBYZI/c+lKg82XySpgnVdOWDtI05fzFLteXMhJDiuoBdmWRdhwKshdfdCanaYf
BL4e2gHbj5WAMHTmQq3RnThnwN+8BdXpDnf8S7fTZC2+F+CxIOVK7oImZdeWuPLS
Qi76FLrWHcJe/7iYFIq/1dYiHMos/c+WhwUuzWvPmHAw0rK/X3fKZvE9AxB+Gn01
q82gH5r/uxp237l5kxDhhNRQkwkvmBp93sKMJABD6vtsggTtVFztO08DRVasYHBQ
thKKSK2w/reI+9BvkJyDVOtv28Je2lqL5/ThsFAEKLMzFUKVgqublVUMJph8DNQK
Dc5HV+QxUJoJ2qFcZopOsIqtIqZjA94I8RRB43e8REERgDO2nWzTnd5ojr0dsKD+
`pragma protect end_protected
