// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e4rmU/0XHuTolgoL/kkslAGL6ngIqdsTv7GmvyTl/cU1E+U+cYjzdcDKMVAI9V+4
IdCdzuVofki0fa2ZDt5OtZ/EFdSuKuiSkqvyA5FJQKXgPLsIiP+dB+wSLPnQKHOq
Uk/elIGapn9Us3AhCq10T5gfgKkydZzERgLfJD/LbCI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8464)
RMw1BfWKMKt2Ny87bRxCs1LroMZax/SGeHPxFl/WVRdxlcq2ZwZc17JJkdKYw8yC
xieE9mxDSeBh7m069Nn00limcIntl743KqyD5dOU/5wdKC377RPmxPBsHYoaNMy0
lWv72LqCeW5VpxJRDm9mcYGdgnuBv3A5OGVtc8AgvzlQbIeNgQnwKJyZ6Tt3atIX
lD62BFGPXUSXTUOA64S6viHpDSHOjlIMG4apQPWNo5HoD69IhN5l0XQLpEr2gF+n
0OgpnGhDtp9d59nIIRtRHmtdCJAzxJvHDk/Zr8ExXKLEZB0oz1zEPxgzq9bL9Nik
izAA9ThVeyDweR9YdJwjGhKJq1gaf/gROZBIv9RkUmFhP0n8Z95yClpbkD7wNruS
SE998lhYXSD4uzcKejp/dt2alkdQnpEAbBbjD7l4B16r4QB4mVL80AdfEvg7Lo9W
apOr6LmKRhqCoA1LutC9xtj58PsGbciDKtmNvDKHdyyGB6liu5dj7RR/xP53OXes
m+0m+AZeEL6jCEuW63g7bviaAiPTZ4XDervoDm6f3r1o1BHlVda3BZqMQ3wexKZE
M8PVs1UlJX7/rsqGbgptfaEZrfIolguyl88spJ9XL7Qle39pzc2uIj74Eyn3axlZ
1yGvOb8IVHhs0L1ppZIqKtChc1XbLGy4FbiSnUBErtUVVtVl6+61PVFNPKCrvFDQ
IgxmxmZmZMVazrBXLRfQ8RnBq2JKdSZJYdDShCjCea/EZ5cPaWi3WrRIPkT7c4fV
p8ezRvK78E9gDIvl/bzPS+lQELxI4JIyt8K1DENsQnYg50VQiRNAZuKFHNdonTMX
Oxqu+QNYEFFtVMNm8dXE6VbTiBeIrgqUHwLgzEdCsF/YnASivJTxB6rCWviHgvjL
uYvwlLPtI1yFPORVoaPKsrFTNqNhMLo6nX7ydSJRSlDSORP7p/3sNQiM3jJBIRr8
R3RlY8ZCR9MQRrWo3ZgLLcPYtu6nUwE3ovDifXGHZJxMkbJVoJJErRQNOBQwaVqu
ZyqPZ38A89SsdgBK5JqM01lQLrEcluzlHqs0Y5nVGNOQmuNj4IlI4jgJHjl7Lyfo
VE2SLcNyScOEzq1nl4VQwAQFLXmzfcSq6tbyXqixIwqNzzU0z9rNFt0ojq8WtmDg
2pw+nFeSg1keLKbQR0kUrDMRJ311p29o6kJmMBunJQS1IUizBGb5+XmoEaiMOmSl
Ujn4oDRvev7GoRPCMvrZuoIstcU+R51b6R18t4iZkQylnqJS8R1UzrXQgjU3s8RM
+kf+Z01cMITLOoxw63m/FsGs4X4991mWccXluaqclubgPvFDCO+m6XUKafcE/o5L
jydecYoNV/6lxJFnKHqMJio15J0JpXn8EM83Dm8clIVbtU0sr0tKquZIr2jwAEab
sFgXlEdWgtKasj907AtxM+C5LF3TMqqpK4Z+DnFhD4QOzUoa5FZZ+4AdE5FRkN51
bQHc+D1BZGETDUUJAXidQAEVFilBA5n17B/dwpufXNumvMwMyS9+uPQkIpdncYhW
+T/2rumP1iurYbij79RuF6BDk9z/kKi5hECc+p8Q30GGmgCEIY6kg5SCgfbpnT8g
nPlXJtr4f0hHVZrMK7BBWIWXGNOD5zUd8eLtfycCjb6ElBkKGg16zVdpjnklFzGF
bblImoVHNLvqws1p896S/4i9TTVkJrkQA86b64fdW97t7XO6hw17XettFno3IH4N
wO7K1STL/Yj1+c94hwKC/OBwyk2GMaMiOOG+Er5wENGyuOgarGYMBirj0M0le5+d
JRSR9EZZ8hoZmukIQXl0njY17i/GIvJ+cR8ErOse8Fiz5ftwGflcRH/kYtXiD7hW
8CqWj8Iw5M4yUAUeXuj91MaxrvuhaPY6NgJvbCmX8S1AcM+/o/TjLBHluWE2lbfI
AucsgX//O4BZfD0MxSBNcW1Duufs90byvimDkIsdNy6ZbBYT4v3VVWan4+wvWElP
hHJhlbiYWckgIPsNj0SceZpSDkx1ubDRH1E3pjoPUFXhFa5NyNXiLHrhbsvJIBoo
3Em2GSCywZS9p2vcHkYoQM3FvxKDcwqyBx3uJZ7u9N8SoO89WgIRkvyAHwNq/6HY
S7oQLHAXpGoMJ5tfVbxIJB93g3tLa9Xq1TKivtCYl/GplWLd2itHlZgwIACSddhO
XrICR+cxMspPwgMCnuLl15AWoXDcokh+8o8kEJ36WaLe0KGU3Pz/Fx+43fufbPMx
2yyXq+vNfqkm9/hgUIv4sSEHgq04L2zvpztENr2O7EecO2GGr1dfI9xSMHFu/3yo
NoK+5SgKflMhx9sSS2i8MuDof7vCRXlWsT4+nHcd/A3Nv2+2dnpbqM7lg8G0VvlG
2kMkj02jTYSaq5kEMIWIlT4j/tTGAXt0CQj6iZFjAGCCeyfMW2tEVIy4Sov/gJa0
IGWbTGj1uu8+mQ3766ggMGDL/PhGhxsXaTx+x5M9EAihuSqb40RiEXUEO6XXH0Q4
6xJCLF0cpSLUfaYX7qxjRA99SMi+DbExXX/xuaz1neOj19jp57tmLhSc7k4u8KEi
GRIPUzWG6y2y/rObM4KDGHYT8a5OktZfHD+6kv5hGqqYtoAjMuheiqKigTru+eov
GOYo3Hea/8VSFstYRvECWp7WIGcLpp9Aur5KjnnlJVsB+5HLbnhy0NwnpGWIuCee
kncq+JaWRY1cqysCC/3oo9FxJrowJi7h/ryF8nF/Hz21x0nKFGQ1OC3rovvuuXcG
HWk6E6cg9V/pqWzNLiZyrHfcKhAI43QRqqL7QNCQCw8YA/rrOFLxYoMN/3nJmz/g
EliJHP9BrLtwc6WG8u8med70/tT3tVHU7UvMzPT80Idj8wcOSwUAq4yHUqWlCnxF
QsDf21gMHO7Fr678seW0nAkjQJBBvWtJJNIvfJYzzrxAPyFdQifXHulzvhoFOMR1
icvOy+3hwD3StDN+LAJJ1xipYYRrdkJy9CObdiAU8tl1vqfKbijxLzfDbdkgpZ6+
W6YF9btKdHobroWIM+7e1OL6WtMkxHAUQNTbKNd0L4nYTsOPk9Bdf41QEAQ1cxL8
S31ViRZqaHJGvPwc+YaLwt4r/lxihG2aQMtb+xLc524AUCOcipiu7Xr1W7K0wO82
4qUcTTeGIGtyWWra7ViNQ1Q5aZKeXXtPRlSSg2UjHw3x6om1J3v5xVD2pgrVcRpE
88suA36Zmk3umRrvDXKfJ3zz3ipTu0CktEAu3ijHVNALYvU2ut1kFJHrkXKd2Wxt
WM/wVdIHzMd0F4Q2wIW8lEUPanqAEY7fuvFAdgnAxnE2ID1gYmr72/HmkWL5A541
3fPAHC0jjFAjncmTX2nMgbwqy/a3WvX8GBnMsURKblQh8tZno91jgB5tVrZQ45Zh
o2YW8f4KOvX9KwPiQV2VW9esRdN+2cXdk+vO5H5yZs/7D1cIBI6xLUQkTmajV5hF
ZqIgI+252X/N62Yeyq4/eMsGrMAJjPH+vuH5h4BYIKQyn4MO+0dxTwiyILmnYvOo
yftCaIfw6RZC1lQl7UhskTow+H74AL8UwxkHiH5gI+Fh/l7COXKwc6WxoSKwkeqf
2h8kgvdDN/NbT1yuRcjeYTCXFIcb6egRLYgJ/OFCrn4IsZ7yuCRaUNdODpmmtwfB
PIMVIb6SwDiJTdJfoVWOxGnyZ/tbn6M/weKjusUe8lm/WacXQ5qXNYv01ykHwcYK
AXccTULrxwl6NmqwVTa8ov3OD1x3wVugFK+DSYJcRt9VWVQtvKOem0BXgEsF2Srl
5U2pH+Ddn9wKynwDg5WaYPOP3a7GDSKQuswDjTk9cqf0fwKNMrMj1qT9f81zCwC7
S8hTm/WIlVm8S0A+zeQ14IwIGS8m3Hv/ps6iIiuRPTiyhadVcmE/NzoTPPE8RAes
/VvJtQqDybkiLE3L5tEPW6Bxf8LMld7UZMRr2IvnOSmURzpLhZA3Y8SCJR2zTh5x
aCSTo0XTe/3/Iv6zJWwnEMOdwRMCJEc5RA3AxwbL16M4ZlOwuYQG5gqVL1YRLE52
UtlNonZ9pcyx3AHOjt/sXggdYcV+fD+M1SvHAtYo/DZwdYNoiZLtpVGUcTYq4d84
abdV3d+RJ4p0LPUDxEFsOr3rrwWXHJ5zNEadiV56lvSBgmafeWQ0MChnAUlAFgza
nyycxaYcdF0y6aBe1GOzwgZ3UKnC6x7iYn5jAhcuKca5xYAcAQCLKL2kRt9uyoMW
Ze5nwGyOR1nIWfv9tj8DNeQHgphggYZPmaYcdLDl8joawZepZp4/uVJ1sC9xWbPw
ymz3goETh8tKc7hwP8sMBbzMTCrHrkK1G2LcbJQvQ4kTSmFxqXvC3i1ByE9d4uXT
8TodP6bcb5YikPeTS9lG6bv5A8sIhKwvULypdJgeQyeGH3SWRcwbjiB3fIGrTpsp
yDWFJysZ19AvKjHshP6EgYkxDoZdNydaiwtaOV2WN4QyA0DFHBeGBeUf5KhzXhq7
LxhfOq4HqQoGYXl2czvurXg62c3ZICkbCaUZ4NL3vaVirV+UKb+BytzRuCJcTkZ7
H+DVS0BqH9FXweebmspTeSWEEPIih0bQly6/XazGXmKxPjh3urkwc3BB2fINZbDk
5nqETtcEPVVpSDEEuRRTnugnShZiVYpfSvCrZzkMKVM4zQXCablsOl3bRlxzAqfQ
RCEPUyRPRSPlMMk1sGRSJwKnxY5STzhNcQ+eBv/CG2Iyzwft3X6a4J2OhdExaE7h
9pS2Nu5fUEv/Bx8s4pp6biKqzsl/A5bdOMRyFA1ReX9SxZFeu+AIcG63YsATKVAr
BIYFufnfVl7Y9if1HT2Zf4/aJaCfQqgSuWkXKfmx9cZoHWLYiIGisUAFGxsUj7NS
PeeubK3S7ECC0fwOc6YLcojKkXUOnpT4LyUmNxGSSfBFww0iZKHOa+mNbI2dPu+u
iUfWTnhPonN29Z3jmtRnvvAR0KCTiYov0ivhQj4iYjLM5n56hAb/yhcE/nlq668K
kA+MqCyNq7m81kww1RXA5dvjr+2yMsA5Vvi510lYAZMDy6LWwFReBRvBxzLGrt6f
Fxd/Hxl6DEbCl/gyt0aMAFyiMQGLCKayS5aw82SBNuwQgfzTdFdcQzH1PQw78mvk
MzopkhlrBW3DwmiSsODXHQi/MYrk67DzSLDBW+Y5kq5ck8oaygTmXyUWS8AuRV1y
GkiSZnbdhznLh+GmJOQbxubEpJ/ih9aJqaNd4UHbPC9zuksHhEp4ikqlzw+OKB3y
dCT+lmqGZfhEYro4d8cM4IlZtmD6g0VL0PoFyMyYOz517s3ESg7ZbVXFgRZk3FjT
YlFpFxXJV2J1eEBRlspSCNWSjgyCbtNhJGGLF4muh1Jfg+LQL3xMfV3apvnRhomO
7HAnpBflpF/8qURkG5Sv53LtD62v/plNqApRMBDkwhBHOjyGbQUjDd9LqbpvY0Mo
iyeN6SfSfCCA5N/NMhQnNYA/1HFaVF58iMB6Jw2c413alGw7H6/OjTSFaBXRPlaO
grkjzqK35SMNVBkL9iuFHfJ3AF50F24w9S5paBAGfEWcb+y23ZGBib/LtWsh/zqd
dlsPACa8shGDKnTS3JCDHc1lurIN6I6Glk7fN0wH4EZlcMbyq6ciFbbI4/JzYfil
VOsPh02jzlMqr1IPtURiKAeBQMHB9zDuPSSeP1/K8idXV6UwfkAXM20a2htHwCTn
5ffcD1YgvZjeqHue5Ip/ywHKouh3/B3Rov8rssD+EVlslB5oFKF/K5bi7s7k6Xnc
EAy/5xbb9QtAt2ZBsmgC5Qq5U/KLg8Doi9dUiaHoDblkvHoPl2xDsvgm8oI99EkV
6WEi+a+zA4MRrdmad7zGT8D5SRHGWZ621AmCqtVKZdJhi7kS3d0J3rdD14OVNaHS
0k9pw7wYJQqPphzi+NvoYWa+72h3uguXeHUhhFVRohFjXFJXkgByIZAIaQwd+TZ7
UfZtFB9nxSpQDCBTAsxohRk6U0yk83e/x3hEW9zwPRkgtkhDU4HV3VqohX2/okOh
ItsJz8nTPp6ZaeBg9epHB9yc+dEQwPob3HUmngg8p4gexutnn9qMNEvKEDGXjAVf
u+9xz4xPzuB5TGEhwVR6Qtsuuo8woQHXUXQLgiJ36CWs3yixrx4AfWV09C3ildKi
X96rleFUeOmVjSUchsiZzjHdBg709kjbr2fYws1ADgVOPzXVYwL5OuRCN+VeCCcT
MLiumsabOqGr8eP5+xwPdofH01fByxwhEM7PeeAbsNSRLU2sL5c4pi3GO1KJjBNS
SRzknDKWs5Yw6Hn+iH+FEB3iaTQ83Py5wQugVMq7EDiWsnTHAtzKLn+tri3gtuCR
MJ10VNCWRQi783vRllofNYm1ooBB78ouBig8wvXNAQLjFK1K1FQSamL1XNPt1SrY
HqGOa0kgNI9RWPBa9evcm7DWYH4wNI2Xxku1qdzKosiKCtDJknJDjof7tRaXu15h
1FT068S7tCuVsYJdtNDDJxlMlD0owbkigURzZekSoT6GFhOmbyoDQlir7egy43AC
Me7RuhXkzDxOGU9NRlJbYPkU/XmAqo66++c2Wg2DGObdkXUBfcxhGwghjY5gr9I2
b/1+TDXydTsUU4/KD6o/znwc/iGmH/UDz+kIM/CBZ1btYDOm4kK6CCPh1fXkEzL2
aIuCyix7Om5o7ZmAEiYUvUYfqW4KsztLE/ffnvPnq706FnN38y3j6fPt9YfsimF+
xj8kL40MfJvrYfD4Q6tL5kolTTXyR0Ka6NAilHctRjOklaoxNxFUWX7jSfyl7ifW
UcIqQ+65tf9BHM1OLE8w7QLS0TA+nO0eUX2tgIkyP05GrXdmN6LHhXXYWh+2vEFS
i57NwZTDq1IV4QJiB0wObRCa5rB2FvX8r6fvIPc7gdETeE40Rg7+IU+MHIvVT8SA
hTaeAY9El8MlKU/asr8fDCwTWMrAunIqzNrngTRCsDRnuFsHPag+RWW9QMKOESKI
HAZY3vxDh0YBdITq3a5uNARrg+1oyTcWKrv6TX7SWoNrtiHrRnJo4UXVAB7gAgP6
huVf4wnXBIJUn6GngeP8UWFg5G2FCNIoa+G1xcGcw5vc0waA0Jmuj4IBsNmQhZG1
e1LWRYPubsURbs5YjgZIFFZrjyU0HEavcfU3fAVxwPuHrImM1UbLUc2zsYKdc23P
VIy49gp28saQrBSzx3RwuVbpt3/KviZ+EcwZte+mFSEIvuUptceJ7iCGNPFKPot1
4vNqOLuH/32VVRdqR/51gtJe/7/i845OBTKTCO4grgv0gn+EVZKa0/fv1gJlu1Xb
qTfFZm0qhPyeaK5J4Lw1YZGmobbhC4qjQyg+EHnfu0vJQN5Fgabn0t2ezzsTEeow
yC3sfNkxkFRtV1PIhQ24BVSXzlrqF9vQZwVnw3oc2/qtiRruAlifASl9ZpiYUUDE
I+jHl3DDyRkCPtDrUX7jxhkJeWfk1QDWda4QMHzWcawFXZRPvHhd/ZOZqPuWOyO3
WXCbKQGUuL9Q9h0mQ2Kc0mdI5NCHhpUmT0TIeW0JFxpOpo+V+pG9hHaNze1MiQHl
G73iBpgI7tRrEI/AE8odIqGXFAbuFdTo7rYm9Os8xkcV0vxgNk3hk3Ohe+5KvYyO
k91dYZ4oDB65SZmjH33oYi5eWX5gEZ88tgIJADFiil+hsCMUlTF+E8oF6546MG9/
jiGsTcrdR/NabZ18hbtGORxbhiGrRDKVXu7eOOeHN5nxf3lm5q9cGiiOB4/8kOFM
MsDhlvnuR/+LJOTyK3bG3w1QWWKxRM54+cqJcEZ2Nr9ZvEO5PG2pstEZecotmTJP
Z6lwoyjS8bImDW44ZZgloSLqKnZ7TCGQy084jUda1kmB2KiBlPCkLVONRU4vHtvp
RiNVMbVN8Bv0YHv4h/qYphyZFP8I3+UawF7Gl2SAC/fRWUx9fH9lyJxAXGo2Cbop
j+2ElarplvCrC+aQRPO3hI8S80++qFSQJWDVMQdrBNEq3bvHHkZ/bBJe43b2+DH6
E0BGmvMXmwMzTpq9q3QP4NMMpKRPAc9DU4KUC4IG5jNiQkunw2bg4JP9pbKw8/ZE
yPRUKY+6OpdohMnfB6EFb7oPwJ/53pxTfNyP/DWvKwpEX2dBmCZ0fURquZwn6pIw
jB/kctjr8X01NksMTFxuq7zg/gFKfDSqwBqMRUZ71VmuOqfRIt6yWPFcgvMcGLSd
pxP34uP0TEcp5Wt3xqaKx5B8DvVEaoFknJ3Z5fbrLLhX7f9vEnHnyyGk6t+WG3em
2pvFRRdVEFNogiyuLtL7gEJWj6g3GwQqYldD7yGY/AZRJwopQvLu+LBQxBIvxInl
PY2NZQIJ8mtXj/lzhUNk+5ZvEGheWvCTE5AXyYgM2vDR3DKbO+miGNyj2ZwmHUfU
aQKKf+nGDywC2jpifOrysTgejNyzO7RBMRIXvZkHL3axLuhAAIT0eE7afAA3mpCQ
SFJg9TE/gBczH5qeLoA5YxuxW9qYIHiTktSj6ysQpzknziEn7hc+ttZGV4sEUdN2
9DmXg9qcmwvv44j1+J1SO+jxWIQjLDnyw+rsuaDyjPm4O63MZ24M6ZLu4m4TgY0W
zSSCgYHPUeI+I05iokFdNqwY9aJRMWOY32POd1LCXrUGRZLx/Frs0hdgDJDOgDNE
rke9hegu4QAzrq6CRKPZRnjybz5wQOWzdHxQ/UD38AwJOOLo5KjLibTo2O8mxE45
Ql4T20YkTSVoL5zpGET9tXNozLxqkqJYkZL3CyB/4k68H6IgbhZDquOgTElDCLa3
TvcV9LWv5OhkJdMAMOcTbdRye8qLlWKYlzz0bBK2OLq364v49/sC+B+FaKZAFGeZ
m53bMYU68aALFSg6up00NLfX/91m2OWKB9fGlpnV01fzWwpiaLQzUonVi74HZDMh
T4TVBNvS77C2U9wQdqlFhqKMZoD2gNzKNAk8d8Zh5k87pkeff0NMlDv7E0kurjja
iLdmIW8t4sdnxQdy51WmPU5PjJ7nG6OAtIsNhqXErL9HXNixLae+2tKEPObuWs2x
5SdxKXVV8bCPK/wP4s5+TVMd2h84vz9omY7KPpGOwOveQBGDl7ChhZJNngUuOckK
zXjPXipnVvvBiBoXW4V4e77QpPzakMAnZlVpvFWlELGzbMBtWMXj+Vmowsn6GbNF
np8ZioaWIxEgUX8S2C9se1H5tS7bTiXfaS1VvgmBqVznETQka1jXdizr/tPihw1o
0+XUVRsDpYlrdkwiGaAYQ9VxmJYt3YxFBTfFfZLp+gvIArEN1D4geUlaIJ5cgWk8
zJwdszZdYS/yXE3N3fohnj5sOzd66wRMz9+txXbrDyTKWIRiPLa+ejo03X54adrW
Y+vI8mqHtgFJszX3mzKXlAjuNM2f71Wu8qitz/CdAlK6niQ1PcuQw80F1Fua4VEz
3x7QxIGAOyh7P7IfVu4cKtl5XSms8iL0Cq5jVbN1Ddz8iqNsXwZ7EKk2JaEn59Bh
RJwE4OemNWJwBB+cuXrtVk3jYHd8NL8Ri2iTomxFvjsTukWFVDQyYsyJafTxSnSR
2b4F22TpEpvGR19ENgMaod5Ph8rMqQraolRvJAMms6LQX+VgjIlK6y2YEgD6KkMr
8o6A2gDjlr6aiv9WT7uQ5nrtySTGW9gs6ADvjzeixCDGxhLQnVf2bkoUwdpSlhYN
AI36Ba4e1aVWf+FTNw0yDCEst+YDmkW/5RW8KcmQySC/X0mYSKgpChPXlBhuwGWh
G4XhfFcM46213CHuI5MlJFhH4lKDla8lotVuufobS+btUcu/+65Wp+tNjANKdA9u
jfpmM43f0TpFZVfAyCwH0N8ZIB9jy4+gHbgF0juHBYBwFJfpLdmCUxwWCOFR7mk2
aVj6h3Fa0gIK27Qi1EzAkO5SrP7NNeL8LouHzJRJNgXoa4VLD6BVYiGALwHFjenc
WOjb8P9bh13kV99zRBE66RJxoLDEtge40E5QUoEsfMHmu7Aobk/2IXlx6ecCd31e
4yYbb2VxBP9TVJtn2fYjnoyOaftVXFn4/6/pKm2AWZZKKpU7qZVvv1qzzQyVut5a
hJcNk7/8i35GM0DhAAWIKuQXyagenss73tLW51yk7yFTjTuPNT35EUCulI+nzCxE
PdwqTcpkPF2zRW1tyy6Kh42wZffDdwqWC3w5mfVuTz5dStccQDA/PLFE+jLclhzB
nB9fY2le0Ufie7j0z/vXgLNgMl+QPH6S6LG+P+c+o9Ni9IE34gO/yXP7atGvzGY/
J9G3C9Q/F41AL101Ubur9KQcJx/Akq1MY2LilMZ7RsMDXCcXkWP2N1H8pil6oLDi
GdAmHifKB0Fa09qIyCOMAj92XDBWWhyKzVG85sweZHWzu9BKjWASpEo99X5QLUd4
3CfPAepJ/b/9Qb1ED3h8ex6mKuk19xcf7MBIvLQTCkIrH8I+zu3d9ne6k/tbZMRO
XJgYBddtByokVWwY37cfvDMGpV6029MZ0BQkZBnDTPCvvZkQ7y0QiovZwxGK8xD/
h/GXJf1SBbfku8uptDn4kk3xyg5iF/QANzMN1J/DqhizfCSlzOm80xdhtPIP8VjB
va8JjqeMoCU+uMOsh4O++tJDy6/wPL9PnfGI3dAI/E9C/dAW7bW4JIjxeFLuZSRt
vOhtNd1A6+AlU2kJvJWkuWqV/5q3LYvowGofsafjdMHEnsC1DsvABuYyU3FaxyKt
EuI9SOlvVy+n14KwkQfocurbhOFjFBArvrGWPbts+GAcNkzrhkR/dNVDbwZ9fSn1
SSJ3m/VzOFk+ENOAsP++pXy40mgBP4ISEhRMEIhG3UxtfWiFqvhAb8ckBABu/eqf
TwbgMwMft97VBf6ObquBkC8STy7mz2fp1hd69tWlgXuqH7hYQ3CREGJFM5LVBcoQ
MSUNeDfZTo/XsD0YoZTkWm1TP2tAxNZ9Rr3JbYyGAiOU3MIL90JecKTnbVIL4F+Z
tw9aT+UHelbDVbJSBkqBahERLuZr98AE7LOIgR/l52VV6NA1CbCPQdQcX9h3AqJ1
LHlnhMXiWD6DIAAeOkgjIqqJRZ63WGj7xZ/Xl4bF877KDIfGICi5U7LuHRF2aoA5
hLidwun9G7H9xQP3nr83iIXKWUcqJIxMFctTo4x94DGmci2tBLieR8Go+r+/wx31
jzepN2+hYqtiz/zJpza+uNyt6iOKTdKW8BARPAbWHuOl0cqna8jCsSNHOODLSb9Z
V9hE6KJc5F4avXhkAxtOXAcCf77EHqx9MkSwVihvEaToZkQaNzMXlTVpyMalcwwx
TkBOP3ltPGn4IkvsZO5Bpw==
`pragma protect end_protected
