// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eFKxt6iJxUpuGUsUHi1O0ueOoaV/G926z0umBRPsPb3xZ76Nq1G6qufR70wh081a
aXDYWwwTThmgS9302iQA/XSfrX1akoRVr8rGKC2od+TJLvidxDiEcPpSgwOOtZhc
Mu8c1fxIqS6dmNzbEHJHKVEgnbGArpzy9cOGtXCzu14=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19504)
PKwlDEEyq0R7PCowsUdVE7xuREDmDHnPRFn+Z35vyXr0nmiPq3xEFKeugtWvWV/W
tnePWzQAGsaluzCzRwQjlUs0MnykVdV9TZRzaeHUg45lTsfWcCuL/fBF81uADE8o
1OX4Mls/8BzZwKlTM2afnZLNfCxAG+gUgI3UFTIUft0ssq6dKlbeL1zzRlefBS9Y
XUwlXRGhPeChn3y054zwIufir9dcI0LdkAychrgSRCNQbEa+A+WNehEN1xS6eVHD
nv5VgRvQr/kEekiXCLk0VaNVMyADbtfc2ypFMKuwOFdqmNq3N8BrucmcdOrf6WEz
K2My+LX2F78Eu6Vn2TxfMUytvjCgbvP3YfyqWD0Je+rogFbjmSfGG+GbGF5LcA57
Qs7cx3yW78GEm5dn/qDeCCKe/3T8rr8bzmcwSBxNz3pUKhlyjD+xiwfC7TB/xWN6
CzLhLOkUzGpWp602gvrjBXj2ufdGaUFFXsx1r6kk/Ws6qdMSKIJezGU4ijq83lKy
T13ga/BxXv4YK0n0HNp/Qpzy92aYnU3ob4U1olxpx3J5DdwXa2IwhOMtpipGRzqu
p+o7dCEH/gj6ad9N7MTO2vudlxm8Q8EdI82wmBZqh4YAOKnfC6oGeLKNtD1/Q4wE
tjbJV8ZKZjM5LZbRgPRzHGmRMSDMx4awDX9iy7AXp+Cp3miBIVvweDbxf3Xb5ir8
wbKUTTHIYFpryyKqxhUIAApOh2RWnJAuIAf5fr2ygb7E4iDxmHvCrx9YS4gyUQqY
i1go/Vl6O4ODZf8y3pN23PSLca2iBjcmvJP5pO1qtOwIe5Y/E5AOarLj0jg9ttIc
A5EPsawsffJNrQWjBxxlIfM3UXPSG0Y2Y4BtkzrdImXidI0/ExczMEbJOu5fAPr+
Io+npkqS9ABh3E4bRSYuPjVJ7HgkXrl4zYNJkjoOwu2CgpBZ7yhCQBsOd8Krc/0I
16LLOtIrMUDEn380M+kEnRm1OVQ6fVu2h6BKQQh8pdf4NJyk3JJAQkcpqJClkwYv
XxPSdIT33aVfpvYby/yZfjj4sVw0unrXWnal+HWkUqBZM/Jf2l5fImhrl96bOjGI
D6e92b/UnfcX9qXFG1RVej9LeYZrXhnaXtt+/A0Tu11INxbvETS8JVJf+93tUjwr
BIau/mG0fZG7/lij2X8S+SdVi21847BVXOiFUp9CXvYKjkNpYa9Ac3s8YPvnjqcV
GNtOq8mXlaSUoHrerJyPBtavq5R4/wCYWfkrTyzLy45D0dJY4SHGwecgw8pz4spI
a2VkeX4laq4aypjT2aiKYOuloQWdMTnbBoM1emKcPM6qkuQuBSvHGi3xdwYIF8bR
KnK/EJCkHXxsG0VX0jtHWjt0NwiMnnX3QUTFt3xdSFJhCOEI3qA/4LySTkWZqP7Z
3KhpaBBhdmuan0v4/StZ+0HkJMjtw0k/uYG1zTDv4mVr1mUT4hNequ9NauvYG5+S
gWzkOajDonN58jsazTgL87DTaJ9XyZ26ExMbqrKc7168wqv1dPgw5Bmx7oBIqv3h
BbgGYqQAyUzEdb45gxevl78iMmgkPKJ52xJiYTQqpVhxAR5ImvOQVcoXUGS6LxTH
R8OmOyvIxwFKkUzJmMyytTyB/TYL8SA6GzSYxdfznFRGDT24JshTJgbNwsOBdX03
B4D8ip2sGM/Lotq74tGFqS7OwIGHj1mNaEw63Tq8bq0q8j5f7LkSun2QQdyoGPq+
8fzXUvRdzGkh5QbnuEnId1KJiEH3XjhQ5afTk9hDl3NjaTv6P+Ymn3ZXpNQrogl5
nPSldBgj7EtKaPxC425Bityd9rwAMz5UiupZmpl+EjQesJUymD2TiEMs00pMgW5o
+CKe+oSG3z9fkQpLiisF3HHw32VWP9vvlOi0B0jvT6RsDzl4huvteGjYAPJpkZvP
nVm4a8KTl1y3SJc0yR9DSiihjzh+uWq/iYiVKu2O66M5RjB+usBQeGy1GH7T+xvE
+9bur1YjPKjeOcUuLde5Rj87HnOB2FYTVbLHIw7Xn350bVY7vKfmiEuSeoUWWzdU
9SNFdVcYuL7yaNsW4RchiUYApfSWtakOiB6/mg2xC+YPF91WwHTf/IG+w2Mq7qn+
5N2wPxKid7wrqnxdcYMXuRoUrWbnxYqQli55rYfQa1kMtgnBKnC/4/iLiBSeD7RT
84ajPrJH+3dlfNpW+Qs9CpibsAVsgI3usREt1f0sUlOllziCOplgWkVcZerU96nt
B/6Sbs7qsI+8lDFL987ByxjFoJBRaiBxSMWMayMub3eiaKG16nQszIADITYrpz1U
vSx10NeleDc4nWfI0D6tO1+Xnfx8wATHZlXsnq3UKhFzwH2iWoIJ6a7hOykkNfZI
T3QCe3eXV0uIG55LkzHLdPRCz1fJjP5p4Ydlw0onx6HFAH0fcmJQVQ3l2vyvv5GX
4OamPIftkApGEL3EdSPrhimX6qK0tD2Muuebt3nx1c1VMwluReO+L4iq91uQ9Qyb
ynpRk8N/d8w3fJ1ds6czwt4C8sv37NpqOVurWi857WEQ0nNvbOHRI5IM1LLwGi5B
aOPt/muiSo/LgCR8leSjsSrHqsWxPD1Kqjz6RlzySk6nHoqxH0fY11R7E8hNvj35
omGvhNkYx09XrSfGnZH9HxHD6AGo1zFeqpvv5uS1G+rAH/R7/uv7S5fWCrRNnZ+j
SwkjjW+m3d/wayFZQD4ly46ILX7sFddxR2KJBmg6ks7RCOBSW2Ppfw59gSeUEDIB
wjnO0ft3n6KyrZwpXlLkN06CkSMT2EO6LI5dg0B/niBI+iqBcI5vahmFrAeSIxJ4
2Dp0C3/gmClq4gRV5+9412kTe+P7KfUScJSW/52cc6eqGYPK073LGvfwrss7wlYv
637Fu5+qDuHWCpvlgPOHVSwtfQN+kgZzG67py41esPGjD10oVzgTfrREPp8TFCu6
29REHy1KJRGtoIXOVZYG6t+QXJ2D8ry77TpoA2Y484FViIvB0AHw+T2ubThKa+CE
P4gKgf6LSfGesBOJWOJiiVF0wQHZawJn8qtnbiLQhUOVHVee6eHaaDOXYNzY3aos
uRrqaE7zFP+u7Otiq+2i9dOB510O759V650ej44t5OR4MCEn7qnbe0dqbeLbEbFg
JNaRVdGII7AMioNzbd1G5De18H6xPCNaEfTUV0qXb3hxNl1J0D6xARN9v6JdpN9f
JIrtnrexkVog4/WbggAZHblQmZAaGCjYAtTyq6S+AJWmdwmasXgqbbPkY2+viUIm
10a/C6oVcwHTA83WtKGDusb1oaSGFZJfs2KMkI3H8sbulzbz8Oyg2OfLkDfxkiCB
vTg8KMBF+o0jOkUAvepf8sTS7gxCdcxUyDNb28Ia6F736ZnRvZ62NeAVSLuJiWi5
lgcrQ58vkST8wEYJ2px2iqsUSMZ9YrsQegFgSMW4/YIbVT2iyhvuvFYlfZgjYEjW
JlARK2utlQV1cOIuzKYrBIwyI8Eh5JggNAYKaHF0DPLGz+agvMnh2PNHbqT+FCYi
HBrPKc57bdBVFsHy0BdW4WIGXNtiZhchVLz4BPav482hnCzMc3GYNCXnySDdGbji
12j+lpDC1FFlB3CNj/Fjy/jmnTkrUsuGQZhk7Ef+nNaC7w5PS6JT3KoMaadAUtev
HCH0RHmN5tNOQqvJ+8wGnHQqgL3MmNCl1hpKZc9BMLpsydnmNtWmh11/hHHzQ3bQ
ozyBKNPjzIfGlAw9n1pevqLFmfW0dgrOYjuG87ptIyCo83MhhiFZZt6y6nc9ipT9
B9tj6lxRJ4xk9pfczXx7QrqfhUjwW3lsRg7Vre2gDuJ+rd/8/gSdqOYGikvTNE3B
juVWjzYnelaJ9u0BFIfo4vMmCdE6E/jFWTjPt1fVHNt82jZ3txluLX4/iTVayMNk
zJmmX3x4AEhCxNPBByGCc9XUZxs/J3Y2nJZmXNM+pSO2rJ1GQQUzqa+Regf/VBwr
tsXGnT+WKvuq3Sqg1dplFJ2k7iEnKqxSaocQc4T3p44ndercXVJ7GI1RzLM5iIxn
khVA2YMRZkXG4kbKtxc3+sC1L7tUPFjDcIjI7tX7wetdNGK6n7Mc6LUJ9ZDM0cyz
nNv5YC1N8ZmLe5y9cFBJwJWgyNh0hddiyWnWlBEooCqW5CVMza4zbLs0LYmIo+0l
8dttoQwQuthtazj+340YKMV05FkPDe4Rz8JodHqOna1jOw7C4FDsjyrasVBpF9Zx
bUpQtnT7libTKALOYe9P2s9/97kDUuSqh5LXwmM7FHE1ALI1eXv8w3MYP3Ncrw2H
7eBLPB5D8TolIOZQGvC2lsQvxg3ffoVDeSEQSRpp9ZsYZAw8wCYbdvZMeT0a0qUb
fcxYQ/vDP/WO0k9Bqdd9pYmIu8ybqLXLunMkIayHnjZprZ1Rx8BqSxGtyw59kZyz
6ooOR39moO2Fkwguhux5FN5HmHgHedh/Yvr5qaPiJAJrW4Jbsw8nhaNrYAK8k8Nj
8Z0BpNE6B+JjS3loiAJkbsktcNZFPKiBRpKwMgifGWP0SYYBdOCP3uzK0OfLy0GI
uUYr73X5Ds9U4QhTebaSZ9o9Fv7fKL5yzrZYJPMiPgXxQ4rPpMNn95nwEqv5OnN1
GuJYBtKv+sWoj+gX3XGFc0jEeQAhdcFjiaUffwZ3ZZ7HWOxpBJXm9MR+ABrjXnbR
/FSHRaeJ87W5QikRLtEgYAGLHQ+BZLErv4UQ3Ebm0BtXpeD/ENUh59wQ7TLbaRZ3
dJHuDCmo04cGegaP3n2yN79p8/UuWeEIEK7YoHQr0lXd4sQ+yoNidHE3NWu6gNyW
UrJt7Zs4Zoks4DmdpSss2dq66nFNusByOjMw0bLoYixkY13Vkhz8j0BVB3J+RS/0
ypMsNfVdXVI4wnetbkR0iGbYVfPsdj+z4U4CSpQJvdp/dmcIIo3OlgguIGOTaTSy
JaphNrh24f7BEwxZHGLFDVHQah/qIieHiK5UyTeydipAYpdQ6FyXg2hfK0Bm71DP
gCkFseQpCT9LcyndCSFGbMkr8fYfUinGXRmQOHE+GYkT9AiNJTz02uzXF1nA384Z
HnNBBUNc/P7Bnh/nj8DINlyq+YJU5iI7jvB3ftwNiy5UZnwO0eh05vPzdY/GUlD6
hmwqNccBlKJAybaYHkYT5ClD4Ip2MTntNuHy9BmOeNOxjPyE5xZtZX37QGJfltiV
FMaChLtddOrpDfqdXhDrhMImT45eXeKVBjl185en9eToEaRiPciEzXDn7C06HoIE
maCPyHLu39eZ+8jkNIkeTipFEe5iaYdMlOMXpA+a9hO/REJcntYoRpYqoLNp5Gvw
iGBvE3N8P4Ckn/EH0rsJcQqJBcSxjU7GauPG3N7RreD+WqWRmvQX3mYX9P620rxa
7ZHOphuy4Kz77ei6AGkuL46IFFqUkCMXLZMn62CCfbshTeegmqbnRM7wO0yRL5cu
lv1pT/ix30ZcE353BF8/+ub6Tu0NRIGHBXSvo8HbFSSes8eQLl5H7Kb/iZqws037
yU8HQZaqSIwqnjerUvUXvWGgEVLsoQXBvPG5JQWqKuGwNzShiWevu40NTMzMy8Fy
ZpQg0m6lkEKlGZxBQK/x0z6YYSbp+ggDqP7+5WU5pQa7yzosnwQADFxkr0uiUUy3
Pe56QNLoSPHK+na7hO+SUw8YFwKmmWF9TVzrCwyYo0PjvTIIjmlVrR11WQn3T7QE
HczxioEmPFvjERz2Qcl4hMGBNL5No9mNoBgv/x6u3oxmSV3gG/VlyXAGxwK4Nv1S
HEemZwouTn+oMeW9FVcZZ5EOk0osY3YcE6IJvrqBjqjBgDS/H3BfxvXJWS3JgWfG
Q+t1KTczoz1GEYXSzhmPQuVoqzx3/nFaY2kxT7lYF3O7oGOQomyyDC/uxuXaLvNO
WqVRunKyKWINabyhKNkkdri5JqTZV7JAbG2pk96hzG2HOH4WjsCOlvbF13oDlaoT
35XDJeIGOHuRqYMBbCVaWNSUdjB/ory0ttNdu6b8E8Z9AkvkpQ/4EWUWyDgn11ep
XCYH+3vh/fNe6Zx3Qpi8WLg6gfXJf0NSLAbyyfkptyciRQiMUH7pWvg2zIfrRrbM
WP1Ctdt3HjDaq0pu4a/WuBfnX0PWDYN5TTIB2ji+Ow/q0Yt65FSyzF6yUCQ1RiYm
PnGHlTgqSVPjw7CF1N7T2jgyEsGqDdDYyRU+kNiZoGx+EpYFKdRviC+E82mG9WmI
4JcPLqSG6GCf4ZXWDMRv4NK3aaVgungMUb5GnT7guybh2IgoQHIHSjISgyHUKmdv
c7OFYwLqXoJLuj02slPvm5GBAFCVWGDapvwhTuAlYy5g4ZttwP+Iis1a8iNnuF0G
xdwAVoTFEQ8HpHqrTsrX6DZl6sNLdBqluIe+tuzK10HM6ZE6uz2/BvG3bqWao8xn
0ejL/amjgqRZ48haVy1DJOwQhOOxZk8WY8dL6EFPu/gsI1n1GqST+/mv049GEehj
vlPukXfBvT/2tHOzMDsGWG9g1C4wUUOQnQfF09XYd64VFspcPUyo4Fz7auw+kUMS
oBuMAn776OdaPMtAJpCqIWeeprZ77CAXQDKFLM7NLfwNBE45GHl0c0awiHh+2Nqw
meVCBaxrm23C/W2a8mJg4kInJN3DBxKgfJjtJB8b7WsjCTGUEiZglB4aMfazJqiT
jAOORdcZmLLdBkjRBld3Mtua21bkfdOKaxGIIHLpJwKgIQIrr8JVLZQ/p7Xk6DBB
wxl/0x+IyRAvwBjsmUx3KW6CPcYUpzutQno7wqE9bEmTtUvJjwDPAo59hheZ8Uua
P0lC9DnSaz+YwSStXmkT2zD5FMVTdeql6Nu+0TC4tNuD2E9i6kgHh2BKMntEl8D7
wx732CeHZsq96OFeqEx7OfDpIgMw9wjiGjEL8xyD6BTJAyTKC9LUcFAnwv+YQOe+
gXxB1wrVsR/XTZThmQ4cdhhQcyWdVpjPiyJWkkp55k6ocx6q/xDyH/fd7n+W60zx
5nogBzQ9QiS9hfClyZs0ZyaepVe9DK5K2CMzpbTngLPXHV/JUmY5zIbj4TjTNGBg
ig1Y2IQycgexCNbIvLkG8lPSheqMPvLSne227cR7eubdl5QkPkME2eCBQiDg9eb7
J0z24KZDR70pZocJlKAYMxo+3zPJzt/jyRMAWj9sthKVp14iQl461FQmE46yEvZe
8IdKrv7bsNtxTZrpGf7jvcHO3EQacXY9aQnZxyGnicAkazgbKCUvfIUfXj/yBN1H
ISSh09MPwnIRApMBmnxAH/wcprPr6MzayrTXF0ygpqNQxKM/yQctlXFN0XyTahH4
+MShHH4UT13mYr/wY3rXylL2T1729fnRjlXjdAqgE9wNXFwvUEm1dRWhI/A8/pRp
zdYSUzyHYND/YgpYD4n+G6UjUpn4+F1odqpddpkeAwe4d39MKpmnYV4E96UXtdQU
pXUI+gviQJ18WxsVOqiJThmk06LyPPb0cwTNcCRQxjZxetSEqqEN8vEOdNjLnSUV
jaPoXsGqEoNF0b0Locj8WE8CSFSA6zWQJfIADSZiKPHUIRb1spS2MCO3ajxIPjux
7ITClEk+1UFka/6aozxDiea5UGrYPADNc/2O1UYM3v3JEzo69TtILTf8UxUPVWRm
MPCuo/FJFpRduDizzIq136NUL2fUXcJHAMgfcTQVYVlvld5Y6TOkvbidw+GCrDgi
6/Yu4p4tdVV2AkdPpBJwZD746mt2ZAHYWE5wAn04HXcsls/wXaZUpdi93GI+D90p
2AuHFWgx7HlmGLKHB81ev+9Qx4ps5MZbF8L+vKpyn8HUocH77O+iSZQoI9kYDgdn
Hs7VZWC/fU5HTGdhxu26AkBZ4eMavTX5tb8aczUIvU1VlSP7ayMtiLZm856ptrlT
VNpSVTFlZookAIwdraxLWHkKp8e7WTdAk99YRHQXVu5+Aj7KDhqoPGVQ6lgo3mFp
KYiDuPVj6wLDLO/NYzpAEx+s4gdLFO9mThta9VNawlmZgZCaFUxKh3uypVCzs3IN
8Z3Gbl9q24gXXr4TZloEhwflPBwZcYSVMvpTqPpTXpYS12zZ3sajXD+YRtS9O0H5
Nw0xBMLAnOqu51V/l1dn2dnKGCRzU63ezvRhDUnq16S1vL+aWuxsYDjE+KrFhX8F
3CNCfC4cNb0Ca3fQwL5hl4puLDKc9O3NtzKkc7885WUcGt17guIsmqWApwimC8Tf
3B5GCJd1SVe55RflBWr/Xb5RA5caTxohbdwH1t2iRRBsMI5e2qe84Cutc21cx/kj
V7IHPq3n4gvBID2nXrlRf1PayRL3c1s6h0Og+4xNDKV+6bg0iXvdoh5BVooemxAO
RwBvdK2uYNw31bcWIp5v5InRIlJtoj/gFPoi26v1wnuGg63lsk9afRqTvO7fUrnt
rdIgcECm+V17wVSiXLtGC2NYcbmaflBOgM8t8i7GSEpf1LBp0hjGsQPPecMwWmKd
KRtw+zQ5aKTktXdAwYZ6EJV5ai38FfCiaiC9HzLR19ZYT/0q+noylDHiv9Dptt/+
DmWJpK3g3/qYtxhAixlkDuBqtNrC+inKFIMp2LCiKG6u+FWSNFlwazow0N/sIyz1
75daFgcg2eZRNR71CUOehnH1q1G0wu91f8giNo328Is++15tqCGh+7gq9305bVhD
Wh+RF4WOOni6i0Gafa+4vEqTFBAi6vyTHbaJvjHRu0e3lIC6TPoJNxQIqTYZFRgX
K/FS5BbY1KVHT0yr8BbGAJG6orUagqdwRB/xIX4Jue8rT2ugsRfRH68oiToIG0R1
tIaxuBys+9g5u/qmyDJu7XqzTCZktEvK+gt5ulY94ze2P8jrGBWnr222hPdG5KGe
903goaiv3pFAk+YRvs70KJ7e4ltp0U9anlGK6Y4HNfQdw/gQmeq8AeIfxpIElDTW
cGYH1lP8zEzWVUj+NN4Hdwf/nBv9/76X4StyiT5YaDAqBiVNif88wcnTVnFx2dz8
86ZXWpgEYDYEOor0Yj+B0KB561tw4nDrsQ7v2mMRXlwJY4T9CYjqJNTH8AFuIIZl
qpswQsOrGyP/U913ZDheQk4/1ibLlJNDb/WUOkrJT/2HjoSJXOvnJqI3AX22A3yw
CAfYniwqPPJ2BK+mlxBxwIHcEJZO/OY0t47FOHlmGxeI/+acDq7HWbGsRaCd0siH
m49Dr/sSB6+EBYTVlw6trBMtFdzcrQ5MtMlTMw8wGuLJHXY8f5jMOZrD45GK0i+k
Gjjlb232kSqELpGemA1KaUMV6noIm44W6UUwmRgTVTLbnQjw6Q6aDhp719APZdeB
WcURN3xAqGOFKjesVXD22GsVJzh+s9b4iebH1Zqdqidmg+P7bt+MMWN+algmqDUi
gupm/hNT33NEXqwx3jpY7VxAsyXt57MyxoA5b4EC+EDKFJKw/1LXoPac93xzJBhG
7vEOPMtnqWq3mP9jNgtet+U61NMYxTfue9jXlwAmp0ZAYdwSiToNqMl81FHodZpN
hj83rB0ELszaCJ5eWEjUq8yzlQuQH6qwxuE1lYaGwRGF1NvNEJQwZ39US01E/MAj
Xj2F4aFsQcM5Mid4NLbUP/9MsQKkdktmaPopLzdLfmvg8BVbRDsF06lYEtqLq9K+
jjaBkrreybi2MNcgN30onmri3tRN6HcG7R+pSkpnzrmjspOs2Bw4w1rpzkGRjZ69
WVxiLK0IuXAvUONL4+qcGGoxrat/URFBM526+0Y3Rt4EwKvb4N54CRb6rxcg4jIO
fdHxiJMkBvDYUoH0lx1BRykx+rOfZHdoY+5MNnEasA0MoOVpUtmv17MlFX15qwJU
8fj0b0jtdjILgntUuc01Ss3eAaaoLkm4xU+3skm5JuSnKPN2PNSfyH2HpvcUfumj
PjlEqROon3EqecsokxGsjLJNHPl92XVlCatWhBx/N19ebSXWiW1isFDV9mp/L4pG
9KOkuyCVjat5VAodowWL2GtzaP5Ij+bAxsa1Tv0StPdAFAALkFry8z5wH1wPgufk
jBMYD5fg1SIdL7pWW2g2R/kCFWgVFcvyPr9P7fMfrcI3MNPhKgSkDJOeT8pTUJWx
helVguyI33+W5pGA6ibuSp/raExIF5iuOLx6zOw85UN0ocey10X4BBR4gtiGqICZ
UAren+vpkRJmtmmxG2j1/JA2IvacgXkEVNi/SoMzArfab8wpMd9WQtP8gM9NiKwU
qAOzu0hH/C8/rACb2XHP/ZLtknZJzWMZNYiojABVFIzC/VXVMgpfECnJNetpMENw
7pvVXQw43WWg++3NrVBgBFgC3J3bVu4aJi4XagHFDNChnlKHedJFqW0uV4bM5prA
sHm98vFBsDi3VGSe3hywL1Y5ldKVLPa0oPxom8r+UQCHwCqdBJLA7DbkmnRFTNYJ
6aJJ8NjoDAGr1vcOxbTywU0pw36zqHYbejqY/G0BPs47Z5gHKFsSRYz2f9uNTbL5
6twcUGxSeQqF1IauDkS25Jh0MhpvlBracT7Ts+IJYNjhzu0Y9ilFz3LpF2AlPLyh
P6PfDduJ6R09zvVUPInoz9lLAGCwyxjmieUxEPRXsnVSBtzLFdiW5kEYU4za2CSE
N8IPt6et3vzeUz0v+GJhYlwH8H+iQ43wSKDiCAPWcrTZgxPVN1FWQiq4YOAA63vX
npHuQW3mFPmaauN0+W4OgkktMrH+OaCRNhKin+xrP3bx6Zsq3O/jdceP3YOQNX1R
S36QJPM+Tse8D7qQD5C6WGpy9nZJn2vtSIVydXKGKjAeFO955beQOmhE8Vx/u+Oe
kIwbA4OI1hAQ1bYORWz7qIqS7OPdGPxfYRi+Be9fOG4erJT4ISacFDxWLMtg/kJS
mTntXBhq/8nKtaycu6C4mwbcl4D362hqMRHuJB7Xu/TWoSi94cRIL7zhRoJVFPLS
/r+9mzikkJKQGY869XiJZ8CeuESU8li7G2E2Q0q0hl5YgCwvDx5+VPknBQ9ac7tx
1GWrS6Mf2GqUvJHBBt1ZuUZ0Fu4ASKZQs8Au1sTiSc9SyWqj//xtpOnNJwhHxrAg
L5mwZvyUGaytZv7blQFgFLXHLmz/VpmM3VEio2OUYVa0xDabmMxjIP29FI4Yx5J7
jgORqmxT+5RYA6aBVoaxZrBkgBkYlQQHX4pRBgefvIzERYkXK8ixbF5Ef7UgBFHr
rURW2oXy7Bx9KlDWywERJB6Shj9cwqe+zK58cvW966yswk8uZUzSCknCll8vSfTz
nuQOxEsJgbgyYB/zol7pdzAKp48VsY5jfG0lS6TRAq5ieNoS6tLNgTAedy5WDEn7
wbbvI0lj9YHBiXPWLUxLMkuZwN/US73rjcc8SlM9o87D0FydtpccKdiFhGsAZPDg
LMmNfRVTzY4mHZmXhYoNJWDF8STCtjdIPzVuKuVcCvnWb3HVKOj7rO7k6m6vQmyQ
7kjT7Ncb7aF1lBO+S+5h+dvW0Gf01mbhXdFyvI/sr9AjJVJwdOgW2GRvkNQWD0OO
cY9DUSKZPcHYU8javOLgW8oQwdFjI8vTLF5b2DGAsX0FDtQe560xgb1dIkBrnG+w
hrkNmWN4G6YGkdtLTXyCjnRTWQVhcqS+EzgQrpXViiDgbVqFRWZtJl7mi2eNta8W
GgtDquFXFMQh6QwWN91sCjYAqGjz4ODUabB+NSORpfZncj88hmiR95YxD6iGC6P4
Lfyll7S5Cvchakeu7SDX5V1GwLEnP3AtE7rY0sZHFKdX4kXyr7rGTZig3aQqFSnO
gtjDXFbYSCwJNfi+lq3fNhoqv5qfV3awCRYBTaLvE7EyjQaa+cQFnCTB1wAw7ClY
B/1xVoFlaCeDTAa92UNAw2XHLG6qmGsfz73frpUsf4dLwd339ZxPspFF/GLu33aY
axbkOk75b5HNATRV/l7SMHrkTNv4xUb7WedMmwE6+3TunfdGlFhxOd3RqvUpBBh4
gskf2vYN0xJ1J836Ar4rSecqi9xI6+pLE32K6xN6JyiZe7k+x+piCbTpNMc4wcov
259Kda9ZdkbRsl9zioX0F88/+7hLqEZ05XndZRiQYPI7SrsL1ltQEpN3n9491S6w
RhJphh83cIHZu7qRwpGaU+UbZpTh93f2tvtr9PRLDOTaYHNDzDZZrx0oaZ3yHS8Q
vSSAJf5TBbN0JOV0QW6tI9eZ9HPhySY0HmJW8IAcYGecGj8dq1WDJneGcGgrFqMP
+e8z5sRxKXfkZXKAbkR5gUvjhA+Uc+CWtmuNDEE8q6x0C2BY09uDfyhseQpshofO
8hgBOIcBB4Y/BtpWR+Qj51mN7tXEGz7dIpxi2lqHc0PqI7MWm19GyjLS24ykEe8A
KbX8IYOFhZHAc2uf3pHgJM6n1ILOMxTdbjN5oN9nPdM353KtMNlBP3+5TgCxcgFd
Wn8+TPk0LBG3xQAEEZtG7BW1fvEqA44sc+wo75juPkpCdqasQydqhUKfof/iwJZQ
joibPsn82qBJoB/SSdAFmo1bIjYxJAobEizkzWK/N23wFTVwYvYDXM9s2tgvdTKT
7fUFL6xnJlt6CNsgKV95D0+nHb0CdKw5X7Jpv+x8wwP1BCs7GGuaqh05RuVGcu3I
n4kCoO8sKbn2nQQ8Qu4bYJ9/kFwIG4k7/9IKYu240QtAHP/eChfjt764IMJ7HzZQ
xfJ2mn9A4GeMk0VBEUAkZeWxTKMilTLniMCi8dFOB2O2F+zY/rqCWI7ap20GpyLt
lhC2xprcds5Zi8NKUEtFFs9PVt4+uDBj//lLIEsx1jzat0JIiTilNZ/ibyYJD4/U
zbmgNymdhjhXHViRUoG/mLmMSXDfLkBIiKqH89XZjK/JC2EUoSUVW54S21/s7jz8
mMqimSwb0OecCF1dV34Bhk7DY0Clq2GjaxSEISXX1W67r/sCy4FgHHdiuD/3ijo1
JT/nH2BqwihcmdlgRhaLEjGCqxdD9WSKJ1tL28rF5m6ghlGQ/9qjTH60s1SisTUY
rg/V/B7er7SHUdkIU7Q65ZmPtVagUyO8e+57KNQ7hvsACNtjgzzb5UeUWNTvUxKO
den6C4m1yylZ1Zu1HBSRfH5n41YOGAn7XYuD82UepTHsbWKTCi04Rv/Ku5ogi9j7
Q6PL0bCpI2OUztklit3VPmYeY6fg5aakmeay/6PGrGKC15VPO6qlp7nWtX6vG+oI
4kjwU3tKTuRuMWghaIekas6/dCsDOfHSlLyRqx4rw83DZOGwa0y9Ps6iCVaaywyL
jOKjuDPR5oO9Tm6XTLh7ZY85Xw7jJL7dqOwhw0Nzuskr/FYMrQ1yIWSk/HLUyUhQ
r+7+jt08SyZAaEoryCPzaXU6R7zrmbDKaLWMvGBInzljmRCtYAGLn9XkMm08Ml3G
8kgpcXDf2Ce05P7p5P7FEKE668JCARim6wqtZIQbs/V/1+AsD7Jg3zMawQfqVUm9
SXKRXf9VpAtHJHHXJ2O9gXKVBRqHQYaEiPHJEXL/orGGSSNkRrX2oFQe4X50Axy2
eFpwjgPAp3jkcWwolwvYznx3Xtq6QyO5xkcANCQc1vFiErnURhQcPV7hH6KD0LGS
xkEC8x/FibmzpNYI2PukWIbH4C33Yb50uT8dHOpqlL2XpIf4JhqYpJ0c6e6oFfaF
PNZ0PltlyRM4TXAQd1cv92uObmzQLxhPmqP3w8gZ5kUw8SrQAckm22Ac25SE3yFB
UOz13GLgrV4eZ9SC/48owo+lYaWCVeQPGf+4Qywr+ZIeec2vjRBmpkWQXaxCtyKo
rc6jsQXFI/dIf94kQrjWFhiGW74TdY/y6rCghoMiE5z/c3gB/vL97mpLUFZ/Pgu2
Ce32j/AHefip/vTCR36UposlIdTe5w+kMnO00P7WqBAiS5v8AF5EXXLZDZTNuQLx
JJSp8yJTU7SFe4tTXNapvCX4quQ5aP1+bAzyQT0VHsaDdcl8fst4tJtZLl2lW8HN
4XUCs92u/jJpdLS/OhR1/9MwhQWD4h4ZrpG7rDfoaLfOVB+XGtSigPg8C5PYIGJo
D2K1Z2Dng01BxReabjEwJta61iAewC/ZQdc6B/XbeXJf8/QB+YK9R8h+XW5a6ta2
aj5mVn3QSwFl/7r3kQTrTswFR06KqkGNVkrTiHLF3dP/sxbYGggK9SWX/kU44sul
/ySVg2smFk2LS13fLrvKYE5l6o/OTdvIGxnA6grSDtEAGH8a+tmqkEuNzLciUH/y
x8B4CvlB/r+2xLIHQ3zfsYHmkkjB5X8/yp7KmDLYF0uvBJifPO5nCFR82tW5meLq
Oq4cuYPwDGaFU/nGMblUYjA2gRSB1ImA+GB5ot/Os880xRq95uuAuKOabVTImJL+
lw5AU3swFXfsbyQArPYrfo5HfSPnXuZPWoItpmLEUQ70LfQGZLMFJQI1R3qV2qpj
2ljQrCosco1MLoaKJehbDMIj6WmlXVAhxv17AsfWzgfjU/8GgFzDxZ5q7vO/s/cs
OEHrPi+LGmQNuOqkCXxhy0e29ehVWV7baWp/tpZGq/PZT5O6i+aup8UK1zzjvuYH
Xz9Su9UkudiElzn31f+W7TfxX7XOcV/TSTYwGNttXho3qUrw7dD/lxldr9+dd/R+
s0b5w3FmfKZTC+iybX75fGBIE/C3KeJ8IUN8919+Mj+x/3rxb2BKi+WnmR7+HGwd
oNbPT2ZrpRdimrtaRLKTe4L2R3FfDHCs6j6FREm0/wgWlUhEkoq0V4x+N8jW5WDY
2QBNok6/pRiysrnyMh0MEX+Kczrjq/nLj2R8s/MXm0zE826kSrCPE9eELRaBCBm4
hTOoRpUhJ0cArCVd0aicSrnHS64U9w5YJ1YAbiWTphpRaE+akQhkvYLY6hF8+ROv
Sbq0PVK6h1wDVR/GPafOZjD1mJj0WTyUsMfWCKqWkonApNj2Cd47v1zkC9Ns9dx5
LHpMdY1lW8bFm68KJVWdJls9IsIbfPsMSzU3k0YYdcyO9/l6LChaGm2Y/D8xgF6X
dgmIab41zW52OH/BLDUQTaXF7WEzv0vWmWIQkpNw9Opq/757MoEVlregS9QllRoq
onslIphnofbLfFY1QleOhOLSgOpaV1iqvpSmUispQVF6vZsZ1vpbonwuVhI8W2dF
iVxrUxdIFIBs0rT03UHPD1+vnMFKBl+pPLL9xoeR3o1rcQbqVT5zxvNiPYlpxsLS
8KDIgvieulLSOOKfqvohh8gZfGMzjSaMllRfT5AWfcVyMg/RvzEQ//k6Mpo84BsY
6lCIPaVFO1FxuREJRWWpVI2mORbolFB7Cb8SuIWX50IXpc840PVbiepywhk1wMK+
vsdzHMgEsVr9xvTyH9Jo/C0VNoP8Xq1wBUyktuqxuurV5+dAJulv8QgDhahD/9rD
brYuvY+uuLjgDcguQqNqi1Jn0rMzI7RTlB41JLNOBVEBvzxWJkVlJnrVGr8Z7pZs
dfrFxb2QixfH87tCCsiY5iC/5UrOkoG2Fkz3qtQYYLs5H7GMoHRxpl/szup8sjmc
lQjDKM3tslbqE44evI103S4waCYwr5qcjcprHKMPNVtNlDFmXrrvGiQ6a7jqJ5DQ
ex92Or+ViiDN1kJuyf1+P7swq4L5h5ObzCw75Kf7bo+A8DPOz78I8qbYefSGMhSm
F0P1imlVWeoD/yVVXD+JnCj2+WtuhMGpNkN8mfqYo/IgePPtsr0Y9FzD/Bk4tylG
IbDsO3Gz3vGl/K3wHjD3XxeA1lZYBkd80MEpODGEReDYH6ZUwaM3cUHVnjTMLK3l
Km+3TqeeT2BsEAvHjzgI6CBS6YiKv/RjxZ/bmlPik83RHmwjI9pXoW1DnPqGVgg2
Ezx6CfKxSNbQAfEyDzVwDOdq/O+kYysEqtp0L93xSUcJc5Gjf9b1EBJgeoWjrs91
cXeonOcG8/Gk7eR2pR4L8z06LGyTCgkMt1P0iZkAZHztXlwde7e1pomoF+N8ReUf
yFiqpShpFlopuWUZ+rzKX7oCsez8zkbF/sIybf4KsUDRiFUJiVw67xOYSQuc0G16
alKeJ1erCIsT8IZ6REoIOewlIrOwQOOjgv8d0NJb6i/0najWWeB2YqaWmome210Y
/ffZt1jbpt6jlQjgzjVZbvjMcubu6d7eqmabRIiUqoaJhqnG/xKOv1nF0y2qAEtz
SQHBsezbhevgPRZHE0uamPD/Hzv9KZwEzHTrgRfTAMKX8UC1TP2bGDv0BM1mFDr8
7BeS8d+L1aIXLkZ6Ii8RvWqh8ee0GuRXQV0KC2YOrZMlhRNs+VTytHSL1C/hugIR
d2/glFJ8qTd8y/Wl75JawP4dUncoOAzlzRKkEUOI2g6nPaH4oHV6BECLJ5+ccZRJ
fAa9qrdQR8SiSUWYRUTTmryAJmm7P8/dk6kwg63wDD5DmBuXm/ts8CUnWyg8kw4S
M4NG8doqzuX7KzTRh43cXpWqLk6xFD9StHC8AiU0ywdY8CTHnOtc9ItBmkjI64cC
R7Oi2Xj/d43EvhCiMqa0shyY7veqS2OAeh4fKK3jPAA5ltO7wPZX/Axt3lK/HZiu
c/zxwJbHwUXNSa8cJztRo/k/qqoWikjTAkNTCgJs1Fvg9w8IHKheajEkAGBsmOsC
Y4JwBlRSHarxaJR58/R/96cea2AuWiQ/l8AGae95Y1gDmsMyMee1bMdz10enWcL6
QVWnBI+nQeCJbl72ZLiY7JJOyok2rQT4V8WCCCCbQkVm50+UOHkIF4HaSu2bqGhW
HhVnRDrrwBwILnp27rYiEQv7zpkpNANkrxpmmUREnt5JnAWDxyYKSX5mDboZw0ds
T20QbiR23dOEwY2QtfkoEqxSZAjBF+nuvct1NdG65ivlw4Fyi7UFTXTQlZUAsr4U
FN9xXdsggHY7aof6EI8WiVbCSF4oI/v0ey6U+rZ+KNut7wvvUAMfEfQViO0OJwGm
pEn4mMJWfqcJv6DfPiScY0zh4ZGmrQWbrM7WOHqiif5OISnwjfgy3//zyQLYnUyv
HZLnto3Z1y4sXJm25Wy9K+sni2U8yTjhRzuVIiIyViDnYOgnJfDmc2u8C4F6WOPT
1VNiL3fKaN7lJj3mAc2FuLpu8FlefkQrcAYUHO3Sr/Sg23sdSKBK7fkCwGpzeio0
a9zscVai8lBHtx/7aiHx85QZAmFd+K4OHnCroilVs5678a5cJ+MWNsij1JkrRZQD
Im/6frJw9JhDMzcYSzvuJhl+iJrjf8lWUQvjQvy4GapWGpnRl7JXTnZQ5lD+ilsi
CUBxT6zyaOD5HkMkbPjQ+rWyq1Y6JARpQaomvCZnX9kaJlzVsz0F/97ml4q8aYCN
VslA4UlzPwIOomQrm9fTTqLSr59m4mtQ6KFgCfTmLmFcAkJN3HzOqoP/b059ff21
AyOORlDHSJv0KzNrqhpe/wQyV9sM+n9Unxwzz2f1viSCNuTJ6BGuyuAUmLUfrX8q
ZM2IPX0epJyBgkcmowGZCuGs/xer7TlaV/o0nxlnB0j8AjM1gMi+RcR+E3JRLUlt
AnVyRLRo9RUXi7gaTKRMQ869b7GKbJFzNhDRSe5Xj1owEfyFByYZV2NLy1/QlOZ/
NFKBbIUVEONKluzlcCqKL7miySN82+ty5+unn3mxcuriJ9pRMHOh5jmj6MY1jbWg
uQwk5Txv/CGdHAgfS2w4H+fpEoB6eaC8emyOBXDhqgRz0DLms6QMJ1HB/9cSlO6I
5Iq5+VzvXOg/VG+ZN2521+2EHZzGXbQFFH4rIZ0tlJ9rBGC0Nr6OimasBeNtIxve
RqqOERCE2b6cscPamE9V8uiOeV9NpbI60+gIINWiKZgxU/UY2E8c/KajSAKqO4UN
7IyUCeTxYLVvM4xcNOEzD6sV8GUUfVCRI2+Z2Hsi1pZQlM6JQ325B86PkqgeLPka
VswFlttAdIcba9u11aKKS7w9Ykxso34UVgKagxA1WWa5FDOBsmYqvCYU+iM2YvgQ
QeT0fiWOHGq5kP5cl4N9gAnk6HXvjw365KJ5HZsF8qSAaNQf+mzAEias1NJm2JbQ
eyA3KpYjQSUVkM2IXWVvI95a628jXllhilDojiXg1riu2IBTpBnanc7vutD7q26i
yUoCdZDXKPoHS+mWHCvdN0nP7GebA+DdddcAeyHUz+0FLkFGIqZCpJrIV21oIpJY
mc9jirWjxHu0nwHhCDZQkiUx8N3q7CniTMHjqnhePO9gRmIb+WTUSVsm8ABZFO1N
p2v3VjqTm/28DN+QhsFfcKk/ouUsNcRdnHOCQVpYzvg4+5ySSqRQr3OZc+cKdmyJ
/Xsh28mF2z+D1trnvUa9ne4pOPlFcvU0IYdwSUS3s1E0PwVYMtNXE2hG0OKFL0dg
6taPuBhNsTcz8qOPh2EuX2fBtpvvSygOiKiLP48LrBJU6GzJlxotuHfXhGa5C/v4
PnQZddHEA/h5IGQMc9QTdKb3Ho76HuLKmRn756A+qnfW+06zxWuza7yfLU96tZw6
qUVsTE0EMbFz4e0mjHDmk//LgrHuEPZhDbM9hQxSpRKYEr2Dmf6yeOnYVw4wn4Zz
E7Z5xl4JS+8goyIXYdMcSD0Idh0hERz1vNg1udXBskkaS2GCYXi4bnHTFbOtdQqs
7nqqv9rg1tKPnFemf03U2x2flC6GUHMfZsjPrHq0RO5jLVowN0fPfJsDYL0l5Iw6
FDcUM+JwwGMwlEKEqRyv+hPjzA21t9XvCwDrF5ia7jJoQUzloJzP82VHdLtrVM9p
kMgdLsJc66hgXc+l6ih6vK054ZNSzrYOrTmhNPYo+/ybGCT1OFgZRtieBRM/OMH8
WoaQh0XHTdI/txoP9Zf+lgbvVJPJSBjC/7V8a3F77FzJHpqWW4orsEwn999hu7la
j+i2aKB17g4ekGTrKs9522Dc22jfJiTaF8IkJ4EPKu8cljDNNFmxxrPlX8zTk1bn
Bp5u8eHBkZrZ92cVWJ6KFNFD4ZjMlWNXRs4jSHs9Hs3dljRKI9m3H/c3LC/v6b2T
i3PtdEEHFnLNaoIXCIO9hwqa4t9du22KduFh+iinJdGVvjj5p6SUYBD2aFuTeVJQ
M8cz/fOWefURmFL6/C2fUEQfEQEUaO0GGHNVBpQcF133p95mWO72xA6AN1cR0Sud
INtqZUZ9XbEr/nqu0DBhUwy3fw2tyiOl8Mm2CuXX/GaVd3E3SyRdwlzUeF0AZRm/
D/qYY2rroEJ8uvpbShZbxEJmZWG+Spx7cV9b4v0ePqb/aUku1Sm/MVGz4XrL2Q1v
vvNjnCczHxIf6wpZVqxOP5EvVI21qKHb7cdR7Bf/V68rSGw4hd+0syvScg6LxY3T
pzpAGn5iK8OwTfpr9vPoidAgzHE6fN1l4J66EXPt3xZl2QENx1RvpiDkBKJqks95
co05oRtoSo8TL+8QzFoenrPRqsfZihYwi4xFt3PRY2P5+9o6Dnb1G/dWtiszJd3r
HtlIm3IR2w04IAHc9mSQXSHrQYnioIgTkU1vH/CjTpbi2m3DXUv9PXcQtXyV3Wou
/RvdpLFxgak22i5EWMqs4WO2uZZhcrRudQEhUoGB68UKDdJ+m06JEVQYlezpeF5w
fgI+g95nGuk1eGxwH5Yt3wgA6pJOsereBAOtCAEbeWhxdA/MTvKHlYbQwegz6b0F
VPB4qmm60kjxxOFttdf+jcP6J6nfY1Z9NnmOsyUaTu00+UldTXBQp9c5UXUA9ESU
gJWJT8g9i2/z5rGiX4PdiE3RA2uHSgPqDrtmqfwwTq94aaQMqJS1E5nEP4l3MOKB
e9I4QYvc2edDBaM1tAV6BbGZ7xnPy6EcAch8G8WypLjgDbTdAB9grPsk6hkKQdOl
vhllPTuUygT3w8CunSjQ7awHPBqU+WkyBKtTSC+Hv7+DFemfJ7NraVA58YIUVw9S
JjNxKpCsxmUP4+5Z6sFjiCz8U8e2IkwumDbfrbD9jWmxMPacQdzv2e7KKUD5bYkZ
Fs7NmBK1RM+2im9AK6Z5v+6uOppkyLTUNa83n7x2oa6s7kvOI9jfl78ekJCBSRgr
sxJ78OaZSA/7qpMHH2LZNKrdN0Ofy6/LEI6sAvCln2YHSzF7Vc43yiWKrPaEGmJ7
W8+AYKvwyQb9G7UFeU1gm617JKQ8oS2PDFBmdJ2cMCRqABm6bZmF1lkxOCQ/80mo
FyLO4+892FAtdCOaFaFio4DbwLYTnv7WBGS4kmFxvCEF2n6aThCGDt6aVbusydN0
ma7X/O9bxt7ER7mtuYbsx0K7cB7GNttdhOyeHnhA+qb4G1KAkrqA3VLCejwH5ljB
XqQeI3m2prn+A7zV+wt2UgXxi118WM39998qaIC8vhTyq4v84Qn9pKlvawqUwvRO
wGkWpfKBfDG1kYOrcigCUxr4+7KPwuNqkeYxA/llmHSSYcMz3wkLmCCr+BGesE57
Y3BGoyWn63uNPBk/+JYgB51dkN3QDuV9tZ34t4FIYhJeJkH+wrj9I3h2o7LBwChb
iI3b7upuVOtmmtotGpqspDrfbUG78FxIDxo6bBuyX3bw+gTdY9Y0fysaAK7LUuVb
KHP65MNAlChaemb7AOXTUSkoMBfGX79+x5lJForEG2xm546poz/VhtXz1EobvhxL
whfbX9B44aLZc4CqeTd+uuikkzJCVnAKzJYSPuAY5NEwTIi6zDEkFaBfAvxzMknX
FcLaTu0a/ydoqwEJv2d2M3//as3Rm52OnKN0nUxfukbUh5V2jOsc4qH7XLfikbaX
YmV3mJthqJy0i51nFTEjs8POdNHOIXniwV3SDuhKQ19gqCPINvo9Ib40D4U/IV5t
Wd3RHk0zitw3ulWEXZrno9ZdFmlTqETxKHPiGhwkA2/nRooa/t79FljagsI6Ybcm
0050fHsnQeoCP14sy3rsBICasrs1MYlWuT+XDcGYKuPoUh3x4PkEkdQtcMqGkHAE
rJLidqXN+7bYLx0qwX38eMpNeETozi17UDS1AbwcoNk2gPTArzSMxJrBMCabuHnT
F+Qk/l+2H4vAz+a0toGez1Z7AotjbmfPPnSaOVAjBJnZid+VZKJwLh7slsigZdgN
0AjoKnzGssLr7OCHAdBBapCuXsz81h/L1/Tpse7mASe/2WuycgqFgkt6o2VV1gNG
YZeKe0YlYcgF3Goz+xpE9WMhfzXnc+OKmtmt1YpwLSn+iumysOIYU4gPf/wjm2jA
6LBpz5nl7IugSnktyzd4h60p5Iy3tKA2xG6alrbvgPvlo+rNXZALoWWh4SDnxDS6
jwjyUonQvYeKTOVuqGQQxhOQBO7Dmz1wWRb2lcEIkyUN6MHE5sj6/coIqepPJAnc
UPNurqjAir6NDbGfCpHaMrY3sSfcwggXOjl0TkRTiR809QMs00zQSWks8OxQjqp3
UYSuuFAm/9kf7ZiRJKojKW/gL2IlB9QFhlj3lKBmqtVfeIgNMm7KhoeEFzMCRzcX
1DD18OiiDYi7qJEZqkuOq7dZ/qhS4XT9h8tpdUKY14dcToLCDtG7NBLRlbNJLn2v
ndwOqgZZ25jANfyfgOZkVw4TMYYQn21UHJGlanfMIwpe2vN6Fl/EUPVCKF/1rc7C
TduvFcFXzfI6QpI+sSElRsHk2M726MrWyTxavvT2YFuaLCo2JZD8oeBOE84C731/
edxwUnOElj3AGVoDdar8zN8gjs6IqWe6khLHKwaRL7QfZWgbPLK/27jWmBCjVkZz
QWAbUqEGGXct9CNxok2+NScN3irsqKRtsRmLxyRG16JPP4Imy0JlJFZaCs8rRbwP
S/WW+I+0Hugy4ajAXCx/l25HgNuamlUEVG+FDNfELgmuaT3RS2DF+nxbkZcKk72P
9TK4i6XkQrzKbzXOUtZlsuWplw/CTTXGqORYYx1UbFnhLZmEqyD/ucOg+VADtoB2
s0mPJnhbDijpQ8qRvubKUKYZkXdy491wKWbqv4iY6LEIMw3yA1h14AJvMiLiO/sH
Lo3Hh40GO13dLjKmuI/sarU7Q2CYIIE+3V34AFRWZ3s9cbGqhhH0EWSPCGxdzgd8
WTH4W7eyuQnkcuJM9kvaIDQIgUPYFSjrqhIgisXA4X5et7k/bozYtEzlhFHOQwSe
AwUVcv1O9YuOdlDIYNb+bwDG0SHPBvBw7kJ/D6J5ZvHtDcVAEF5yTTluQGheyoj7
3Y4Xua89/9B1ddiCMNSIqdbhT9Dm/6cdtxjHlzEVgtH+e5WQsQ76bwW9mQhkUyBz
m/gtyaINEcyKLPPzPDsp8OiAOuhnZmlcV2s6Ds0fCJ1K7wGHQv9EbrlxNXT5l7re
6PmMdjB/MRQ8IEvegQyfdCwMBSPFBcB/A0ZPGhYP2vnexLc/xJYUTXqWxKN4Ka/2
1gpxIoTnTm+r6qDgj1NyqwH0gIxvtqNYqlv+w4B1F1Gu28YHjyYL9S38B/PRr0c/
PmUP66Nx4a9FRSo1XKKbw8kcs5KGGDeJgPMy2KnrTE0sJZu7TGctyEPwLQRLcF0A
mE0MT+jy7JX5ZYjKU4q+VGRynWSLLXUe6XgPD/mVFHimifk7UiEe6Es5UwiueSP8
0eynqssB/W61+Wzvnu9K9XqlmKaTiR6AZfPX9Kl+NhQ0t/s9GNIOrc44RDR2g79O
3PnhOFUKetfU3qBsFA/0+1YRm+CA69S8tbkD6ZOF1bv1qrkASKixM3GRCiQdu698
QTXHiiyTRStk89lRWhpA8WGn9ZbE+gg5H/N7/d+hdj7Ut+HZSayU/8oN+lBlskkA
vdXonMvABT4RJtqD4HlRcFp4Ls1g/4kG1bpKO2d8KUZuMN3+p7Yyjxg1X+ygCimW
jeTImF53OPYAbSwgslrDpcp6KoCE6rcLfv6UxpzfVxUA2TA/CxZsJq/EMI2pVoXU
p0gO9Qx5Mpozw6oWTmo1ur1tqyGGYrKTc5Z0I8AZoXB8D9pvLO77X8QSpaNRq4g3
L73+0nPp6Y+oDQ0vhdqrsSlimwsOyJFghDXdVrHOQ+/7uJPNVyaG/nCIwyXBJWnc
avtu9MM6YobQ5UQ+uIaMmbxi2xggAwul844vm5EWwlv7uOIqeGZWLzGKYgyT6dVc
9FlxWyrWbA5p9LrEwkLFS0usVzxaO3LsXE0Iy8w8Z4rvpWs92vvzez7XBOf7de7k
aF0LZXqMURlDhCpiUtvGTIubJUtJkvUvpHoXIXXOX1/6cjbQFD/syR6Adb+aWmiG
lAtfKtNeEGDA5uKhvqx9BsAlf8zYvc0pXGVasCOlzEtmNMHU4sSYtJeNsJkYlKGo
RgqGAcUct1S9qok9MKbBPwUMmVGCofoX9Z0aJKew2qvgM4uQVtZlZSzG7gPH7FWT
r6mjVwFT3ENEv5MkhQW4mPNUyj5dw5D06ChqwzMw0/FxP9xN8iGL7ygKRFiLNwOC
q2VDyKU+ztzXFFpq4iLX2z+BNlMN8T4ANu0H+NC3bY4YCXtYmb04tbD51oC+sAAr
Ren5rbnCwgxsyBythBmKJPP+f00n2OfJtlbFdyTF1YM4gpuIX6PkQ/5AZqeDG/zc
eqPUxet15PZvaTlMABmL3THMV+xh+67QGeOyrS2G6MJIfizYw2Xb6twX6/qrxreS
pR9BD/Uh7++xlv65piQGFHR4FPpIlF8IW0+EBLBqk4P8s6RdXe/5P0DooGXvq/iv
gQ4uAFHjcLtliyPoMyME0+MEForZ/omAVXQoHyHIgqrw4hlhwBgm4v89pAx38Sh5
M28HToBbX1CKKwWJMhsJp0Tr+0VhYW0GglQtj6tjFTiVfKBgo3k/p+vM1Y73edvf
bWUnapVDJlv4iuPKyREu69mqsksFOQNLIvRqfY7OLwmkvmyjQsbxXS0qHcEurRBm
cJLWoikzQwXS15bUSPxPamApHlHCPY+WN3qzqek+mtNGInSJlR72OTYAGOWcdExY
2efdPWCqAHro9U7/K54l+TQTPG/KwWY1u+VvonfUkA1cqdvDHMBYlldjfjadhaKH
JrBdZ/SsLyuZ0mv2Ytk3RGNOQWROczC7NIYrHgNlakDFs5f9+7keGYPulaxA3Fqc
pM7Ew3hgk1t1GcXA8pwoh0JmzNg2w9jwuFMjhmIO+Rl08rfnZFMB94Hq1qKhQIHK
o82pMSV7CRwVzu4Ma//f8mr7PzCTfKcG8F8p1kcvIeivZMDceSeckve7quKj60ek
wxPhikCVJU0mPDOHeUBIMGSV0aGHlsB528TWl4e6kvOTsIui5OfJH9Ig12Xgbrex
Klwa0OlIyCxNFt8N10Gqgfm5RpTLntvGwRnhRbYfxi8tWj8/bylZp0GknI7ZrCeQ
lg6mt0OEvZRbSozKobW4cbsrqXolJGi0srLAT6LVWj/CinbL3hG3ondfcTK5MWt2
f8lmqDEx3RFEeS9V15Y86T8Ne7gKH6KK83fGSuobrdiS/gGWtCodx7BPd2lyjaQY
0dS6iUFCnE1JOsZJoQ+N8eN8XiKcBZCUJcwBfwUlcw5kPv0LlFDHIlMtNIsc5gXD
qiNJS+JNRjB3oiYeklBxx9qw9Sw5BBvBzoqxEHLN8zvst7o9QxcHal/FeBiBgOOt
o2otmSzt/sRvCiVR8qdzfzM1FQeCdqA0Szy8DSEKoTk/vfkHZ56gzrAtzI0izKYz
cP+7foxvm4mSEfGPwdTbiHIcRsJHJvRZOF5YOX6l8kE6TX+OnJXkUXGtoAtMq/kS
wvPd7RePgiVNqPN7pQXwKMBVjxPzmmqrAb1arqaNQVk2pxY/K1dQ7ekBKjwQjSO0
nowSuSmty34RUweNRdYiptdDrMozTgxR0nXoqmGcDL+8JnoyNAYpg3aESGXS462U
KQ9KbYqJOx3jTv8FjrDoQviTvI3ENm9sxiMxjyGqTd0VSjJFiDsn2LVFaS3vQpf+
+bFE0cLW17FnoCR4KaFO5/hcReFS6DlyIfzuNS4iN/XKXTgjGF+zu6eZGm+lY2C5
OsQilD2SjPveQ8B6pOz855OTeRP43EV8GwaFf3mA+D/F4H4bSoR//uoogCudAYrW
Y4+XU7w5MOrBCtyT3cxLhqzJB+4qaoMCM731G/rTc/SasPLZmFkkv8v9gldJXoKc
JCUHawANejQ+v7TDXkWZ6+0AByqC1P+qyyXJgH3mjp+ERWo0FRjoppHR3JaMSOxB
wWINDMajV21IHufwsWsVo2s7wfdfQPiH3wzfHweYyObaZTi3P6uL/pZCN293ynkQ
WLSC5DWfXNdfFgxPJet0gUGwBf97ac7ivvFVImrIojl2dAPsrxV2bq3ONa51zPZd
1BQvvczR7rucd0Pk6a2/db1hj0fpl7GUkM7a0c2QZqd8qI+heo9TjoR5o5saiOtf
49+M5nU4IRrJhW98hCz8R8OU8TjVHZzWccbEHg6nQzbJV26UCa1QYaNdgo00Lztb
lRhY42F21Dvoqoh2Tgizo4jVAD5opHIgR6ZM4Q53M08w+z1+CfziIqSmvaKX2VHD
VUmBA9bZOOZFLggSCMxon6xlMWVwcZPMu7Z8WP/cifLAZufkQXGmFfdfuJLDCn24
fh5V9Qj2Ui0Zx+YVHYKRynK1lB7dpuR1+SzZ2qU7QYo/UlsfZ9jScPOc8kEGm1Tl
xQH7F1euJEJ6gE8H4fP1uf0kNKhugxx6XsZXGgDRoy4PfAhIfI7KhuYVFBUqaKxY
VnAfxFytHGRl2axMTSs4OtE8dly6FEPJ/m/jzWNKftAF7A3RGgYy4Z7r/e6/8HJV
HWHFUhCRbZV3fRD4ZZCjKOWvROKay9b4yLcZEN7eCLgU9UgZ7XVe46jf40AW9c6d
ES/SHo466ywNmn3j02JpxHRiVma5ScqiC1UVOhWE1114xrhBJ4yq9b9w0fQ7LWaE
8aIOPMkDsBB8RCzxmhqdwNnjFtj8XtROHgDn8NIC/J7QlJH2yMLVd2lMCuVYF/qz
0fDftod59od3eiAM/mZPgcigLdj3mDkJMNhff6lSklX7ZlxeIjh+mcywiytctoR7
gFsV+21rxyXEGj421k/qGMhvDQFzAE2prkUcjs1yJzuKbQwyvTr+FtOv3VKAYJsR
UuqMPic/q186HwDjAJisGvRcOtzaEhCZ253MPjHxxq9SJTdqrBSYbjA/oSC7Vhyg
wWB3Z3j8CZBJqgzJ1r2egy+jSFo1oBfYc5TWa52z151WC66cbqj/kv4Yt7xDrj9W
4WcXyBXNNCkaOou9zub/uw==
`pragma protect end_protected
