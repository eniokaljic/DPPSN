// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Fgvn+KyhfbLDX+r9FstlKVl0DDY0twiIe1IG+CvVWW9ekGYbakZfDbobd9FvNimI
9jd86oZNt4mgWDuDmmfNvFiyn04gkkomXPH8QygojTPOKb8uNoJ6MeI2i/fXsMmK
vY9Flz4sbzQCgbEVOw1q1Mq7nkfKW93YrP6DfQPpvW4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32400)
h6DNVCj0WWQhprjYl5cgp2SSoS6pALqq+7nnSJTQRY+QvFmziJVWT1hpGWAfXZE0
EH4ITQq6n6VwOJ1g45DLuCnhlTten17Eg7gaAy9g4RcChHtqC4wikc6ycbJ0tkDA
0AGdkKMdM9qzqy7WdOvoUkGIVKbBmzNF5l40ibaObIN65wSoYMpiegMp1cotRSYp
LjKn3mvvkD5lPmey+4xnZY7AQgZjMa/vtt3TIjYVfbYv+IwkJfq7R/bSC4EB0ujH
8KrVExwgroGAMaMererPXj8F0BEe0ALTWzAXqxrOi0FxlLLfx9Enr6SMecMTojZo
uzl4P4SJmvSfzczjv2qgz3Lj6iWbNcyqQ3RVyPkbgHJS7kzzINXAOZ3E+53mtc0X
wsi9Q7Fv19r3VwPu0KxN3peL3xQubuj4lq1yjEWcSkbbyJddT7+qTQwE+1H/oO8q
O82P/Fsq8cp0EmJgyjbP4qxNqlo11OVx7h2qr9mV4SVYlTRY1VcYpG6RqmTBFUKL
/Wd4cnEiV4KkFdqCUFxAvqOu9yvkyip5RQIWVKmF4ODzZsJLCQTIkij2/zxoxH3A
6ig0OaAuXRlz57Nul+4Qm2+YjNQ/6/2yOFb6VCqZ4Cu+Ag/7+31YLYFEW0Fk7JT7
UyjWkzb8ps2B2jafOxEe4goGGzTJZOwU8b85suRXVJyzJSYaVbcOmJgQkQq1eU14
70/dM64wEIxMjtd8uR/uB4pPwU2yNbe7R33nkQwVKJLJa/TsIxAaUXvCM3I8UoXL
PoRF8zMoLJzfuAah4YPFmEal+yAiH63gc9FwuWSafOQbwuzlw1eX++R4Yg4QdqEv
K0coSHF63VUXZReyqKJwm3U+xXgii6WhfDyIxKW7kUA+8YWdZ/yMkZGLKLwIXtQP
hdtIMWoRAYru4lDWLWuXi92yHMsn/lpmppLY072AcGB0RGh0DJxX3PmRYbJ/NObK
w2/HSFdC3Ajl0BKvkWzPfbCeig9MHMKd8xkuROEEw0iGoXJ27Tv2PkMwTfosxCJC
N586l3iYHGcrjc1hhJ0eeA3FoVrcY3aXlH9+I498+bGnrVzXTI8PHcCH1+3XgxcM
jI1wm3VWRm4K3vZ68q+I8BYHqKXrCDWBJGZEtOm0oo84gCI/Lhoywf9diC+JYBr7
5Gu4TZ5hoPlWzKzxZv3zmLuW+xdM+uSKqtXxGINLSH6nGvRmqfJnRaRN0WQoEXX0
x4Ywqko+93zEG/9/b/D/CsCSNSHun7bcifQGwHXFSeGJW4KMloUnY8JJi77aLqa5
9FhLEFRKetGMOU7lqA3+DfRXeypx98FwebSVi1DoS3AKnqmrCpbr0M/mUXppHg6N
7yKL2xForL6VQ2Qs8B3rvUU46f7sfEPBiYQQL3UEiYEqyNzWUCzMO7SltJYeenOL
eCZ5DnFhDRE+7aaIWfgAAKBDBvv5DHHilExMzoi1maCUEFCec7PqYokJnWP7WOpO
B2KJ5EGz+SczZBLVtkGDc1c7zpZWI652imTd5AIuKHepxGHn2VzFnZF9kFujZdRb
aD3VufLi2HyMvtLnLtG5GmnJGplcsGD5hw7YTUm2gQEZ37hhlt5b3rkiLlLZlRfO
BHTyn5XJp8/GVz8ku54BBTPS1elnuCaKMNR0IYsN3ts7aay5aagmYu45AkrGXNJQ
38yph/Lsh7WeNpHONvuACqx50eID9BnwcpRAGaWmlgTxmWr17IMoXqzgjwtzOPuQ
spkS8ZkwcCY3pl+3yqtOG4p+XVWo63oftQVt/KUxjesab9717l/dJlAJj2/QO3EI
PzF8vFi6VvD/ghd2HZNo7ISbmYt9rhO5LoJXy1Znk3+l7gFemi0QgEHyLtKWQpud
W312BeEj4rLNv+Q24Mq6OOwVH19e73IuTjP922kO6yqWF5PqJSltKgoiuXKNI94w
676jilzB0hN4xk0lLZepFrQuYL5f1MZO0WwN2GhnyACO7sEAslHkBURNciOOq6mb
+RmthXr5YWRReWDt1prt4qouQeJyMaiJRTgRd0Xz+0pvl4FLbNQ+N0tnALuOnt/z
wOo85POzzjZIdryW5ijDLCjg+xhrTvTs9BU7qE0jfRhsX1X5f1H7FNJwb+YCW8fP
OqoE6H07AufFv94UNaTtcU3vJmSWiNEYGGVzZyAraM7zngucFO4AKzmOlkK7zisS
Iuch3s+vRPx1hlZGdKQaqH0olJk94YGEoZzP8LoijbXycUg2cdIT4HN92qlSFFDP
fT2BLrU3uQwa5vSWZiuDhRx9J7Dh6jkdoGesUpm4NJSJvqjbQ6/LsCNnCYAsNnyq
O84sIDySTme5TSwdGrkG9rY8AHqqNQ2VmjQqz8fl3JZUc9G6tOQecVhYhp2frS+W
DM/hU0bFbrMiiTnAL/g/h8UdQYWqPgsOerYbW8y1zPR6xsSeG3ltOvpvSELI/Goz
wnkY2acb8zxcKXKUgBzzWOV1LTjaNkp6XdbAqXcHJsThQv2toDlhZw6rS2IAIfEY
1K0oTvCXyRLlaWFoZRaNUcfaRpKSXjdbIlXRZrFw4EvyU+fe0LR75CjZ08/1qRIk
u2Hmr122EGl8XzEV/b9OPKLIdu95oA4Fujdfk6Z9HkeC20ScLPHb8bxchopZutO6
GKNfCQ59/H/V2WDxqZJoCCM2U1nNPHHjE3N6wYn9k2+3HJ/jHztLVOy8dmuYhuAN
HQ/Fc+RwVzds4tfbZP8M7Zu1KTrdCPehvisLXn6VPO9yjIcnqDhJI77oIy8XrKdl
ey0rMjM4nDXnqbgD4tofKcdXgjbf8z7a4BBXG1ZNozzcXP2yvA2m/pmCiV33YOib
HDwr7T2sO0pRGYrNMuc2vNeA5JmzoTnzm45eH2OzEBGsQasp5mbdv/CG4o5R9CRh
vTzmBLVBERINN4FL7gvxWWfgeQrwy9S7gb+UoF7X/o2kUlXInphNVFEb9/JQlrP7
28qAwLv5KArzv3WzPOWZMt1LR0bxgnGGIKBZdNCOIJHblKKyzUPf2Xw+ippEdjLQ
mZu3fSgWtgRFUiM/JI3rTnHTzG5NECVTmaXVeHOjwtOkMEVzba2q/CrQqwP8CCrU
xOIDB4XJ2eZusaHS6DuyltDbuy9qc52Cjbe3gRXcwxsvlCCKLWyH/L78LvUfmjyb
EqQkAlhJOujHjG54+mMW+UsbwylYSnkfZ2a2mhuqC7gfXvuDmZ+/x7aWtRcv16nU
P9IiqQUNSt8FGlj9LnSyzBUQyhwJ/2Oq9dHfBs1XnA7+kx1iMjmK62m+EKts/IGj
e5dkkUTeiTQZlMCQPhePWtVb/xkgq2bZuXNGEkBiTkB64nN4pbowyzKxFKqsBeOd
mKr5rvHnBv2DHaim4yUaFkF2WcB1Z/iyQP0F1yzbnKvRiOfobV6DTOQ4FCW2fZzk
nsaoIP7Pos7vZbJIDtSI1GXm+8nBqBjYdWBvLQ/r5WQMCSXMb4JRNiGVEeUGlWSq
1MKw+n0up6DLV9kjpw56ESVpEPDBA8qVB0cFc0k0w7WxoPMXs1BLV9To8dNP+k5L
91Zj4hl9/g/sphCXwD0WiBxo79T6ZjAS6ZFtfiSMT8/vP208vBw0UeO1dzKU3txf
JM5U65Kewlz+LgiLwcT2a7ecPq+74MpeulSDy8pSckUoC0pjbh1TFNNQFA3B9FeQ
tMcSBMM7KO0TwVmHxG+fv2W3upN7LkyA9MQlVfyGPxdCbJxSdRg3NF7mFlrhaDmH
PrJxJmGhaLv0iCZcyR8Z0zp5g6CQGJYuciuRXQdXycOmdCCMu4NOLlRdc7aALqEF
ChRXbitvsjjox1AGTFn7j61Om0sAwBldxWsz/b8jEsQzhv7UeRbTXeGPmxB11Rb6
GQ/SuaRiOQMBe1eqa5FpHiagy1EqR1sJn1gC7ZrZVjLVo/Evwr4JE55qmvcdshUe
3W9/7LQXazmhoVH4eZbOFByGA0ioM+ulaXZwZERibmYw8FbQ3uvOXV6rij2XEup1
oDgmhWFVBl1hWLY984gyh176UHkQU0ySW3kZrxBaFWfB3AXHRZRojVyjuaUnXwxF
RMn4HQdhrcRLxKQ5RYa4XdGBktsQWnsO7uKFvS+4O3k1QbAUexx9uFxDlvuhxWVl
vfPMJKq/DjXdHSeGxtFqF+kRx309r3OjjRDsjGEnO1Wy/zLXQBzZ2bbYv0WlmIie
yI+yA/pbdNeJQ6Sd8Taw2/N5+e5pjarX70eyWeZrQ0RSrwShHO/gvmmX8QQK6+uC
tFfXVQCqO+BA5aYygUh1nWsfSQgliqbugvqpCUtovsraZjdu9aCV7yuN/yjbJ09X
S3mFexnsT58l88Z9RSV/SwRZkqf/U/emrsZGiUtq/K5S9LKQi/2JH1L1LYCeI8fm
FLt02jPJI88C6Lxi1IL+hr626CjBciKNNBd8lNwVX2D3NzBDaLBiz/3Ky1+lwmQR
tzaTq0jkJDMU6yFp6r6a3VIt/Mg4HmSjvYSqBMtYwnE/BbNrSXuMxGa3qS2gf9om
ynYRxKDhKqURNi5TmcU182VotLJvGjrrPGie7kP/0nuAv0butbp41RgyschE7IHc
EP5cMHpSXwhFzWtDjmmTl9Bw4gvi7gPI7Uhk8JAe2Z8tEUsJsxnd6pdoW0z+iVdA
Sk/+d9XNwfWmnADYLCYkYUtDI1kHt6MTbjyBsq8YcdmTdW2OCfvBVduS9Z02rkcW
PIVeOQWGE9KoEyXV4jHGcHOnNA1X11IBvbuTcKnGghOID42VBFVh6gQgNQvjFAum
8SA8GKa+wGTn+dOYVS+j/ZTlMXT06kkCKlVTwubznDcfw9U0xJ3CCkxUAFC8ATky
9BngKQ9Kn3UM3WK1sIx8cg6K3b+RAY+Ce3yXOGhUvTO4jDup+KDbxV6Z2hokJ/BZ
jlosnrEBZbrTstfBEDbpAcUgxXCW77j0sXemeAMxWDSiAsM23Np81z2SzzeKPRsL
GMjICMbnJ9ceOJrs9YSu4NiS9pv6656uCczV5Sbd/D3vxsM6KsKzXXwlf8zMBWP7
60+2fIjPQk2iN39C8z6ykAF0AeJZKbOT9hSRq4CtmfbKEJMhKpQoYCt2CHoE67Yf
6zRtPut12Oet+PBwTqfARfL6zR9aTGsLlQgqmip1bffL6JrTOYkFCGmh74jiGh0f
JH+d5xIr3WqBUjzTcRN/zqm2Km8a+TQyLgZeUo1pI0rKxCdYNoHkQalR6UiYfdtL
80pPUStAhHhseacvVXopPD/+UuWBWLRrbKGqlOJHVY8dDDDtIIIS77WcOKTovoD4
r4jCnk3sGS9zV478ogKlLA+COCy4M2FFeUVNt+HRQKh+eBoiKdiEc7tr0gdu0v6v
OvwinSc9S22UTenWTzzCZV4NGPZkNgbzBuSWP3GdiD1y3RmZTvfEZ7sOUO8Kl6sr
atQfYR3GcdOWZqa/d+gpgjFDzUAKJCXzV37YGBUn8+kb/6/NZkP9MD6wwBETaIMh
9qEne7qSYr5bffL/iHVFizaOgcl4d/Fhjjn836+B4U7oZbZ43+jZSXQTAcjJO5U9
MY01gbr9UMeJvxlOfgrLuey+5qBo9h6L9osofFOH3PJcT8ZejOGGPMeup6R5J6Ah
ZeyMdxg5qpglwgbxvjjWbn0vuyy9y2xXjkI/H1nu3od8ZyWlCSugAYB2+YUb96JU
wO4j2R2zZtu5IvZWTLUECyuhpR7XVdHbdF490WUhmf209tIR+e4ZhCPQoC6rgYWo
ttuqS11clO5ScsvTLP9AvFnvec8vnLPBUzEhKFo7iA1li22h5GLDNw176jons0q/
6P2YY454tkUqWS7A2f64uPX4giXWdCzfOkL67ur+zRstJibV798g4C6cxZA+jkND
iScMpS7reAdUOwgkevrUv8kaBDOZsGtAJdPVeulrujIoEoXs65MzP0w2f3kerkPp
Nq53IRC1LpMaQclMeg45EWk88Um+0YNBjbpDVBj7guLA1Rx8nwrXEjHIxyush4Dw
7GU0LeJSzpK0QuS1GGsvygAZ6EEUCer8UHPi2tO5pdUTSTHDRjww1knEqTKKoa0f
75VjFqjqGME0dXXr/EvdlUjFOyMJoTwNwpe/am0RJwgxMda6pTRUe7jrRPcOIMjN
87cRb2h1+5Xf9GMJJxcWiE82UJdajtEsdt+TRBfj7nYFc+4IH9L+StD/Tr+myXud
78BgtCk0iW7liQJzHjNqB/0bkSlWy2ljF9SYKQxjjgPybxFTVZUXb0MdtVHilZtG
i5Luut4aW4Q7TOttuwfjRHrLC+qo/fTSMUUGEDaTzz5pxnC3g+8rK3fvufHtCaDM
fo2e/+XCMjsFAi9IaiFsD8MWydG/MGQqO2FZm9ixEXuuzBXzScmE/R5AOtqEQ91c
qACvPkUntwPpjwMNJ5ubw8MB/zXuvf9dRknbdyBMSH/1Zp/f0nwbqo1myu/dWxy+
WQA9QLKb0fXhGZwx8iN5dSNVNwCA78p3dzhbBkCiKK3FcNWBwoOaaW3VQ/PVxMWp
dW3EOsmDDm4S5JO35ydFUJZUXUw02ZWP8yo0wa3/shtMFXyXdRyzwJC4pik7oCIO
KzuulKNUqmjGdwFRgKm8hODV5w3xik+w4J58rs3eLvJ3L8ZITs3FcGtc57LdtDUP
V0vKVVm6Lhy1nDDk1yn/NuxecSvAO580Oyn+HVzGBRb3Z3quwzjWwUfoD8TCk6+U
kj17Nj7QHhsA6sEAWcNkEAPcOEX0aiP5Vu/uIyQTGwP1OYGzzhuxgp1PMnuQwFtA
3n9F7dHORhs1jax5lbvS9HQ2v/GD2W+Q988+DY2JaxyvQg3oeU2i3IcxtG28dHTQ
M/bXMFTwbQt3QNxTvcX31edB9odfW1Rd5TWSGN2aHc60dDeg6Fc7tXhRWX3rAzem
5fw7NpvYIGd0CroIjiGtOdvbjg8faLIpnY4cEoF7xVe+TqhwOTCgIKl9i2K8FCM1
7o4FgifWcTo1gshIEvAGog19sIpEP0uk1A7nWF+L7ehxMGVdNXFbxyuL7m5VD1kk
RvPkJcHzTSFC/AvmKk33IngZrWHR36RFK+pr7gDFWyeIdm2bwzyPixr6ZB1Muvhp
/DLiav5AmvuPiyIehdTf6wRyz2bD/0bfkwqgl30aBaC5K6Z7fVC6MuAuN3E0SdFL
qGCYDzVTYbNDAbbAhehK4UKHS58ucLPYyX29vcq4tDMBEFeHeJk3KeJ5LrLYytRs
FdfO9yiK0VU2rJsrH8wtub/a8OCyFCZA265SIteY5yWdfHqILAYEPxFOporza7AC
aA4mBad8MZo26K0iJ1HSfzW3cKO8XOVtM2Af5B1oW8mZuwWw2pZIuzgRkXdR6KCM
+7woKWeCVoPh5qVTVk93QKmfDobaPNXO7GuTaMlDcm3yzwzjDtkab0gNd1vD30nB
DATg+Qit4vUsSjlY/hUGm0UEQbw77GlyV3FvndvwDC/iLtZnVpW/964bXJySBWSZ
xShmAd9qforwwyQ4MJJ1A9dayVQfE5z+sHrX9Uhcr3onMo04rN9dp/UQsA9PcFju
C1aGaJOHN/F/TZ5kORZOQaG8bqlFROukItcFnscKt8YdoEVp3ARgThmXxQ3+dJ0q
AOyeGWsjvPS96CW5I+oFLVX0px8GP5fPw1qiDUffMJN0c1DghpuxmjK+R6Ty646U
Tz6Evl/FSPoLfFCyyL2+2TmtwXaK4JMxhVhbLaaMYVSdhuTQ1Kp5J+phhVoSUgDL
ybM91sqvSNiwjJ/egGT85CGwsaGYHut0w17VRdZmVwwdlT9eXTqy576rinDe9/3c
b7UtBZACD66HQvxS6MXZg75v/KcFIDGfkuclJ5wyVNc3yQ2qpAqB+s4AOfAmspcK
ABM1NVpjiXq25ojo5jBB1FJttSea9+Q+HkxJui3jOlNgYS0JOl6yRh2xBQqYS+wM
OgUo43AO/aUcWFzer9qsuByJ2WfPl8uoErljmTIIyU/M8HCf5fXSt5TPwer5RyAW
Aj/LS5qAgaTrUsHsmLVEZSd3zKoHxWj9m7e4QUcyN1e6CyLQ6HePQb1Ir+kA2TaC
oMYh9qNqayRVMsVy/25J766/v0RB5nXtvJR0r2bcpOtuHvsnGn+gTjAj64te0PfF
bbByUVVSzTXiYXPBnooodVIq99NdwoQTHN+AyLpzK2Lih8CvDCE+YkYgwlOy7Ghz
LdZhVhuT0CdAZhX1YwSvTJJNZtFmruAF+kFSLvDI7xl1huC/KyixrO9yJzJopkou
nrcppkDmS9YAQA5g+cin5x5ogaMgyheI+sTZ9j2nBwtKi7oFBatgMnQSO7DXLgD6
nwrdF2qgf4+MD0YFJQc0cZN3D8ATsJlU/eGMSQu2cLGACErL61OM5F40mdkJMRBx
M335cMuSjKYV0ggHWtdW+ojbwlCQJlBQ+tPaD83340iFU/LwEXj7e9Fv0RTyOpyR
n8MQeObpf7VMF4u46LYLA9BiGMFEciTu2ivtLUsxWyRKuzEmWS0u8R0FHrWqvimp
dVqL0oOGP/+aSpBZCPDeIGBpHPKnAIucMn/ahUhuADaJmFMplaOfIx3F8iB3Tic6
EA22iS9vbl5jTHtshjUxIaMDZf9QMfzLE5S6F8YimBKr8Y9Pf/GuP+CcSTqsEoGf
eD+mO9BeUkUuqZ3gunoAcEz1N0KtWg5Dj5FrSCHexbOrUlW1myMEqGcw4U8qH81M
mVR61JqlJt1RnrUiB0FHmY1eBaBEgH5snpWdSc5ze0uO78CaeMpYpPdB189FiOmP
iOyQ/M3P2JfPEWtkwFQEgMiEnuYMz6EgmfkncEl4zrJpbIe8xBlX9jyDWE0c4Giv
aewTuZFL7mRqjZJW+ipAkzeuaK5SounJpP9xeYLtqwhRQ398lQZcY8TpxHl60gkh
oLzEryU0CC/rf0uFAKO8ajcwyBQNNxItydYl+IGLuRd5RrdvnhAkFZWzlIV1xCO2
n5k1FmxVt+zbcld8D/bcLJT1CYt9kXEYPxOO3mM9++8i6Arp4Rck5nZa3Xo0WijL
2zOXmt4mj4e9EUUe8ViId+kgE/A19S3Dv1TKicceCKdC9jAWguCB1sf4WyiZqhqs
Hbln4oqLM0fkfuXoUAdpbXEmbBrlvpCdQ6b8ICeI8G9UpG30/fu8zCgfE0Y0uJ48
XNfF7zqqWyLIs3WtjfFCzvVqgINAD6zHys9VpP3THGPgkLfaBQssrB6mWGrkWAzO
eig7m4e/7ibizGCB2hWlQRcU/C0kP7E9BSVw+oSkkiJbOi1qPNGMDpbOdCulfKBd
Lvv0dIASb5tk/MbiPwHaqvwjTPAJmwULuQZH4vNI8VpCAWPPqlX0BZ1PeqysGNuw
gbDGPPOAePHLQT/9jSwzwRlk2KlZoSa6yyupWqigD1uS0YcWN63z5ZPXop0AjP+k
LGx/Vhk/fMRYOUVsxI1W8koT1k8IWujukLjFakID/UCdzNBnJceLiV9GSs3dOWb2
NG/fdv4jD1d/VhtORsdSLiqI2eWj8IdSZxfHGIIuRqTS1PZSMsP/UXdctlQWLlm6
NrlMwzuG1W4oVdcHainNrm9nWy8W7PPuOkFsGKXVobDtl67q+kcGvExhaz8oK47F
2B4GNPYIIgjd6UJZwILbc44FD3pMUD3e4eJHLUEp+a0n3UQN+YOt1VQe4FyUaNGV
6Sez+eaz9gnoWejQocMxoFoT3gaMfLZS01dxBl2qdFeH2g1qd9yonqSP6CleM82r
Q6QWxIpe9SLFNiZSXRv5lFUGMkIsc5rggSFE6nDeE7zgNPLhytfvpNedRtiGn/5c
yRIhRm/WytvM1JLc1ml1OVe3VumwAH1/TiHvEYKmQLjDy0qtgoZV6eE+oPUT2mi0
Ul7pKhyHvQxFSv/zs14OVQCFJVSRYoWtSAdgBsjfBzgllrRgC8ToBaEJoqsSnXzD
kL5fiveimOTLB8S8mC+00HG7lZgGg9RLJyAtwYS3ZoyVPN9Lz6VfpoaCAThrGvlf
cZGiCpXE281IpzzqywvwlYWoEub1vD4VWeoxxXR3Z+RylCufdu1+Egr9UScIuvgd
YlUdovEZS57BXST0RbfBD/bDttnCDo1GHJYfaaDESx73oJWqlCCfYJq50ur/14M3
LiL/qA34/7ydqNw8eJatM2rrB//6xGxTsjr/ZCdIuuSDo/MMDCa68HiW7M9KeI/4
rtv0IoLYs7ldHW7ZqxxOUTVZgTUymKzFGywA9pV3XepoqcrVFPjhkZ1msuHGvbEP
HnsIDlh/lj9TJBrlX78wCvex5hbkajljPIOCRtgR9pNCBIXRaY9OCm8aCcNLUYqT
Z9HSVZHYvivqcdp92kPhJ8W5m4hhwwTyOcPg4HWyBXySpD6dfqYYoqaTVLGP8Hg5
3TftT1/udWSgChb/sH6M2ado7O5ALQdob//Qk9/M2dgJ1qeqhTF8AvUx6POKX727
4SD5FnGT5ek2IP4pTcg1KtZUV/bQJmBn+jvkX2jLHJ90pVA7Sr3+VGfdnmTeA01O
8VKs1VNZUB3GVh2fTlHVRyE9MkTozlfDSFEh0uu1rzURq8s1ekXpnmFzAzaQMQQ0
ZgcygqR+7D67G1hg0K9NcQD+L0iPe7gBRn8sONcGCDGfYa87ady3TIR32ktTWkDp
YvlM4dBCV9Lc3WIQrg81Atgbe0HzFJX7kOmkgf3sFaT1yCbAAAlMsqfNopg1/l6v
3R+CYkA+pUjHLT3cPYa4QbnpMi8E0E9Rii3Fb7cVUVt/3cc3pHSOcJ+wsXYf9hGi
rgQ/153Bx+dTS2S/hiKszj+9fhPgZoNkLKWzLtl2P0BTVRZU5p+avUhEjBNEsEwX
l6FPjVeLXBlgUNYPtI5iU5YUolL/YsWD2QoExjrFDxRxsl4IFSvW6AWBBbN0+rUi
r4koE+qh5NDxR/n1SfM9oIDA1PYQ8EiYSe24qIg5bif+MTtd+uN+VPwDmaoa/TXe
r0UjnvSff6YTR11yd6R3rx50FH+Nsbc8MBpk8lZ3j87ywBuN50fyVMQ0WwRoZ3MT
xAe1KmAHgGPe31l2I33ovvlwjiSzrxkzK7glvjxN3P9Q4fpN7Zvpc4XIJhVsdi1P
e52eoYLxeWOdwJGebRej8MdsyePbzEi5MJmJ4tQGTgJJnW/EC9u8Dse7XZZ7+lQ9
GxDxqRvqAKUclYtSBmqxTkg1i9FJFzVA5a+tb0W5QdIMJrJoKHiT6JTfRQ5SRPF/
xmrxWh8BOZB0vrLeFj1tPFVNq2rM4NQ7podd1UXvtM20HpY9CINDA/pORELZk2po
Nfc4FQs7lOojNNlm3OVharq6b6kf4atpccfQN3aTFfhH//Qx6+6Ts0ybRYWxsTMi
0kqWogt9G2LIsiB0/vaiX6MrxMwJ2VAxjEv5la3o8f02GdyngmQWSjV3HFGjpfTH
3t2/wavGsaQ8IL655d04zx8m6K/bL1VoYKsEbYRys17TNR1QpBcN069Az8wPcyN4
8xvuVDb4jgH87e585azT4hYN+/PNYj4YxNfQwMy5TMNDH2t96TU/nfy8CFw84Nm0
RJD6dWp3rw2A8W6vvReABhGdVMXOuYs2BKepEzTbewQwMaHMDHHWVqguLVEyCNEe
4MTXco917vQUHTxrIV3YZ9wWt18+RY8sZcf7dYUyFFFkcOhwyC6iDI6KEMBRxDZj
5jTgO8FfYNQbq3uwiESuU0FMw0EWuGyqCVuyvYeRb7HuWsSxOPAtJlsurL1gJIcA
8kfr6kW4f4TR8AqxBWEhbb4vyssQKCSK/FVOIrr4IJasnrDqND7goioq8Ai/gR6E
IgP0vdb6r2eT9cgffNOdA+ASA5rFsBiyiP+3G8tuksH+pcNZv3nN7dWsybYUe8bd
10MT/pxdSxZT0DEwcB4CVEdAfra+0gKRuAWHn7lgJmBIqorhI6RhX9NFFkuMnlUD
SDuTDQqzrP+VLWOqO6oNroxMmiC5UPXMWZ6tZuIWAe4BvtZkmLUXHrqwUHqMOEcz
vWnPbEJBR4V/GO12GqbCgXt6t/VtTEGKwpUcKOYyn0KY67sON4DuM74z9gAm2PDH
lm4fYDWw2c359b29z2ckJd8ABTRkZZHuyHx6wccWiap1NklaGWGKakm5yUwQ5AUf
eeIMaTA7mAnqr35MQwQV91gJib/2hib+LjcINVCkzJjZtPdpnROTD0ifMc3MPM8D
DX9KGIurvO/fUpIKag41uDfk2w2/aSjSDzYpxHlMmwzWmnGxSHKtTweA/CSRStiQ
iv7nuidMt+98sjIq2vpctu1uRZ8uB18ofCeCRiUf5ThoYk8+6/5SSOSisYD04RvV
8lYcYxBt1V665w233IQbkZh8WF74tFU5xwBM8Oi+MgBsJnLSuGwGVFwyA4szt+Pl
ctQyu49L1N0LG/mA2r1mGl1rA/GbYgOPn/c2rLJLnJR12V5TZ8V4m+fYDoOREVAR
G3r79BhLIWcc7GMiAG9BR08iiVpvPf9jo4xrsUazK9g9QxUf2adFLg4TJxVx57gv
LxpS6K4vGkL85/R+Ln+OfBtDHzzjQ1vyQeEBbimzNljURLCVVnFlKlVVAliNZUVv
iOGt8rH7yNxR+SgygbYVFIeJXT58naLiBr4aWkDuiELZfmX4PvRYEZ5GJ+L6EGje
ZpTI/b/jftBk5mRbHdIPrhOE9ADDowEdrrZMZ4B5vbKjXBPe5YXXx1UErWMI5S0w
21oAyVzk5mY25Kj5cRs7qg8qf//KqywSejg4vu4/9A02a8IWjaI6uk/sIju8t57j
CDeH8dQl7Zmbdq2DjOZZBw5Pz3Rb9YZ+0WCYpfu1ylZbHP0+11SL7EP3P+t+XSDL
bwwkLQiJth6SI0Qj0+aZLVIWodSWFV/VR6LXlD25YNIIiEtZ5jDPwfqZJJyhfpJB
6w8wFYETI8S5qQrj+Ut1OPMuXr7WWW9ljL/yYXa3mEzMZcHhsGGK3xvnsKfE8VxU
MxlEzIObwB4UnYVXmPNaa4bDOnCfwcJ4gjwcOaNrS2j7CMPi0XCMFzGEToU/VIUk
HMo/FGTuPAXI7futGw+nempneywYDPoX0bT7UOonL//c4zK5S/jmwaQPNOTW06sz
h5BOnP77VUuUj7XzoCk33DqV+ocQZBX94fUwKydtjaefM4raFjIlI/IhL707Lhac
Rv36vu4x9SKhRKa0+3lntADKvXHPkHvBV2wIys1rXtj9qiytKEotB+shx7uSInjl
ObzJFlkSoaxnAWXmewWqW0QuZ2wIAT47Xqi65YlsBlmzC34BiTCKKR+I5RMdZGNC
yARNzlic90cktJO0ckuSFOhCIWs7jtjJx+EQSrjqnqMwCcWISZL+LxwWW8i4W7mB
HPHuHXnxK940b9yKanPBax24OGgi9TU7zHUK8IAHVacysReZE0D6P83RwpGF+ZTp
H5IRIlxalr8uxHSpOE5wTk2hLjycyutrcR5WLu0hvE74xUmZ4xHEdQPoWLOERlmd
27LyWbPrKkB19emtBe4ZId5pBI8CsVakULCZ+q+CoCPku32ftghcCrySL58eLGxF
oskOoEzij4siNOoYrDw9jP4Nq8Q356/blVS8INhPxiywBLTTwW7wmVirRpNkfOhn
+bSoR1aMdf/uDBx0AhgvTdSpTrhVZVjBlpJ2d5ccViCr+Yf7IIRE8tV95i1QMDCX
0YyKKiWsYY22dkqO/Pf+hmDv5ziXTTzf2GlG7mge6XR/l68PTho+kHB7iTb05eV4
pUZs0X7I6FLm5BkqhlGpmU0H1eaA2HdGS2wsZfWxm/jVxrnGRH35chhhHRK6O040
YW6112tlEz9SQEtiGa2oUmL7p0s1odzOay5IjUQAKjNfjZrHWMrC+rI1y19oG4sZ
MirBi6bKQGGP1Ox4z+sZxHr/Gi3Uuca4wFaU3yV/e7NeTMJ9D8WiH2JGNdnUNV++
LtTxOaQVY9IC74sd83UA+as8kVXZf0PankTYN6oBY/fnMCcMhvVlBkK6TTaFNJSh
1QLBBcUrm9rYrGLDELujZjrwtm7HzcNu4TEyKoB8uiIA2+dYtqUsrXCXA64Q77Yx
cYy04BcxF2gzs4+R4USTYcq2jLtsthSrOWkFNMpx4ipH6Pr8G4gD/ePmyxaH752X
Ro3xycPPLZNBy3hzhe6IUwDm6hXfCdwzAFewxyuFhd4hxFK6kQPr/Rhd4i4PHsyo
D7wegaS1FaCD7QUeRfjyIm3H3Tg6G1jlGT79v+43H4wFc/uyuVV3YI5R+3G7jrqn
gJbGAuRcOxwG/dJFeWaYVUOJRA/l19mQ7TLVgOlZrP2cEGqpPQ+TaGT2esPWHOd0
0ESWZFmZuFd82mnLt3LB9MOxbrzV4tLWfipsfwDUX7zRAps38TcXklfy/Y23SWSA
Qg06/jchxTCjSZLdqC6xLp8ggykwSdoYh7ZSbjujRB0KajlYMRk51bQuEAhZ5CQX
0imOfagQYrZ821mcVmFcd2J5Lnlu+hLg4lWjaa0Xl2HYI1tfuPNpdK5XhiQF9KiS
vWuMfOQDetflA8RgZ+YsPOmRmHHPoNPPFu7Bpe6Ohnf+37wV/LL8x4vyyLjdX/4o
qowKeHD7oefrtohVaxaMkvvsdetSOvYuZstPOGAtTdAL6kMmepxF/b3dTyfXBuPG
nkpPt8CyAqjhbFAxx70r9FMkGfzY3aeGpI8qciFRzmrl8QMI+U527dESzFYO5mZP
LRo6WXJMqS8fCjdFgbSx6ylLCBIBEA8pHEyxTmT7rPq0DrIwgXbmjkuT7PJyd4oc
0J3SDdVj4IuiZcuHaSyjegzhguXuqIbCoaJvjmkrd5UFhLM8GApHy+7wuidTrXeD
Shob5fquUzFWbz5XymTORp8ajvrtogiB3MwY3B0xkQx/lRqne7d6eEJOcrOMYL27
bfi89G9ozWpxnTpenr2It4rzsojjehFwwNdR1TGQB5ii67LB9rSpzohhIwv12zwm
32ilXUz833M3U6RyMVvJAleWKdtBXoJXhmv7V2E3a1prsHE5CckazLTvcLeFG4tt
rC+jYRw40N170OnZ/2KtEJf5PbgBANueQ43WMgSpl3d+Rrq3waEw/cOEUC86GruA
ArB5MEDzgd02kxeMTkT5w5rvuT3Fu5Au3Q2c6wu83CA2ESla+As00OSJbenT8iwV
rexRlGI6t3aAqy2shGtcfIpIh/d5ooA2ScCcZqzR5ObV2aPsi0Z/0qdlgr+bGc8a
JNDsQ4DxbO3ctLHpPUCl2u+VnQEz9wcgGF1LsM0A+mNF+2HYRp7i3pkZ7bOLOt1K
yR02AvVBUKhwy03XlxBkBMMylXzBzyxeooeFSAUNCYz0uglyPxTSU0aWrYdEKIyl
vhy9z/EmkiUz4qsPpIkuR2srLsnQJxmVvTN6lXgtYysO0eGkYGrSSeAkmAy7Ac41
4+g5e9MMzLWX/DtNMlRUUyA6lRxZoj0btRUKmhnfjVO9JHwznh10YjFksZzcAKQI
wkzsg33sgeT9zacd6QnMDPZrBKHw6q/Z61I25PEoXaXelgSsbHBAFZvaKpB/FO9C
ap8efS9Cb9I3io8b36wDMtJafUYZq5WDYL7knKK8XTaHsC5suTLSSpYU9xHkuy+9
sFcLqFu9i8K+Z6XCABSKhqdsVyKgnl1daQ6Ttr+BeRSE3ZkOmThQuv1+R/V6hSOa
faRflEgbMDkaIAlo6h6aUsEvirVNjQkCOqc39oVs/FSPlrgvT4PW8391kKoxMIrm
slEQNaXYLiNnodQ/L0xKthcO424Kr8XJ+k2rLNP6pktKSuzwDB2drh80fBeaEs9i
YaGwP73/on00VA4VICLMOfY9jhBmvKQhNNK8blAJ11BiWw55thiZQ1Y+bR/X6zbe
DqN3Ju+cxlqXMu4JwtwybmTc6FAZz4Kzurij9JomTCnnBAjZKigkBNr4GFQTUUvS
Rs2kyU5Gx0f+aa2SHHzJEJbeRG4cD/+BGBKfAPONtkCOzRHbx/iuq66OmDFHNr6H
cY6DOv+vSi09ASHxzn37fWaJPwy7NoC40SYSJvAQrsk0JXwOSNJHjzoFuKxl3QkQ
sMkreIa6rsoouPNFEylBQUs1WG3/5Htbns5s0ddtqHPKnt/MSOV6K2XqAIstdZkH
g+vD3T0sB9noV+xFjaTrs1BPVUIrbJVqU34pZZBuHQxu4P4Jz5AezTVqUVsKToXi
LWl7UO/kk1HO78bD3jkWSblQDpfBDyCkOtbLvkz7GP6TcDXAY7mDHGTfae/GI4fR
7KxsH40WD/o9Sd9SQ75+D04897oEngOpKN/gIGB+O3xRTV429tP8EZM8IcQzmekK
b3u5jAecqHQHywb6SZSBmy0Q0Fuh2itynevZNwywq5TSIQ8AG+xQv3/m/9Egm8eH
89mz2H8ct6+26IffsXkTDyqOE5uBCLw+CX7QtbTKrQ/73I787jk0t2gFnteI2l3b
4Guvaw48+ho3SJ8e7I/40OsCF+p1z17/FE/yAhobVvFYq9joFwGBAclKsYzv9PTi
UfizVSu2DvAWHJwFTvtDGcU9BV2y/2S4k3mD3FsSsYndrN+A8JtTUH5a9irP06/D
17ZJqpOyQ15k2Y6gWqBcSw4MfEuVLyxSPMIY+8lo2k57h/U6LRpz1KFVuu0wKs/X
+1B0KwDlooH1vfPa0ec/kNXDwO7xbWyQGxN3JBITAYQo39fnTyrJTiKIGHEF1siY
oaxI52IWIY3YanPMlcpvDzKh5gIMB5ICyG1uHoruReY0uVWQKRSHjIaJ0pczGw4F
H7ERYYzYVYP+bin1ep6uj1+JEXNew7RnLFCb+I6Ul29KeZqsu8K/cBZ5Zbx1ehH7
4s5JwQAG4t+GBqbkigz7kvx/p7ggIq8ZQ4JyK6BITDOgRtX6q8358i0azmbagVvx
ZugS8X70M1rT2CFmkkt52LeHDkCxRz8PF9BxFzBQrP8GFen8amEaSOI9/fWag5+Z
Vk+orsluR4CmaBvLq0FwS3O6PSW0wFAQubonAs4q47FpYzqUlRw7nY2xc69lU+qP
yYCUSlDCVWVydcDzfHxZQZGgXaY1qTPH345W9jb7uUBTeCr1h3YA/1BSw7n6fvvH
1b2L9v9tGELr5/LzoPJTro3kpRSHEoLla7QwruT7JumIsxa0KQXUqzdgmZr3WeQ0
YCGSl8r+h/YqUfN8ZsAXOsCDQAkFcIuoYKy2HaANbho2Cp5uUlmDcyRczPXe0JOr
p9TVJ7yUHnF/yzi92IGgwMT01WvADsqkhji870TYH42YxhaeEtCn7cAu+Vy5O3g/
7jp4jBgE8TLREzoE1gkCQ8Zq6T/vD3XBIwCSZ4ZTqEXi0LDTICphSqnpXHjcreuQ
ir5cqU4eiYdes/OhdwECA+wHYvGkl4/ptGZlVJsBhu5MEewPOx00E1RU/OOzUnVU
a6y60lwk3T8SDQ3mc7cecK/d4sqWmEgbe+pyRq4AklJLE0zt1SQ0BV7exCfb2Gy9
FVmwRt89D7/kuG+51wgp6wp9TQrxFJAl85CdOStIJ7aHoC27UswpBBJtUwhtSzQS
R6p1WC0S98L1sEwLhl/M8K9qPE+CbiXJFthDVrkjXvbkokMAeBsKIuD90eW29Eeg
sbbWoMwct2f5xqgCbu4JfczayY+lL4k9vHB3z3uFOJPuEmfLUPd8ux/FyrTHs1Ef
t2LLobgu/eJkWhVZhBHQtaLbqxfQKM1A33jY8qY63cl8sm0wPicVw8UgS3vivNhD
NQQjktAeHHjmuUe+1Kjt7HmiKjwm+y96LGd0j7Q4Li+74D3E3bV5/hhu+0IiiLM+
NdVKNmRhGBMl0FfIuVsSBn0NKDt0vVAhkII3wdvRAHT/1aFFZGKKYN+fsWRP/5Ml
PFMru32+A1iGi3qXyop51T6Z7//lv3HJCN0gYK8yhPrehOTKtNFMBj6hVCDV5bB2
w7811kBRgxSfdT5MQtf1aAg2lFWs7rmSflrWB33s81TYaHB2rAE42UDEp1mPLa3T
tP6rUva5H7tM8wPpo5Iy7B6/yNw4AmO4RMwDjNLArlj03kBzaAZcTTA9wfs/jsCs
gizsbPl5JIkLj92liNSJriLOP/kPFJfHgA4EqIPUBQeFBOZqtBhQfsdFsl1U+hna
9vy2cUf2xMW2coXyb0BJqRUkG6WXg6QSD6cgHthyIx33q75/7nfom1dUacpRPQT7
h3Jh06RhVPlNvFdeqVetLR1oiRXAKWXV6SAF2QbTzjxHz7vzJqOTNPMkZjAR7I2B
wi3HRZdadMYQeg7Mh5yEmmUMIZeCpMRur8ogeYVNm6q557njlczb2dKY302q29nW
/XTPDhEx5w/hZ15usv6a338APRILKybJTviPk85ohL4sAKT1v2Y4NsSFPV7As20t
CKy4mnZT28czxAJzfsF1U73kGfFQK6xe2Xffj2FHsLbpBkkRKfbnqhmsfel2LiG5
YXcfFRcOJUr+A/AzhcpAmeTMitUbzz8CD0T+bkuNoDszpnEjLRuPpG3RUB/i5007
/1woceX8FmHvD0KnGdHUEKF+Z5miX+jzvphjPYdv9LHl7LFKdVH0bovPpU54P/e3
0OWK60TbUYHIzIxqWzAwQacDvnKs8SOn114H/I9yMrHShikAbnPcAZRVu4zhcKT9
CkdZkDkZKnc992aj/Sy5dv7s/IPn3cEH6O3z4PBrB1h6DrmwE8x6HLoCQE4tKEQX
bOQgGZ6zZlorr+ilQ/Wl5nMlcvBmWnmn73Od/2v+aKeWrJ0HasLs2/ZAPajdLgQv
iLRGKiNnZHh5UMRc9pb6K2fKG9MNvF483kd4qpnm4Tvjza9M8O1F/VrwxgW3FBEU
m2C9WDDNjv1kITH7TiBBPY6mUx112u7gxsmojkFYLT0zao0ovwo0y8p3lRLc5GrL
HmPYkk5BD5JSUAVH57XWqwPWpL1hycI4H6MePz2ia7kmHf6pi9piOr5z7Avv/SIG
GrbwIMagcQb2rsPk/OsLXkrSxUovjyegLHtC7e3+tXTPbhg5MtD0OXbM/NtSxsb8
3XmngBxPIvYnJSx2SOyNB6OQsgohN2IDPi7z0X2/aCc0G2ey1OwbVYbUzflWYZKk
lhmlWY+QPIZ+xqQ+KPpl16aKcrBs8PaL8YQFscb0NAGPyovQg0h97M4ZDH9K+Tnn
j0LLdqWx1Rzt+9pOLV0w+1tM+mVeNT8r4BLPa4EOGKHQNQmZ05H3R5gFYzMeGZ0J
vmfTsiF+i363vPwnOPDZ7IhDxo6817D2WaXYdBYxzKyvnWWhnVFqGRUCU3tQ+D/q
T09UGKMt4SQ2yPfjEbnjqIAxtOQcTD9OUkU6x2PiGLV99it50C/cmjODRdtIMxE8
HaKm+2KLStzCxqk8R2mz4d8XWF2eWefvNC91tsDrxN4YaxwYD+PV321YQ5yvBlRN
sVwwBUVu+O3c0rPzESYedYd+ohxEQSqiagpkyxordrFyWKVOM3gZqQD8xgL0KFRW
F1pNPEHRZwmnYWTdeFVdi31YAL8RF1BGmTO3OH+o3JnsZa3P0NaeGhG9WFPHHSVU
Hr50JdycEgVgjneoBpJ9wwbcUmp6c6MaLLGXJrfDCuUuEJGglq2AMykDTCeRMeGM
Qw0obGlSNcZO3CgHBwo70hQpO1psGbLXz2QeWLSUjTSjJ73aB5Rg5XsLIjzUqNLw
X+6g+cjGk4wK3SQKQTIw7UA4vdTK9j+RRYBf33CZsv2LuUZ77gchIRiTiEYb96M4
TLnNbtTnLkysqaK/o+4X5thROnYhegyA+pAl8U1NfVy6ehHK5mk/RiHe/EEzlbb8
vZJqSlXdebKYUC3uhZKCfAMxspuryCrDfFCCLQhaV9uiojc2h+ZD0iHHa0lwDRUs
somCiERw5jeIzoz4Z4GDj4T/Hb2ljyX0uNSE5Ms7JCGWcEoaVwgXVWqkLlaMrAfd
1k+1W4QJRakv4frjxdYkpqUGqmjpz9Ezfq13YJzfPfQhRf2MsrCbyfKTam4uVYu1
3U3baU+Nwx0iPI8j2qKY3CNbCaoAxAF/Q1i9w3yGxYUT+UNYGMnhv8BjQx1iy8rC
35GR7Q5aY33m7QwFgpvb54hDbBiU0z1i8E3goTzIanqdaxBm7MrDjoFn5x4PgrSH
qHpQ54QaNJULjkElwuuCpibhqNSBlypBV76Q8EYhk7uu9rfncSSCXiefwMRksfXa
jD4Mjlj5sBrxUx6YNGpJTj3FsPliQ/BVhV4Aj1O38ARwTb2w57WiVP9e83wMc3Qa
BnqS6PxKNdpjooVEmwaVjZ3DwcvJyC1WnioHUpcnve3vfUlFmTrKnmRDp1A8xmXo
rQIhEXsGvU6Qc/gGacTFFMdyo+U70Z/k7gimwoqHmXrdmSkZiH9a+3F1H9poS42J
aow26JVGhOFfLQezRg0JgBtsfREJ4j2BTHHSQrk6OTqbF/5F0XhRH2LV4YIL7pXd
jjqm2fArMMQJ1GWxONhf/9K6TrmaF+MK4dHkQP/u+TJq5MCbmXSOH79Eq3fqN7aa
OZ0X0e3CWbihSnnKMshuiZxDXfd6fW2bQ13fux+1vUzGwwtaIw1/YMXux5h30Yzl
0RZMJzTYiUEmuNR8y4/hi5wwi2PdYfK/A3Tg6WURUMuK+KwAhSLcvLJ0lo4H0SyB
8GwR2D2u64j5Di2asQDpEbMpctRBteWvrCr3GyPIXI9B8qrKm9aGDmAuRlIH/Lou
SUbNeuyj7e1oqC7P2PZA8eSsVouq/n9oV6mnxsQGd11TA8hWezz8ogkTWGsGBT7k
06TecFAhAEjwD+hkJLL29BxQxYbWkM8W43HZT3TCvB8Pxc141XRf7EtiGmd6yiP1
OhpML89K6U4NRKl4z+pb8B+bIli99WLPs6iS6MvroVCiXTP8vlzRvesbr78CDvBE
LGr3FvKfhDCc7TdPZlhXpE5iUyLfl/HHHQLuPuSeCBamn1PSLTC8B3B4ZpJMSB3c
0UlvAItBkOZAIzXIHE2cTs4e0e9iB/NU+jWO9nMeX2RPLGkZZfEYCwmMdLuJgWRL
4Htcy8DnxKDm+4WQo8wjLodfWuqhBXQEEMCY+rchQ03K1RK7v18DX3MN8qFmzq0F
jgz4gdjzH6ESwZFkbiZsIXBGth0erT13ZigUd7YrTtVerEPbYdFSshERTzA0fctB
KpLw1Uy+Ck1Z/dkOF0S7EMntTL9yEQg1rIMU81blgvNlas6/y+FUbtaCVIiZMGAV
rsQfd3SFR+OwBvbJYgb6BGi06A/vCssxWfhcb2w2TxMd7SoFB62cvwPSutvAClPl
UtRg15kgxr/okZMOuKcf6SISFIVLOv85vs748W8nkBCni8+15ewDADIKepgEAhtp
d+SGwfWMwdxstsW8NgyCT+/J2Hnd4AfhXSkLwVoj6jAo5gR2hf2mEGDN5DWpAq6n
XVfUuNDDdabD8tIWfoWoKj709jJplyBuf+puPLteGr+9jkZdaS63NVkZZXPJUgUd
8CgfcrbOKHax8RH+ZBTPRiUkVQcNOopgR8RWOR4VWFG50C8rl8IoZ5sHPSkIel/9
RgELA6FRW3MoSk9PQbcu/0RS71qFhZ7wUq5wxpu7c/nuXP0ZryOOiCYeNYuChl9Q
nvTH5TuzUulzNsnU2GEx9+219D7MRnuuRcnzQMDgDBMIgDbRtu3SyvTqiRk/lFyY
W9iS7FFAruJLZSOK/Eonv26GsLtlGB8oxv5p9jT5sF6qCcQqYmGnAeyhx3p4OOyT
oYyXUJu8o9uW/QEci1L6F3sm1HpPgZ9YMAS9LbGJc3dhKBJnLJvM2kcfbv1rTfd+
EL1rSo6/Hdv2UC5BCtiMK5l6bKg/va44GTLjJ2gxFZ1dxCr3wSBfIwpyrWHH4acn
mbZzqZCe/J78oV1FtfOJf4wBMYnMI6Fjj4hozBDAnont4EQYdJOqJP5fkeL1ix6R
TqyMOeMkuI0U2XkeIh0PtB/B0IZgBBT5xswjILU6ZrP+FSZp6jl69zjsPuvLSiSA
3TzkiV7WXMfDsRmCepseEigOhOrUxYWKRPp8RWyy3rnzW2ovzWMMOyeFemvpC9Mi
R37MKPppvOxgybL8OzVCy5Zortza1+cBNKEViOCH1KS7YNwiZ4XXSGZgXT4rp52p
y3nvK9DmMVTr6LMm1Zhu7QLxuO0TWmF3fD7/+ScO7Ugx0LdaWU5sjQ4sPtH6bmRU
aSVFVoVn+6JpeA0J2d+8Tkk01cJjcGkkr4MP1DwWkbJB2Tln+fCjvvFdQBySLBBN
0w9ur4XXRTL3bOMzwdDd9HX6bw1OnTYHGALifDi5eYTMMUYoVqRLb3XFum5fnQDk
DVAcNVzxUoGSYUL1PxbJD5EQp1BFo81nH+a0xpDfTiknamKrLoFgl0s89JQS8ANM
WG1Wr99YaTU5/ENHmaZg2wzfY2B1AClvOP7aQis2ZQ8PT7lnasm0pFmodh7MlIGg
7PgPYZt/TLPotPoxx8ZnPi2gqQNuC9+QeIAVQC/nPUilMtf2zkbw2LYKXce7QGgX
50iWA8dLfwGC521j3iahMKsHodK18ZYD5WX2sX4kMOCt35gqEovrjTfgT82GC1nL
6a2mJJuNjG+d5Bh4ogvCdKtYaPwxT3nZ17Qih1JbC2n7thZ/pLkJob+jYxeg7tsm
vefs1Ij3Qz5gh5RMk2aSLr8O0XpYFygi9/zqJtF/gmjg0RLul78moRpZml+h+Vip
k/RZQuGGVmjjBC47T9smkxG1EowkAGzXUDOxfQVa/17u5qIqjFilZYAceR6KPwCT
h0bCiBl82o/No8NceYJW3u2wEn1AIzNPNnQQw4NTLb7RQYjBw+eMnSewfAawqi1/
bosdd+vwdgF7j48cLpiY5LN0hQr3cHbScZ42W7L2yZcwkiPxwNjr95bhqJFv4p9b
tC50dW2Y5fg1N7TEzS/mMgwGHizAkuRihymwm8t+5KRwswVlCuhOZK3H/6RI9kJy
3LhHtPsskRKogSTpTEHEhol7iq4fstb/8dm+ukGeWHAajO/dteYxjc+gJ0H/lMp3
ltq7GJJ8AWDQc962SD3Dvu9sigtpUc9XoIotun4gk2cmwPzMQJzzGu/wYjGJpKe5
z6VAGxsNOvj+lCGTdtpRptWpsP6Cuv4ccYpT3p8K/oNyncOzp3+SO/YaZ+kcDmIM
sLtSs+TCA0Yn19TazKsVo5MPyqUaboVJ0aN7cD0kITHIOhIFlaNqHEKjqAvUXmMs
xeGIleoSupzTWdjVbxXP4x0h4uC6w10K+3VNB4vsIu++2ODwrB8nWsHLdI9XLS5W
bJNP7wCtsf82/APKXgSFuntoAPAjH1KDFtIDsksQWmpv7tPYeTolVrdo43CvPnIJ
g77AwtLdPLoFucudca+Jt1XisZajI0wnWjjeHtM3+Pc3GEl/2CD6N7dhdvD52a4K
OwxvCe24nYE0yEYIbFTsMi7dA7RFKrSLY7fWChGT/vrizdP4xMtRWDWN228BXIQw
30lt/QUvfDwWloU6oGA0tjdIhuqma3RGD5XxN4flKfxgMdxA50V5cGdRtK2o/vL1
bAI4zprxNCGGDVe6vr9sWSlt95yNkxvKaIDKpn8u2LbgX2Q7BY9MZS54C3PdNH26
J5P4mGfuvopHmMJezJoCpjOz5Oz1gK37drCN347XH0Bbro4W9pPi70bp5WcMFFFc
rf3IeSuy39Npw3MWSLEzV/zgMQXKx0DLha4Gvt09PUMdJsK+NgfnoMX8mU+mGBP0
5pc5nLpov29ma+qFWrTptnf0VO7VJ7Hdmgr5NuWj1TgsJfleL2HtF+Sk1qbArVAl
W/sxb9wGL4d8VwgyC91FVa3lj3Yt8gAuwPPSIDCgsveL3QB5cm65OPJUumuRwlFp
YgF9LA9PE3+VYKk3K6evkDnPKLPQ6SrFKBsnvRRVW5xanP6EGfmE9vIWd7rySkKU
7rtXG3hcAJH1ui7Hy0dtAlsQI7u6ovjZpfzpx71c3xuIRwXDTtd0t/NXAM9AhUdA
/vSkcScLLX5EfcXxMV9or8/xJsh6HXSaJHpXaN1R30Q5vANFndavpqODCCSMXXQ8
1OJzX2hRakePR9KvsIudVgz/FUqUcydDJYgUtcmDI+fj6MH9mbW1zBwd1O1d2H8l
wvUvLU1v42mxvfH9kRSZPjuZDkvGR/LkHNmBVOKgiq08qhFZPVfz4HyXNujmp5XI
lf2Wkan58TKYVW8AbuhAuL46dgxbnm5D5l9308woivCLtzEAEWMO+lJtW1TknwpD
zs0FS7gGQxGcTVnJ/jgs47Bci4aLj+yRqv8q9Xwn/cGqDec6o6MhJtj3r8dtA7Ap
9k1aYY/sPwOz9IrinAmi4dTciNKzFMLy0mLnpUmLXpIlkx34zauu/IVdW2zHOmkH
skuqA1dkLMjW61cMRH8E+xEad1AZ+uR+nC18yPdzNPgiQE2pfzqCfZ3PiK6I8YIx
wwhSn7SGGtGsBVaMz8RoxdX+gbH5MpryNggPtEmP04GIbZ729mlXFpW2ONMmLXhk
JQm19RW90LaIF4qEM10VR9rUn6fKAoLwDklCzKMTBqzsQ8FZumHS41paLLu7KUYf
gj3e2w+bufso/bwzPJeyRnUWy90bx7200oxd4hU6OdzoQSqZjGrgoD2zff9AN9Z2
x6AjnXH0ALr13VHUoqWz83jZYB58AAlc3ml5mck9kI1laRDJlJXrcB6aTPtLXTVa
Yh+qPR0hlj01xuKAU8hGkz/mJdMzEd0QBVw1tscHNci1xZkz4nvFz5zjPlnh/Tvv
OQUgLBbAvgES9m14/pP7cqzuOlp561C98wqsd1KoIUyQ51QF/Nnz7VDLO163rGq7
TV/qjjP8emqxaLqUak7M6lNoZdf4mRArpI1H/HDkuaOEZmOy6YZHg2Ts4SWdEA1n
qpZAwlurDTDr7n7dv/INK0clOA2aSi8VusSJmSCfl4HownvB8ev/6uF0fMr8hxcV
GiUEXGkONCGhqwGYKe+R6eJgLgCpEKqJ+zuHMr1CQDxevL5JgiAicDsiYFsUjB5T
jyYHcUhALeArTUrpMOjKg3Tfsw3EKW29VbxwqFAN5HFC4gxx8rRAf5Ge+6zEgXMF
Zwn02yuxn8KR4iQF3c+QSToxl7WHMeLLYMCeRSmEqkdE7MlA9iYZPSMRIUA+J3rj
nsGHKegiLk4TNCzHw0gkmShfFKajoINTX4LhfjXrQFj3TzFCvfIJzQ4TsaoNKczK
SxGtNPGNmT3fEiPv+Oq5zlWAUaTA+tO49ZBphMEGmpa0qwdeurIteG1yXnb0Pe8h
t8sr67KpHo8M5Sa6ShplNE2VL7ANVSsM3IGFLmbB6ZWs7OzuJyOa73R0RVz+xEh1
ojy283iQ7nXdgLee9r4HkwrlTqU5tAK8GMDe5srqw0m3ehAKoUVQMsxhqK6nozpF
Io8GzZYHMovJzs7ZOpvbzUjASX+XCQUtERReaUxgk391L6i+dGM+zZ4b0yN/eTlD
kkjrAZEsO/6jO1pT3QuA9a8nCkqXnhlzQizySCPB16L7Q0SQyFTo4n4ZcfEjPtEG
NymW/819TPo7raYCnEeYBOWMAmM+MkLzelhscs8l5O9+H8sLl76eN8KxejwcqhtT
Wc1AauEUv/+u4EWHU/ppKNiWegh7fr31xt97k5BSAleTWiMwiuLa+BocgsNSFSrf
gBUk+rHf4HXdqSpvgU1f+faY45Qa2WmWuiR4/tUhspSP+6vkAC/HqIbw4ZhPsJkF
Cje/s958O7IqFAwjSPOUMSKBX3VAaUz5FstHi0tFGRQC7Tui0DpZMZ8yMpeW5LYZ
YzrOg9cSrv0Lehsdt6HPZWreB5yzNP5apzuLAqb6S6y0xx1M3OJ9kXvYu/aT9ui9
K5DeytXnWO8U2nWK5obnSkbYm4fr/kdV0iVdbC8p4EjVfKtR/YgDFvuAh0XQhShy
W6wFgRvJjl+I8jltvccw+4iFGIHtEuVtUNmNa4f/UKVlgAT6x7JcbVhOWzZnxRF/
SEOf7stnJj6vxhuDAL9XiZQv2O9s9prBW2D6KrVgmlGzylQ78NKsA7woUUBPxHx6
Xm4WbWua1JWHIG8m8q2ZiEHrdQskqoCiGq9lL+7Fa5E5/7bu79bNZYyXfx+Ircpj
iS3wPqNkIkgnsFhp3XtG4ZhWZnpRR85wE9pnBWyYuVNup3ABcrsZaUtYFnYLtqhw
GuTqAbkZLqx6k22yJgIAzDuDkuCe6lwVCfS22YB8A/o6CbUvxJAgoyEAnmePBvJU
UfviBFKTW7oSP/Vv+UD/nA/eycDYZWPddt2vAyxHykIEfKwI/hgpKQoHHm3DcKva
OpL+b+RjiM0EwdZ69lUySqazcaXKfqjf6VDAZxxH8dNDNlkYuvu7MxWhY3tBniKE
H4Lu5BUOrg2hyIQZfKOvPmXpUe0OgOf8NuqF3rwqrKZ9dCmaNASdzkSp4SbVYCK0
bxWUNL2DctuE+ZyyRmGYM9zbvWUFTk2Rxv+xYvuBOM9Fa64xkvGdLatOv2jxmiU4
SSRtxTKxavP9JKDVZ6S2IiIgtPsnpeARj/+iv5VOjOXBkGUvpGtapOHq87TzeIyF
r5vbklCK3nmpYb6BLaQgGiC1EVMBckY/QRkSPJJdoF1FLl4zJ9pNEpeUIGT4/WHg
YbwAG0sUgu+zZ8WvQglSTKumsyl/nU1i9uKxkV7TBLkhaEIYh0hoP/vzdjRMTXkn
uulxCoBX4Bx1PHcbgvH5+gFLRuP1/xho2D2xmRIXaPg4UAYDg+Twhj6mavC8+15e
9AnybOtWeoTsojaAUWh5ixhtuz5H9LzNErQMdoQa0dPRnJ7K1hQ81Ft8ilTGObWD
VGvkgMnvZ6sH+Z91pGMMNfGqQX2NTKyGn89rdyd42G9+nnrLjKNOHw1+JWHo4js7
0vnOeXV1dOhvo55rJZ9jyngzzVjEvdEzdMqkdfxTh7yPw4kkkXLU5scP18u1Kcx3
EE9VK5OHUa8Y0oEHHrF4+I5G8wiuoSd3OLosgcmHiZ8yJ3Do6qam+XVTq8x+Bh1g
LLeABa+meJIQ4pATfW25Qp4HMErrhKhdoOgu8HVfYU7rsFCSOLwhEyvxXMl4fpfZ
QbwwAeS7FHI3zYOv0ocydmAneAuhweX27Rym4rdV8n6TMp+6cexKfR8vl1apGkXP
9ssX9ykiqoOQNPu3lRqPdhB1dL4uKol/qyN1t1gnEHzKl7rfS9I/8+fhRZDGOBsR
+Q+dCKFRkLwUIazw2HO8NIM1KimoPRo2NbDANgktITdeEsWC3rjClmf/anv+RQvS
rKudaDxOMBG5NO7jem9fLipa62/k4jnOZ9RieoNwp1PDOa4MdWRqNhmDJLhf6kVP
VVjQEHMJmmLOee+KD4V7e+3CjAqapkuYY5/WMSJpkIDoBqrGTvEz3b5Dm2nUvYhR
sJPCFJI3jCRZx7sx0Bs/q1okIWN1TLEh5JWbgG7XgSJahOW+oR5L8vDTbjIV9gri
rvOkbrY8uDl9wZTSOa3+n9tqUPLZp8ZZ/Kh9uRhqOfJTvcOGEiRGuXmUh7+nCaZC
Ie91dqPS8MzJGi5zMwoXDCLC2s/EHzEEMoWt5z1hImNiLg1LxClSrYJPyjI9DJvO
nDY4/NNZIi+KoiOtgXruC94d5yuE72NmPVNBLJ+6luV+G3uNIU1atDbEtIQfgUmP
P/fxF48tYBF6BV1j1KhwLrwFXSyZZoBRFy3yubO02aCNfgEbyQaVVY6P+m3cxkdi
yyyOoTdy0Z2mzFPm9tmvNHGnXgoxY5MA/RGanlrPGpeyY25UsXaEuvQFSZl5htXw
7EaahvfyzTsoIombre1vdit4KwdJavvzfuIc4iDBGcgOH/Qvgm2u5f2XTGYETcMy
AZ21ILEziHPFQFhoz2Tw/OcGo76ElP4eI9Bctw/5hKip85mpU3FSzdB8Y6szoWfU
YVY+ifsnT68wgjS5Yx9AAKHGFFR5arJKkM2Zea+35ofwg3D3ZMJ2jd/dxF/H8d8D
vcEqKOwjTpgWVQ+8EgJt/iAONlNCW9hwYC37UKzvzn6D96pXVpqhU4O+j1mf15KV
A/r+yJewr2543l7jE0hRgE2eG3RvclKnlFaMpgLMYy9Cx0iHEc7sA8OuOCU+ONdJ
ip0Ve8GEkZNSqoJCuC5AW6K99XbhVYPch4GPPVF5zTcistUrPvWoRWNwMgnlbbdg
yyG+Mbsms81Dtx32vUYM9tni6yQ3gPxXTOqiIETKlOQgMghfJQYwW1Y8eO0nq2w5
WCGE6lGaU6GMAz10FvTOqtvFMn/FssSNzc7PnM8grZi4472cYXdd6F0wyo0+SzL/
HD8YtNkjx6vD3B9J/hpnl5kuRWLF8T/VgILQD4oOnY5Fa9nFG7WBctQfqd+xQrLe
6hEEC8/Q/y0PGJ/qK9aDV+fb7qrywcwqGFfRpvwliqw7Tuw+nMgSQvOWflfag5I5
LBs2WyOlfslz9NIW3U1RG6KJ87aPKpxX9qXu+hc2XPYqjkhXpWigO4JxbNABFzXq
IAlMhqOhR3AVwWWTle/4n3Oj+eLCuBD3gdYxI0pVkJKbaBwPJFiC+aO3li2YfkfT
NsK7w02RaRujpGwC1j1O7ibkzrxJs7dq0rPEYhhglMzKPnGuh/Hg74ozaniCbRP9
JO8EiPlTkv26gHl0FopfWtDJeoBTvUCKbnIqPJbzUTokyMwmrkHJr38lad+LgfQI
g5Tf4q6qCiHV2wnwIxWTffz0lDWeaOpFcW+R9YPue7R7dRyEbbHhao0aGjN9/EE/
bVrZaWD/DnPn+sVgyQat8XAA/Qwwzu0FMxZO628LVG/mG3cz/G1b3kBh4pp/6gEX
O6S8zAvAAHm4iebrZDEG2/p6ILCUPf3/tpPT/50q8C/9k0H6EKPTguOORn7SXeWm
am11lVrO/Ki19zFgyeHmRrQn3tKxKXN4qVBDc86VL8QTX9RI8tkGZFfwWZAo1et1
Lva6hCgLbkLJ2xNG3k/gqn1HEI2ZWDRDv7CoMwU5REFtK6a97FdyaJ8UqwyZzKcb
hL+UZ0y3t1JC+/E82L417mgejfYqglLjGIq4qMYStb4SwZ4GPXGzsZ0eXNDFqDQx
wjUzHOa5kjRCKCKeXglwsI3UaEinDB87YnE5vMfQmDmlq9IOBt3qwxs3ovsq0ZcM
bB7v4bU1WJ5Xv5UZ/XYvJZgQVNIGmye0hUI9U9JKWFFPeF24zjjhI7J5DmtR65Wn
zq+aBJQJ8U9+dRThzJXdpBZswCtXbTbtTJDRZVTZLvaWL7mNBijUrx7aDuTvD1/R
9wezVUaFFeoZH6B/dd81ypWeVP/d+Aw7VFnNawgH1caJ6uQQUOTnNTvP9zBcTcx6
CAAZfwVd60tqPwkxmIpiG7hDkk2JRm77wvJPUgrl0P7ViT8NUkB0qYbpt5VfF6F4
QbhUif7D93JJRu7jMUHbG9CtYwzV+pP+ziRVbChN9cFhSjWdvQX2YLoLA0J1QvuK
PfsFR/FpC2WP8esGgMvSaI/JKAhU2/RVLpnwhb1iGTC0zO6ATRCtw4H83rHqBcD9
cGlz+Ohl1Qgp0iA5/CrV3IT9FTmoim+wnwVOARrLI4PIF8TKwNOFGwkfKJomlnoS
E9x3YwPA22bh+8RL+t7ff7eRAWRtJip6SIE1NACrCQklZUireq9xWX1DarawWQ3B
d7CBA+qVm6raCLJpLqo0UgnlPr7NlpIcZPZuLZdTvbtUh5Z8Nv2QMmT6Jz0aqwJo
KkPYxIKVHEhdEiVZ+xDCSNe0hfQG55N5dnxxH4ofNPwry3SkQgjimfdcqMEKJJ+B
7sLvwlVWbttbCUpPGeky77F7j1/scgjj8gjslgdjuCtRT0wT1qFQtCQlpimfaGXA
hea1KPlBkHU0eZ2xGqGwC9K9gB3RmelzKTL+3+44KEAJZcQ002IgZst/P8H+zyrJ
ned0T6+meYUm5LnDO3rTb7yOG5eBo+tNiyXPtMFwMY86EU5Zb2o9R58PKHzdj3rp
wyY65kFMREX4l/QU6VLHXiUlc3JafkdVsOG61xYPaQtHNdu5+NdCWHdWQB4Z7/TE
ZmXQ10YFb4/OltNtsfpEg14ZjPTAOtkPxAnrZKsDcwLc8cdCuuj/pXiPoFDiqAF3
ujKneduQ/VVMNNhnIO48dOXdyUwxqTNYBfH3u80XMn/+3cRnrTOvXUu0YpybXiSf
+UUeWkzl0XXBAYVFWrUOW1O8DTDZpX4N49XImGOeZXihtPKUALyP3zACsnqH81e6
41BqydCaEdSHOEso2T0CYhmeUxp3/W1jtByDCyWy+fIZxObHEyeihmQ0JrJcOCj4
+wF9B6NQp6iE42fyJ7mOuA4dnGYU86H8He7x6OUjL9o7TF1VNVVyMfmv5wtqt/GL
T551+9d33D7Tj/a8unZoZ5DD7bIyEtrjoTGmDjr7DRhXlW5AQmqjy4/F/BNxDphk
0ZzFM/xTTfbHODphVjuSRnj86x2ieCfT2M+GSvtYtUE1IJJW/X3HcMNDJH9VdFtq
hlz5vXa7kR35BxWgjJXDA+3IpmVtuW7wq0kDpF0+SgNvlfHgnCp6PzgMvcMNrdZw
N9TVJyXfYjbdDS65XfHKjUynKU7zGCuTKPmL6pxb0W9VFaSiNsep5uwAFfZuLHCD
LvjSCMBLVU7xyX22TyoWjCgD9bwfHxFrVlVWf8HE7/2NJ+dSxD57Ht++TjjgLaE0
hV5+6jy6d3edD1kbgR9Hh5EUx3Pr4Oh3QZh1aggbAUPnKIfS2CP2h3/LGA7cd/UH
wQi+Y/xfAaERv/SQ/zsZZYPtFYGNABRK44TkSJni+mtb8+6GnkrJOeNnWKT5BYbR
bbXmFSkutCfXRKIOIcio56gOxWhSEKZtrKw1t8xz+I+nIYbUNB6YHuim/A0OmE57
3tS98sMsjn3QHZqG/1R1moUG+epLo8jfsmsxeipX+KnTpM1lgsTqbHYSsNfLTVbz
0erxri2bvjfk50IS3BsxmHKwPppNsEQMFt/cfgiLiPjh5LZg52k2d2mUVPlC16uB
IdEqlMsU+CS7ffPADnXWnvyCwts6mAc6WwldIm1T2uFlvK3jH6dBXr1VgNNNKt+9
m4rDUpfoTm0ZIRnrmBQg2uxnttXJ2Ok9YTRUeB8J00GFJPDvLSWISInqY9Hrwdtr
cehabFMcS4oE9uk2ZLZII/BxJVaMktNsZdAoUkCR7/cwEKB69YbLOSRbEXz1rK7A
yVvj1mny9+lLntH9/Lfnqft5SHiiDi7FEfKGwgCLyMXWt61SFlOXRf8Dln7pIA2V
Vlc4IbwkLm06Ki2KFi1+hiP56BjlrkTyLYxfPT5Zx4mVkyYF2mcIqVBZNNQ0QgOS
xXtFZtc4PqYEZeR5by47cJ+1TxHByDCojBjCUYAnSs4MPEeF+9ROGpedGsT23BhU
RsFGQTqUmkBEgNxznl8qIR/9D0BfjCpbIRSRUIDEvfUnBbJIZpdNDOhl71VIbBx0
SG/cCET62N9DqkY0y8cVNmW/QbwkjxMSNoAIP3b8Uf9Tc1uzT9RBYfXxVgOfe60w
i+v8ArJEa52FRnVfWRoALwzXPNqtNkAyaBNjoddf7hHzE02F2Is4juyKvj6+ZkEI
cc/F9KQPQnGHjLi96pIVk98xKIRW+khHzmo2NPcb3bAY4ttZAn86piG9/bmspjYO
zKUEAzAeqlWc7Gs82Ay6ylDCXDqO0uRQ3acq2wwwqfGiHJLHRLbBNXXnWq29qG0k
QFp27jsPc3ByAAocqKfz7zVi21jx1vJvA0isw9pMwqx4XAdg3BPN69XPul5FBGFs
EWE/c0iPlGvLAnFQwuk+1F11egxmfn+FT2eSzUUwcdsCaqM0kgti/V5gaPekayMR
jBigaYIAWMkTrwVH3yMynQBIPKoLNwEqnMz/bPfV8JJZ217vNVcs7vSMZaGNYIim
LdIlkfkApBaXn6y9De5JvFpW8NyLqaFw3cWCczAxDt+M7RHABoduivtSAyjzhvMx
HRlycYQS+KQTlvpaEthfOriu81CyFxrs4gion5of67MFbP+qTbJRrK8qMbxyDtEP
2QjI0Yolu3Q/nWQ5m6RGj+FfZqIxhJKT9WwmdXrrb8DctOwqdIKTB/AVYC9PtfnO
4OVB/H2YbaIO1UpVJVXtA7TUmrZ854X+jFNZOWMzIHVYofv9M1Wz7MxZWR8Y6d1d
Hd6GxeR7WiweXKByPg6QC3JKZK3emF1B/JoXAQLm+I/EIaPc8G1Tmfq/xYHNxViv
43PQ9hf+TedUFVfuigBt41chqkF/OT+7OigLTwqIXRDK2kE72fvLAZUN3Pv6Z9tw
hbMkI318gY5GuHrFLMdwNjA3KTPuWcZ3Nfwm1aoQKXw8jw3l61+mYQt+9oEnl7Gu
z71SyyGgMIIWsVYKKP6tQ61ywPqfkknbFkxewxG61GoZ2UAZYcBwMB1ZNG9nK+FY
VjJrbvMQgwpPQ3tGoFAqynT/2sqTWFDd5V6nOgw43hrba6XwYKLsQEV8F5zQRi7V
SoYKZ1pOq4sJU6h3mEjUqNTQSTD96Pf7xsOxoIr5YLWx1zRsJ1kV2woQanVP2yUR
rpjZku60LDW8RpuURXKyUd7q5pE3TxJK+iNqTji6hu3o3aZwe8JCCZ1/B2dbzrq9
RX4vnK6GgbVFq9xxOkiiW9TSh0gHTCOkPTr4oxJqpI7plpNrIonvrtezQiCmkb8i
5WAXL2jtNpP9P6txkJzXVWrnN7mS016Uq9iEU5MkSQ8nQ/zmuJFoZWTx0/CrJL/9
aoRuRvMWgYVT6cTatXh4SXimvKzeeI5rtMRjc+p7wu/dYpbrR4R5qcjWycaacNsi
Wf/33WJUNo3flAo7x6eDuGsMVb8vs3c7LeCwLuz+pwFObT+Uz7j2+XcP6yutbnCt
KkWjG9Dql2cl46ttzLpCnCx6uPABKHFVJpW4xxolW1JheV+XrNpwDLK2pvp2jLgV
XZaLL6Xo9PKR9RQytKwtGSugrOOsYJm7R4Ue1x1IBCB8HV904cz8p16MaSL79ODS
A0u0kg2zjwxXL2RlnfryJoy4HcZ0wBhIMMZ6CSNH3RQCyw/i/LbUdbVyGWinsM+q
lEegRxq185HIuEe/tvjHWJmqvmfkCUk7tRaJuthyPR2VLVKR8xyG89RcEhJJy5dx
mWGyaxUpESiYsAbaF3wPfD09g/neIP/6Na7h9F9WzYvmZLJHxKQHkVcdZo7cOWJA
PD4hBLa2rH9cfKBIFlBbm/GvZZMaB1YciHuQxvGtI1jLEqI0I8iXya3ueyWSovLt
avIjZ8DoTZT697jrPXeIOHLreRD1onx10jvGo0YsU9X2iqsB6ETHXCQ3ulHvW7Bq
57Qc+xTNWUgKJ8tsiwIc0Ze9VqkajiTHuM7P2oUcvqkpphQkG65OV0X/kuY+xzlz
N3p/rE6w+ExI94szsN3ShKP2SUosna3JeGTVZs3pKoc5zoWvHsOp46TQ2Ws7WcAj
PeagS1WYhJ8Q6JKm3K3ktf3pCBn47VAI37wTwPHLdQ1VJTP6Nfcm9gQ1t0110kAY
wgdcTBdpGniyMtXG9qK0MJ6j9ofMN4Fe7ZN6N2Z9MYERTWCf8LzEJzivlVuricy1
/TgSChGF4I3jTf5URcnQJTNrcsVecttMYAhNz9JXtp3ffvj3ayVwVAfeQe28T+zs
NLUzn3y3qC6WdNo2InuNesYj0zrjLpyJXmvcjuY7k3VXFt29Vx3OmiUcAgzsU0Y9
RdzU7l0E0ot/4d9zOMDAByp6lflM/zkq3yAo8cPgzoGQyZXErIL12gW4rafL3Mk/
W1GsClbEkP5jDkaBe8bo3Apgl3sW4biSJmkqp2HE/RpR4Q1j+PClotVjk56Tahin
bpCCPEF3rCJVGoHwvzlAxCTyrXDl2MayzmEsL1FxwX2HgOkutvlZIBVbFBU3b6vb
8BL/hxAZbLtqRnHH++vDFaKdmbRhcqloP2TM09vGNu9ktSzK1k4L7JZJPNKtnUHU
6JGBwu6nBowJ5SiJiiATF4kuct1y/Z2n82z++bod0PP0hyFmrrmiBJer0P3Gw5V9
94sLJxqFX+P8M9gC3KScpiMy8qvga0ccqu30raFmwXWmT8vth8gKEtwc9zRrKtf1
p/rdKEXMEUExssFe1FsMy34samkXPDQ9IyvW9Iqs6AsjGRAKopcRgYm++JDDskLW
Z5xXW/Ym+bydTKua92SwhIgFtduiEDqrEelBb1kptrxOfzinc29vjEOhrwCuOUGr
5KKSE+G10T/4JtCoYOK8r8eWZBifuCce640qYL4+UTX2rfLKJO52w19WU8/GsxA9
XfxrqQRliaFKBFcVpvX/2v03BR5kUeOGkKpCBPGEjNX7OlBJTuJpGD/vqusK2Jd0
wJyjnBz2UirFhQ8XJd3UQk7rdSN5SdZ5YGdHJ5If/4VIMrBE22fwINRus6JCPSDM
/2B5NASChDg2ceHMbxDbNrfH6h/1T0fVNJuMf/FMGNhpaBX90dzauaO+9IJbvyKJ
Eq7NhvP7YJ43O5T+cYgBuk/PV7neZHf/H3mf+vxY3jDwIOVczfU5M2ZeeziV/Cg+
n/F/C+glbxIuedwE1bhDC7r1VUJBla2ErvG3DXVKkC/O9HLW/OYXhfDb0W7fOmwG
Qh7MIHbg5TO2Iw7Zk3v/OyRQU+GP98zA1kqOLJd0JOzGN5N9tfoxnObRV9BlSluL
ojrmgsXTMz2Clq0aSUWTIS/xLEPtmiAD+ScCl7Il8ShwRneaewNQiUyctezOMfHh
0OPmcdPvZShRdWZqJtKRbyecZxkKkfrW9YSwaMfMIP9Wu+v82720dAhhA6WRt9hv
FjKjwcN1VA3+CZhs6J7q5VZIJxP4lSSq/4cO2t/8bumXuXy/fds/zgVqNfj7pdbx
L0ALlftNCCQ33RcMVkV+L1YP7ezPiWXCUdeyUo09VJbJ4pJ2hupYDWcRBU98SvyK
b8AHmY4YL7soNCyOQDE1IR1+vZh7ZSyz2iZ4Yfuvfu2bEz0rLJ8dBSU5U/q8d6xI
chOJvAhYHzZZFmq/A3QSXL7q/hPJUSLMOpW2D5DzUu/WKGIyuD9IcQSopRYzDsLT
wjKkpZY5uq9FMw7dFzLtDt7v8kHOFaTPdU4j+r0TzXoTZqqQSI5nt1TLffFp0zjq
RZDoK3EyEBqANDb+LM18DvVKFad+AR8vc+/RXoJhDKbLcqLMCntk9raxY/2+G5z5
PxuhrF5TQPhPl+h6+5+F9TraL9JXc3LUasj50IXGksUwmF16vjk/jNIxHneyCZmw
zBHbrPYre54oGqkH5t3gX3FxcAvx+kq0ETeWSL3OeZ0XGQmN1UUX+B/6ntv8ABb5
utx5nVUblfZpc5GmAXogXrZ84kUxG8/GjH4bxphDkEJTg9w1rynDl7nd/cXxafyE
jOd+PoBiyVVGm9qwIoXRsFHdnepvvHOGwpPWmKzK4c0uBBsvHPCQ91MpNhylu63A
MviUiKU4QOMznMsuXvfVSjC4HB/t8YTSfftc2431v8HWHGPG81Bdc/mUmjHGEMNR
x+hWyFDXXvtsguyt+y0kv+awjiHYdaCbOEMUIYKpKoljBUPcNS7S1LXMOjCRTiis
TRLG0/DD+sYuLDEIcrEmHqIdgX4CROx0aSNsQ++YTFggEJP259ts5Jr9XvLX42yj
PRHl59jJsiAv+DN1jiQV9ztSBKOr9/bR6aJ1wOTgufc4a0kqn4CYs/o5bl9kdsYu
5jox2yXAVT7ebVBMTKGGVQ3VZseOuLgiyPva0HFMEM3X9yuRY8oLWtVGQ8Y83wsm
ZtEipqEg9EMBB5xZwgyUtfpYBlt9zUtQe3OmMLuQYPhiYMTzQgEJmIOzMyLU+joG
meIEOHSaemeJKZbj+W7WgSzEx4L75YV6ojW0xvUiRDH6ss2TFHbBgEDSIETSWOJs
Uyxrh7HseoU819t2pZM0hB5Md8uvgzggxX/vwpAonP1njJ5R3lHkcB+KaCzJaL/d
Od+zuEC4kyX1aCL/1aBw78Y7QVCavrI6ytwlPKP1cmrTb6zmujcrb+ZEV0fulWf9
KpA2nQDNPA2yfFs11W7CW6VSwADC6vlJkIRPCn7YnT4MotqZjlNoViHLlJ7y6EHw
zi0Z77/NaIuc9GPJ1VNfGcP5TL9DwYfn3bTMSW8K+9uEgGWqO7g30soNNFdkSq/G
jxujg217kpehJvhs4j2OsqAR3um718PCO50XQx27tHpGUH874G1bsPo6utlQD6mX
w1/3Cb91v8ictgMb+uJXsadZ+lc1OAZ4sf47r6PORSmleR6E893TjqaTq1RNrI2f
/4wyQt1WMmBmZfBbk0ONiIxkMWqirdzB/uQzTIkAPauCCPiiCB1dYwPCEbo3h656
q/bam16MbldhCK/T7hlz03c40Umc+ASWJWPgW0XGF8UllL0LcEx/tMIhggUSpUHH
tCRX8AKEwWYb/v9vtFhE7SyuMCdbJ6LksnS2eYp6nlAfFURUGvYUuX6Un8GTL31W
EL7ULeSckTcY6bBqammlV1vOmxSHnmvPLNCMpOexolqtbDtqOI3LkSn+guoLTrpO
PrjVObyh/G7oWifJZ3UKdJL6CEbXUgPyjoah6Pg6aWJ6rZoeYzjPLFHoIgDtKntz
oUBVSblZZUOpCJSVipwzjtzEeJ+z3ZxLiEG5jOOpciS8HD2iovQ9+LZrrKCgMaoR
u9bwR1OvexBD1XfzfDItkRxsVhQepRhRe4u9gdEDSLAEEz/l1vdHYrkroXtiF1/V
ddON+6eOt0vSkhi6XeBWpoc1Ew0LO2VxmAWaBmHxsW+Uy3kXb4xxWXbk+gZCNEcD
kOUWn5dqJJ2tLrf7fpU3ezGWk0ypxlZXcEz5M6JbLoSBo+4iU/WRfWDLOdwhg+ud
HOnCKibJrPX0NKhTr7ioxx8s8lt/hV3WYurpFXlvCFm3aN7tOiEKY0sk963tBmLA
foJK/RYWhUCN1mJ7hoZ6DupY8vxpFNQ76UkSGxSaM3kNr1JWamfGKh4Ofr93H50r
TfOqBQyyeBz2Str3tqIjOyKArP6QwXY2wv/CUUKWByj5aSF6oyx6bWFdi4o1yqF1
DJ2A2BAoXD8PnR51VirROSfNyiW8DGC0/Et83VllJkl5VwRkW+BJOsKisn2UdgWI
GsORq8wABd8/uKZcupEl9KiiZnmntV6ZRsKXoDvgTqG4pL/4bY1HMFRFNBZWuHp2
4qpSQcnyJ8UlO8F//fw7mQ3sODRH3J5tjkr4TStWwpQlpkmWJClzqgnS7KMuWRow
n6j6dS8YcCm0us8+9gycJtbiqqJWgt2VbVrEf20Abixn+XP2A9EpBDIszGNQJtG4
2gVLFY4eT7xyz21rCO3rnfDYh//UcLVcZlwOmXo4Ipk4+uGo0w3ruVvRIN5H3euy
5AVZWh9e4NeXtsrDK9w3Vmt33lEWsM9L9uxoi9/gBTo2J2yfG66vErrtu9g3SGWI
5KBzAl45yExX5j3YA2tlhR0HhjQiBuiGZiRckl9PvViUSt9LtofFiV0Zwa3SgT5N
KZyG7Zl65seCfDIsjtGBEII3M8+rrAh6x/BxDG4qudqMyYGHEjLS63p3i4fLR5XL
ytAVrPeCn1xg8/8fkzhNeTA3hAgV3kXZnS5F7rvEsPTt0oO3PrYxQE07x6fih+id
lWzAim9byh2UiUBV7vlVhDIhWHyRtmAZYfqyLvPLKWJzDzTv2pBoKCX0ak3Mpwhu
31ULrfzZfq+gCm+mZ7Bd2KclSL6jBVynMC20gOVjlJEFxigOlfmo6gzurzW2nft2
J9YcU9R5gMmpu2Hxful/XekDR6I+WstttOtCM53rSphGgL41XAvUwX7xE2enmobc
fYrF6S0WEIJFG/73AH0Rkv01nhPZVYLInHQFicyglwGFktt1pSjrPjjLMw13i1j4
KCBzLkwbvlEilK0vFcnUupTQ3XQMqxDoWlMHTheSOSuZJMcWPXc4WUmno3NBSjpD
h3GIEXa7J/DCf4vcBsdFtxrB47gEoGw6NVUd+6A4uXRvPUP/j9HFSUsUeP2SZmJd
By3kflstSyUK9CUSuvTmi+YcDXDZ7JfqIwGn1ZBRoZlt1xAA2MgSPW9tiVA5UzoV
QmV9jfBrvlqrz29dn1swR1HPBQAgLttB1M6gBKOMeLXSn0L6ADHGlNkPjkBNh/L6
yw0Nc4Qh08dYfYpPLylTRTYAGNuiB8HpZseKbIt956Br9RCVJDXnG8aRo+ie+EDv
jek53Sme2CIIXdy+VIwq5/jJybUhDgIx5CcXeJJR5RZHLZtJIp/QbsCw9lyExUoT
3wlKz5pCE+sEr4EbTCWFSc4VcwiQaB4IAz0B9HPBXWcPtv5ZtSMyh7ydlC82kSmj
HHD0OddK/Tu1tN6H6WCW4Y/PMOghDxqNl4dFFGH5eVBxRhZhF6BrIrWIollwUqH5
o1iB50iV8M3zZ13ZYiXXqMJRBs57pz6WdgxK/hIABtyBo53tofuocmqiZtfXq1vy
uCQs41aHW6A7UvZwM6v6BGoz3Ct9Ni9EBvv17EVS9xhLS7a1XcJN1EMx7N2OU7UQ
ZllxJay8FGL8Z3hTfhqJ9yb4ZTgMlIjZYQtwVBY8WAwc5ay4o34fyNkCT9XtNmhC
FbOwebMPWkmAn7Qvh6uMe5SqKVIQYHs+EImWZ+BIPuJKfi6wFDsyrNm/JUF1QPAv
LmmHbRwknzAJ9xRyst7+Tfl7pYUMiwYMMZ1zfmx5SGJvdlQUbOYj7eauWvlnogUM
zM9UzU83chxMXFVGMRb3bBLwUzpYAWUIqDNaO6lzEj7fl49vjxuniW5GUrqzwRz0
vjB7lAVvgAby2U51SfDhDWAmOl40ygn9WgdjmMwvJy9VlsGvvGcp0EP3LEgaTbha
5tMMdLFTEgiWONe6xzIQCGLX4SnbgsnNbqSuU+VpEEoUkQ0sJL+ZYdUX01ZFBAGk
3ubKW12llfq6X07FpamVkiCUBIFZX8iCIp1O4vJDyH7U6sq8ZS4H3+yFiJy8q0Am
mgbW1TJrWXNLN16Fil48ZHHWPv9uoqWwf4Fo/SuQ6FgY74nFCQZMRnw7ZfWbHmnH
IKnNmydacxMdnGcARYWRubnELlsq/fJQbdr6wor5k5s2yPgzD9pKXWTtz3RJlltH
0UZUP9uaKqH7/+eP5kIQP5HJLUtIU4iFVoEAqkAcRjphJ2gjrVv40gPYNV5oBe9Z
dClixtInOIuIyjpKzgj5uuCqtCqWx1TCGaPG5S5nFcB2QSe5MSOiS+1ZAvI48xPS
PQXoekoq4Pe5nj7d3pb86DKZPJ8p5qtvcm2akqFB0SXeT+ysvZs67xZO1HqdORqr
yLp+m901wCAqLXmH5JuVnqrL2pJ3F3W4Kf4vzRexTzVZmdU3QrObs5DhZi+9E6bE
B+KEYFhSBeIut1mm9TVEHBLFWpjhk2EWhAUk5sSTY5+fj2Y7SR7P2OwCW6PMlY/S
4uJuZs8ph1Ah+Uca9T4UmTqXVA3SJmNdJ9zEGj7fgKAuasiT5J/r3zN+aXh8Mmr5
J3/3Jr3F9AokYi3FGjaXUVwY4wcqkoDFlXL7xAaZcPC0KZIbj2c1SDEk5dNZGC+4
Uhzx9S+1GKVpXRbo38v2A/Lt1xns5wbdkrxclRBcosIu2cQf+/YGIxBEWE0xTUW8
UdAodkRD00p1uGqDQ3AYP/JvFmpBBha7iC/QTnXnd/D6o7XMFbr6kVUfCa41hRBt
wRHbE93TbARh6jEwWM4YO5RzltXxSDdQq56g2EL+QNveVYFs3zs2GGIhRLAQtpCx
o3hCBrhvoEITs9wQ4xt0vZbaRX3AWyZ4zqT8hEsee5H1gtrE7KZMzmfdxpytLBsR
qdpsjgL2oVxXqkDgbnHvZ3cZf064KwcNpDc2hohJ4H6mnP+IIxio/QuAQOnFw356
I3t61ucTVBDOQx04Kg2CR9jskCamtu913ns0XkxkgRx+idyWvNOSzmfdcHdeTvnk
0hAygT+Q0sll4g5J/z93WA4vbgxC5hoWFpXrSVHn8s8idDkMLg0dXDTUodKrm8xa
lAr4KSeYPmhrF1Y2gJYUNPLUH9K4mytmQTSFl+fD0npGQnYmN+XfNe2Jr/rtwNcW
XXGJlXhnl30CXwTmlxwPyrnXSbY0tRdAB47MT21TYcPbnl8LXbUU8Nb22C8ZckZl
dcahowKU/em9Zb2rglcwfx9Ezv7x1gicm7GXCbrXAV4ZkcgaSM88TcXNrnltt6+x
Jw126L5z1YY4VoQ5x08kiD3KZTFNt8KhVaVEqKzy+swOIRvbvrxUzP7sZxvxGM5g
PAc3lDPtG/+Jhf3yxNDWT+YJQALiIsxp3oXTil9HdJ+T/4MNPjMFPZuO8YIruaDG
b5uCuBmEIH7qWvyHAud/7OcTF/cK8tHgYICgLQaq47qmVojw4cWtQAUNfGpWcsLR
lAjmVnl4Sj+CLLfsQY2VxDN4R/5iUryvmBCnvFn6movB5Pi9xVbSNpUZ3/MHp3kv
ts/QnZKQAlGlHqSsEHCITb/VCaTvUq5qIZNqSth3p6nt7ePeIVXbeWVTgMRVyWmO
q9dxAF2eBfb6WqtoqEM4Pe5Lrr4NCvvpNStm/niNpur690grLjcEik+b6SH1G9Me
ZPsXbZ4Vo7PdE9rVY9usIloGAX7H41SILypCwOQN6wTL1k7u3mdpD+srO6kDaxIX
BLoI0CLhEn9guJF42PKV/cdLtBowUCNA79Xu0AyJoMJHhVbZjLJDtHGl+FJkCATs
ZiRj2mVePJ9SnBXJ1gfSayZPF/SnA1zYkIB4P8a+/KzKrnybfES53SQzvF5BWoSN
ZmBJRQT9h3/SEuMZ5ZLwJnyV+NqCML+9yEQJmbThOk5Zzunqg79kI9v/lEBtLwU2
eVueK94kw/ZrkihNS0KOZIMl4p5bWvkaLbJ1OSv49B9MStLKjNL3vgyt6HmTiJus
zAE42qFXtUzDWx0vsbi004APuBVMloiyo5QKTjhzfBAXrjJxfzvb4FsxcakjA+OR
wjhiepJXB4DFPRRA90Or1m6mOSpJjKGhhA7fBp+H73o8hXnPBOaEo87swQeEcdNq
O9y0mMqcTqBSneuLe9jaJFeJnEZLWCC7IUedzt3m/z4dPheU99l2iy/hJIoueWH+
jR7MHLFEa+S/hjHHPzvrU1OTxjmBSYw/Gkll7YJsP1u4qeXkQldvaZp2szbF8/lq
j4l32ahSMAbYHDSu+1ClL4RBpNlLeK1kfdeWNze0EDE3h+kfvDyr7zs3DBoS4i+W
wd1ZUClDHnXQWgpVhx0MBFXpf1/NMrBU8X0zbKn9NO4ZLh0Gm2n35zIeOvwm4euY
ERBGiLeDLCv2hWHU21RnMleR3z+CsHFI4STnBL0piIOc5nS2na10B4lUSSgDMnoi
PRiG8FwidV4Ag19GRQcTTj4JHohhfOplniauOVD9hyoKPtHatyIQ4YgFU1cgLYKR
fsV1AuUmt91hbxfBEPrSIX/UlcShjQ9x0166PJrskp1MVHmiEJQrvYtCYWSSyHtf
D4OjNm1b27N044ZyK0/TZkYI2oKMzDamABr01Nor87Y8kET7ZWUTJdWqy10M9zYm
L0MdDycavGtOaJ2L8U79uk2t7TqXHreHWfoheEvLpfoe41q/7jogO7ddLS0PoZ/d
d50NhPMT1aI4CFhSkHFzfvV4/DVZu5UA54+uS4DrjC3K7e8U3U5uGno7Fv6/5DFJ
azDt+BcTJNWFYj6PV97y94BsBSE4MJD13RxlipglBjkZYtMb5HMAJ8ZyK3CDNDC2
WVADyp/9XbUZIKnVNJt8AG2q5c6mZ47A+k26/GFcryDUZI7Yw5EySyhFOCw0XCwW
IkRc6IaOO2ptVaXnMGecRCsqdLRg9ScMiPkYMODqPTvZB7l0/qEJHabbayJwKbkM
6U0HLGbGjF+sYskgC8bLRKjTretL6nOcBkH2/lTreSNZr6T3hAulZLbTVuTX+1Eq
3d7ZGH5Psl1gSEhRDMwU9M1o9SI7/8xGxTn4ljPdtjYUABaEE72Z9nIXv7Xo2TnI
BXTV2mE/Fk0Uqz8jOEHg8+t42J5RUfOBZmdJwUUmG3DrhVVgsoZ/Wk2MhH+G+g+I
OQPU2vJDShe5RCq1D+b3kzHD9GnVKjf9YhWAYUwVT2UI9Jb7+yUNBihn6hAhV+0b
PqkMsgttfG1V4AjcxzX1wYKzqGbgm5uUPcDuBjd9vYzrlYvBs1DNAoROn7Gdi5BO
lG6qRQ/u+SfplW1zZ7q4IdhSn3YiP1oC84UThBAGz5oA2m9C7yyPk2YIegccg9D5
cMgbaA4/gEaApCtBcKCLkOLFfqMfV7MOTeCFogdn5al0OMFToRb+5MS74K3XUZZ2
wbJygFxsG+jLJCvYPsbeWzEg43qQM5PZLkMovOjMV33iVNbfrsWbt9mgs4D1PYlN
CQa1A2JLebGlLkDRDZ/o6qCQQ11W2XA8DByQSBvSS+L/4vcrOUv/VCH8BxdqmxLk
Z/yepPr8wOLbLbi0kJHamvNkqdlY3vi5jk/WXg22eU8LQlb56RBsGwnTMpWTxZ/6
MoAwYW6IcwUsPqvge0OV3aXp+Ai3sLLz2U99BITP7kZjhvB2iX78pYjeddpWZAgY
PhMgfhXCEU19in4AofabZRjtXvT4YN8hqf5+V4RtcT8VbmtSZJ9NG/2siA3UmWFY
cODtU4OR4WXoipw+iNzgVt1XVXaR3RS7KU+UyWTzDVbADpolM2CsKhPnviE0Jgb8
5igYhMQ5+v2wMCrGvwqTExjeFJ4R2QwDmkRnZ9o4z9aLPT9cilq8gfVl98MHAYpG
iE61y2ejwHKSMExMDh/GT2tfJ8Lve5oaiFc2B0Uk9P+oXqTlcVqIs8R/EwI9v9Pw
x4nCLFFfZPOvXu9XqsbNGNEAXg/huM/puOJPy7ZHJjXL+pmnHz60dr4dcb5wHr48
KkPfiniWg+XesXL3uzFMPTjhR6QgIVKIF5NT9BbSEHYrmNmQU8as8AFGZH9wA6ek
pYK8ewXFjdZxmPqzulbUQq0/Eud9hw4RXUySc0yuovgLdh8BHoq7OP+4nKubWeuw
FEbA61w3qVNeoJm4OEJV0HUMaKWEeW+0zM7ah6/hTJlQglFxgRJf4Ea2L7Ab1y4P
SGcVqvonzxkCQKxZ42gyYoWSz1KRfpZ5Y2zSZYnIbn2riWH8dX2ioUQi9iFmBa9J
eFYMySeYQbBQ7DnZ+NcApg2FBRPb1T4peElK1UZrqFb76TMREFKkQxevBe1Uj4pv
81mSzD4jvKrdqE5j85js3kQbi0KDzIC1CsUi8AjKAW0y181x8ZnmYVn8tJI0yuIV
l/6JS3EI+U5lNwkR1a+9j7uwbYlRhykGI9Dp3kX1QmJzPHWY+PS1pVy9K9++xR33
RpIZ20aMKNuzT/viY37zVpV66t5USsAM3RvcaGb9wr+cdSGZdfW4AfFHWvHdY7Fg
8bHJQefVBEi6QSeuOJNpqcE5FMUT0cpfEV+m7VKkHRoYUpGUJoYpfWj33zHQhpE4
`pragma protect end_protected
