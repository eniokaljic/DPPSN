// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fr04b0eYAg7V8ofKm0oDZiT/zNzvJHfXCGv1o9EdCo1ntM/bUCtR35itDdI2OG7Z
bI4EtB9WAmSKzo8BSni1IDxpjlaYeEYHvpmjdyM9GlEOnub1mjE1d5TJ+yucMR1f
tcI3rJ/1h6jbQD1VJ9xdlYBs3s/peMuJPOa0hfZJDos=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25872)
CqD2Y1PK5EbocXnuUakim+v6w/tzhcx2Sk5bwctDp1QqyolEd+8q/cfqlSTpdSIj
VpQIR7gefIXpyJGqeVKsunfz5O7Hq8SgSu/t8fRdkkIftJqn7YSSuRF0jx9ynSMr
T7p5tGY9fPeTCiml2RYO1y7C4ze10tRaXq4yQPF37Vm1+x3SOiZtoW7Ty2sn9/2j
Cuew0NJaC5RJ927n4dcU3WPnKVvuX8etVX1V/3V4WqDYdfrY7QpYtBIbgrQiUMVw
DRMHL/W/eVz58PtID8XnEdAbdd6L2ZoHmsDqB4gWM3FmFlEEzA4ClIQr2uBtF21J
+mTaV7Ubt1BgAcCbwyLQVuv4drwsnHa4LrdUW84XoA/JSzWUMimaMheE94vUITvQ
j0OGmfgsJo7e2Jiv/O59/jxlUe7r+sI568DSR8kUJBTaZd4otiaXqChgTZBtlp6x
iM0lonfdi1dSuSyw813gN6y0JGCsoSiAddMoOnAIZ9E91o+wd2mMlLN95GHMFdWi
pOvw/XKTLVf+FXbpIu03a6OjC8TvYZGRlMDT/Oo88LntZiSP3I8003YfxYwoeTKw
eNQTQBJfoNnZ2PAIY2NTOYsZXW/lODbIbsMSYOvFd93pelDbI2ukBP/y2ZJr9H22
ct3GIav0frtbumU/SAQf9LnDZ//tbBh7SHA38kQP//QfhY6lX0n3pKRlhHOLgQqK
zbwOUR3XtjVmj5/77ZrOfELa1xJq3fwwFXMtWuHXLIqVAWnyU4JaA1buWOLaxpZ8
97iEwzEWi+j5oedMRYSeAGG1i7C6QuUI1eSWtxYnOHaJVOVSF9OEOxa73Y5UmjIu
cIE5pkZhhk6yq90HqHL0Lyj0j4xrsUQMwmThSQD+ARhhzw0pGlpPZf9LAWDR0wqM
Fs8+yXbDADJwyTaQbnqdv8zCWTkAXH+y2i17TMKqNQfNhyt+khjCczuGNXl3NnD7
pHlDXqn6+EsvLuiAHTdjT6HAKLirfW25yvalUcSjVKo0LCwIQGtNnEhl8EOlysvN
6aUvqHvMLwVulS9cLDoOaVOAnjSNKIgayn4l8BtNvz+/65imx5tyNpwAgYl5/SLt
dhfDFUNSS82g1tD8geIHAuORUMOCDWmY4/tFYKwLp/qUordVVwy8pD1/GKneOqk3
yTzdgeolN+BqTSJOK5cFrnP8dTX5xDCT8z5/DSm7B6KtdDmQOTrKJNFcgNDh+j8q
SShg2/XPlo1uvahEGKVNFehrhA2EoOJO3N67fDdzVQB+Ss7Zq+UC3kFmPFLGkTh0
C+IVcSXNnRrJdSP5TY2xmsHyeG2zgpELxxokf3NavM/ds+tChlD6Ea0uhl52PQlf
YypUjq9dqoeolZy+Yn4yeo2cZl1EWguXCb0RQYEkXNnGxWKPu2cJcSGttaFoJgTR
wz74TA814iataIlaimCitqwqnd7C2TmbltX259TbIVC9rHoOTs6JvTS4/MhlG80P
Cp/GcGJ/SI/dlukX57WSdv/WSOHnMHDi7d0eZ2SGMSdItYFn+otybTdVO+a3pzPI
Ls+v2lqNyKEoAp/0cShVy9OhyArxvAzzPtkYuGKnTBPJbBw8S+5xZvjg2o9j2YMB
p0zH7W/RVMHV4YZw7dcrQiRYHFm8c9Q6N+Izw6syDjDG7cBciOngwIrvhzdWA7gI
oIzXFduXfrUAnZMgXhBpA5KK5Hf5SlU1NT6geNoJUrgD6Sj+dYKA/qz8hBdnMWld
rSVuTwSdYnheGWCamTScTC4f1U2OLkTW3JAch4OcW+kAgeeQxC/OwlIhzm1PNMmb
4ORuT7FyH0L/e+3D30SWpLOlXgsk9dCm2C6U4mr8xmHu+VIfgEap5/ZE5+ycGRJs
UdilkLWiUIdYzwJnNUZQl1tptrYpRAcd6m3JRaamsHHOv0yW18olm5/NLYL132ck
a+XeFPHMj0pw7TzLv1x5EndmeuHafPqbSfLioygqX7p8e+wFc6nPl+9IZT7ayWh+
DWGX7CenujdHtceDC0As4d/AKaCItANDQGSHA7S4FxbPN7y4vB4tVzMHzO6r0lS4
Fp/0t485sGjVXlEwFVAL4PQ/CVeuLrHDq2CREFV/xQSTFmztV58Lz+HN8QvflAKE
JzBazC3UaoTvIfN+wGIbOqZQ08NZaZEG/DomG2H4D7yZMr1Bnmb7a+euoCVVOdui
4g63lOQsdMwq50NQnTArhbd3HVXmFu0yFsTvC1Y9VisncG88v6l+VYneuKy9GM16
1tyD5JXNpTd/Z4olHJRW1TNWBncYgzs/1/WgQ9xXoIHmMCyYOlbWIwnoKrbKZZoT
lP/+3Wv1p6vgkrCDp0V0GwdeYdNAuA5Jic8x/US4CNnRLi9gSaOUUBYRQRL3X42m
qilVBqpSDmUNQenSbaASnMCWFPmG07gptqq1bqF26nxsriM5aPSpfaVp09urGoEK
KrQhc6g4uJ0cajhCoIWvVG9B3wjsYAm8tRVOeVUTZ2NU5VLF0Ylw6V/Y8hWgbaYK
ZQRq51l3Xm5qlLwH2LbxDoDCvxJWmnM4YFJt0mRNeGl7HMI/8WW6DbPwF3Eof6lW
tbQk/Ko0KTfrBJ6EhZ5ry73NWAIK12K2JnWk7HscEH0xvq1ZGq3cwy8ujpGQhuWl
aXZz5/sbMzIU5XFbgi5mI21Oaly4b2ulNSUFn4ppzp/i0OUK6pMdaIZIW9DY46sb
1D2Yabd/CIBwWsn2Qvz5QBpKN5LNtT4HxsBlNjAnJStXV8vGfxx2A4pDB65YHZdv
ZEhP1jZ2P1oxn/s/hdEPsALAJ0XgSUskLTZ4w2oLqyDyuxKh1juwrBZRLynj5PW0
LZlamSEqpLBdwDtxPYDLGCcggQzMyrur75g49Uvs9neapk4rs6bArGQiQRi179bC
q9f1ebt0v6gIPaDc/T0jJ520CJoeOo4zxlTnCfNNTaFbIAs9MBEYU5D0MrgwHmyv
2py4SbkyLcPR+ya8ytMm3kWQiXQffcsdrGvyvHVLdflDDNLrADynMDSTD4xWbQD3
IIlP7BJweoLfm9EbFOWnKLyqbZel8JOIuddNtssuzLY1z3RflCy6Wku27aec2R00
/zw+0PFO8iRo3PcnLsf3bZLdA5VH74QF/iBayVYFyIMbK6hsHfBTfwxKoOIYN0xU
NVtkK5Da0hprvM7Mu5SXn3X6b/xtPQ7VVv8S4DJhz05ZLQ+sXYTqb3hHhkM9JOou
ojG8p/UaPAwdR0nGFUPJJh/QGR8+m/C4tkk/hqsbg5Z9FPpahKm0s813xszJBiGK
Ltkzqro7CGLJUPFIEKkEgEg42vZIRhya3aByKpFYqY+ZMgYRfvfEf1TYLljfYka1
t/zR34Ol8c7/ajEsJIWORE3sYaT3jQxqqaV+6h9VOeRNMm7h5Bx4U4lGsZd+ir7a
JSuGC89shjCu3MczUCULjlvypM0lLUBAl8z953JBshkXnHdtG4Hc9yU3TmLI3yGz
cy6fWOLDBBTdrRBWbKg4UFKSEpF2yTm+99/+8ENF/UgnPivg5OY+RahFxkICenwn
+VOP1jHJ9UFnzF7IaYT4KcfzIWcjnocdcyr3QChek6wnQtEdRKSA12O+1AGMJ42h
G65BzO4WZzP27b3/8WTEdC0MM17IMLGcHKdwTUBpDQeCWcWAX5F/Y2g1SNrmPRq8
lL/ziMp8MlSwD8EbywUQjOClh9ZMUwToQbS9S6jElPstZXpSF7/SeMu+uD3cqJ2m
IIFdDBThw3it4vUT0bjjgrJnHqDtKuRMh9NRQwVXPiWOkHq04Q2AihPG9K3B1eaw
/pss8x9yy8l6wVUOj6OTsP6srunX7R4ZgzJezXWdZr3KXd7mPPHP71gsuttBAQ+H
FgIcsmT2RS0dzeD/XXxqmtVcqZzCy3x2+hkxDkAVGNkIPTVHf0z+e4/tnwbjY+zk
KoIJEpjL3aLaKMq7PE5lZUUSSnjP8stoEo4IKuoVxxED4FZDXWnmIw/bM3frCpbp
lSiPTMvbUXV+BosHCdOleOt/KsFBa8XHH4oBPMtp8TdhfWWMnW3AKjO3r6nNWhym
a8aWJbntc/fNhb6NzEmxx3LxeW7mQ8S2W7tN2fLCsZJES1EWBUxBdN0WRiG4X1Ma
JTlpyn//ZsM9RMK5VoRpOKjm//VKr87MRsDRJ6HhRF/BS35oEYUW673x6DDHhff6
0zg1DNVOU/tLkZ4ADdIeUb9iOLLp9dLfnJ9xZik449TJ98ibYAFy4TGGMDeNK3mb
s1/Hwf7RtbRmpMP4eF9HzRnuSGEE51oaNeBtcsg7d5beZ6XHcAzvUeV9zMqRall8
jESXbxf9iAIipnFvC/rCipmS3Q1Ow/HQbMr7ZGhl9a2M+ZilGid0G0CZo8gr2i+9
pOI/MQgiSy0JOhIaHOEpnlcGqQ6hYkW9LSmRzi8iUTzU7k6fJcg/v4IUx9RHT10k
KqgWYQKxdmq2dqM9qK44csMuLz/ELWQ4mmzKi60Apkwa0NnQm4rI6WXwPgRFhdCY
jbNHzFEfjTRJKeLeQk8VJVCY2/A52O6Oywt5/f7Y3tW3RguSMRVgMSQm4hE730XG
FHoyx73p45e6+Z7ImVHwlzy8/jpQhSvoJ1FoukbrvL4MhZIGn8fjRyhWbu4sOe3t
VmZPZhQhpc2F1i5epwoKWWEsVs61eXr17R9tPxBMnXR8L0HutzuHlOklHILW+ydO
6qBR/0INqt7g0+8y+XAJEQ/Lhl740mlRS2byDb9uqdVd9/hFMIIklfsvqArz6usJ
NQjB0vUyBW3Ofe9oUQK+yhgb0L20xEFiKY+n5yQldm0wMi+TsOL+wtEhO0Y8co6e
xrGbq8Sy0SEeKEaCLLNtyNQqz6Jbg9I+CyK/+wE/mLFCAFKC6npiYVc36h2OSz5G
tbFl/32634wNxqX6WbUesmXXEP7OWnw7g8BzJm+0CD2BQK+rz7K/m2VwIWqUK6K2
JUm7mgTgTFv9wTe4xazwpqGu1kI10StSxB/wwyucct1cuXvJx8cxn3aKQCodvXSb
qpaqGp1KS7B9Si6J4ljag3q8n/0XlyFqNTjdcuvZzgvJhuQrmNuYCnzMY9WGhyXe
R5WTSLE+lRfZISd/FpBBhOcpXNQ2Uv3qCWCrM19ARCNx1Lif7iRFNMMz7GTg/UP/
uwIXstTyHpgMH9X0erZpCGKVgL/HSuV8S81jG3CAn5S4D6vc07HW/2LTecfFE4kf
uLk0vIc/NWE0Ly9ABu/eO0a0dZJl9Y2H/kKsR6Y8WXfyKeNXPyHbHMQ/at++E5K4
ZkFCTBiHueLp7V596b1ifVYzR0CO5I/m3XZdvcbSDgEozEHjbpW4QoRJChLzsKjV
iHt+ETxfzM+qOZerVv3qNQMlvMHs5Y87JKDe/EIlGadj+3ooEhhOTPn6wCG24CBC
8qdFJHudgzFZEUIHVSqxLV4+0vdnnBTFZMJ4t7bajE87srfDe510yUFbXAFKQrCY
Nnc8v2Nk2DqLJv9ze6JoGUAMhM9ZzgH5vJrphA+/xIW4/+Sd7vP9N9t8vi+JXrSx
DZjzuwJZwO9Ilrh/Tft4VIs12ptDchTI2AVhUg91EHOSDd7q6Xp1QaLIReDj5opb
a7jY0i2W7+VPqMU2TI74HK2WZDvlbusmX527cKBwiMLyyXF+TWwnS5hE3NZoFKSH
P+rHbLZ2z8rsmd0NjOaC4TPYrpc3cTcD6upiqmyIiYEeKQqwH8Fh5gpHK8OFkT9j
P2Jcf1IQCtt4kH4bfGEtz6DamsHluUQGNgA6WGbyH5QiHM9GcsgPXtIMmQKwOgQ6
gZUFxyiHiJvUGIyWXc7EErkdUTAcgd5F9DnJTW74ABANn/e7JyQVJzrfzKKOri29
wYdY1jLdxctxRb8yofFjGQC3EeiK0jsNE5ayKu0vZhwk/hBVhX8ndVepjhygmHtw
7oFX7vZg44GsXx4qxPTMboJeV1n0WDFyGhHpfoCpdUS7crJ2XU/97VK3cf2Bd6aC
gRrBq9NDkm4kl+RX2K2vhQfsnzhWqGUagCxIYNWc2wWk4S8mSluZF5qK1MabhweT
d1t0U/ks7z9OvY295VXatR2mHvzyyr40i4MBhW03XSgKU1PqewAfKk76ucCFh97g
J11LMwc0QSzW0obaedeQmIst07RYXHkIB+IqanYb4Qyna0DrJK9B+LXVXO0Tr9GE
yHkNGe4YwsFlx2uBpRkJbuquXrlvjT9wMtYnQ3kXM4a+FT2GyFRJAVR696PiGVuS
NKzxU6UV1Ocah7cu0vTktUarzPbGLKBw76Y+tnmzd9+PbHYth99H6N1Qfitisn86
rBKyTKAgM4GJzLax8ZA8du6dgc8dTFHl4wcpXANb4Qe79nhS+n316KoUC29C8MKJ
0vSJ48ELBrOS8KA3KyzR6AgUXvtN57wFPM4MYbXI+bw6f7Zeu8g+XDluvi5nN2M8
Bs2Sp7n8BRkw1HDxA8PO/p6eVNUepsB7wmNNToedpO99zBA3NasOchYLenvvJZhq
8Cofpc0IIJ/zfWiZ89OyJUpriXIgw/FFLdeddnQSU7HCsXtC+95oHzcKV+cQrF1S
KVLF9FdWaeS+iWGaYPj1OtDt6R4SU9T14mKMw8U3truVzbwgoP+HXbeCzYv/e5/q
RbXOTYliGyIF5UQ5+nyHikts0UzaXv5CfHQBIZkq8SDx9Y9rjwMgyMUZsdQTwuJA
X7H35nytY7yVTjY8Syrv5fHW4juqpdrimT+Edu6jrIVIj4ABWGgwI6+bElMOS84n
TWBy5JXdI0rI75TULKoQ2pGhlwgyN6m7eygYRJfKwZaXG5MlkaLtwHjZYpV5Bo5D
FqARyO+5He6dSXhOHdHCyfn3XgFFpK+BHi17bo9y1R9xfLyjF1NPoUSqmY4PcqU3
6MIyX7lTyojBGb6OqwxvZ9OMdm2JeoqN3aMQsWd1nLuedmXvO5lqeA1QS8TslGCG
lA5RwEAK2EHCB1FYmsK0QSGglA35nfVd2H+dwB+6cfWsDsO+hzKajBN7Eb+w312Q
FaHaNMYexNrEXi4XN8PuJp18EjWpu/vht7bkkgXcrJatesYygAoS+h+H67PZoQBo
1gzXKTxpR7HeZjsPtIl7EYsOY4oiL2+B/xXlwyBC1jdYdmrkDAJhrGiInECIFNO5
4Kn+LXtu6cJcoyc6uuKs/lUSjFDmf5Aa0t+pU7cSzskTUrwxDRiR9hdk5s4qXvQE
c3d7qej92HpscW5yL49y66ntf/k2CyT/rRV3WgSPFtFGR9XB4cq+Uoee/CCInA0Y
9MLkEU5eHbfECMP2lcANdEa0ylA3yTFPwQid0PUkG1urz1ytWiKcSxehZixy4eGp
f4ZIqY5YP93+PqRfdprK01C2IiPOlZXnbTNTddUU5n+aNJRVX3gVt4xMdiOvyuyo
V/Mp6tvC+YKoZlP7E8rNQjY6rGe+rdoMji+A33oPvCww9PpKpOLjNKgMmxR/bzkt
TmoHk78LLrKCU3fICkvx7XBdv1JAGtwi5obWet4nzn0FgJY0C0dxdy5lWOi7msBX
dPUS9OkXklkmDhwWuyYEL8ySoHscLrkRuScbSFdizJ09PVZ6OCCjt0KMy+l/y160
tc3tdpbEiqBKBrbp/MX8ZcFRPwve1hVMDKIktq3GU+/nc15tU0WFp0xXcsAz7jje
eA82fRHhOP7nk/y/V3kknRvedAUEUnbhbYm2PoxWi0m/+37FLrvRaEIQKsHHKJEf
ZKeeUSqpVw7nLonA0HHLJIqy+moIy4yFofotEAo7tUcRSoCcnjGF7FNrrWUZbKtp
l0JFx5N/09mGEkWakdiif2TPf3PLdiLTR9Oegnn0uhugOVl6w+nevvq1Y5eIEmmJ
32RfHsrp1XYy+gmV2g0wFfIp38JN66Vn1R98poFx6+cKiyR/qGqdWBB/aXkLNA6I
nKPP0kGVes0VoYzZ7XkAs0XqSbrzQshfxpjY72FA50vE23+aA5hKh4CZx1n4DJfr
YIGEM7neVgRA0sGak6Jsc83vZ6g5+TzdkjHGUC48Rm0awqIEWVMpuSZtsfEdgPiG
BKXJ8ia8zMGrEyzWDg8/2bjPCeqanAz8GG21xLCQKD1ZSlQES2t6JQpmDnYUSaP3
AnGSQEFYxVtZLLIC7+dDLmCRHh5UQeqX4knOzFCVjBG9k7LFZMTG4qFevLlAFA41
r4mZngmD9L1qhxW/7FktCjc8+bDJTdckzjgZSDD6/7TeQz0TjgSg1IhILpfHyPSG
7wD8Rr+6ghqM3wkqQOkq1i6Osp6rMDFhnoq6YBZkGs/EL7W4jaUusMU2OVhJAxG9
cqszmwlq8ZPZrabPC+ZKV8F43GDr8JT8661L87yRqQNHdd+8Yvzvwe4p3WnFX+nT
slNX2+8mvGJNXWIhZmCaagyPTWHSdkoI54tii3Hnpwiz+LSaKncv46JPvbCwCgLs
0Af7kKw8pMmVEMpnNdtCfy9rc8BVvA56dRZLfV1+tgLemRfw5ar3IMHpUD9iMN+R
NaMnh1/UgnbGe7OFTiOqaEnhT2kcIeZlHpLQ6gK/L5bkCfE/4A0H7b7H3Yv/vYWG
fmh4ijf+M8uVS7q4tjFaBBS9zM+fIi5UJI4p5l2EqIbzs94mIclUqPUm5tNJEAA3
90bU8mUBN18cIIIBJETpqx7pEgAtsiAOBGot0hnCMFieyD9b2+gUomjneZRInBND
GNIpbFO51m/zLUVBpRR1QadJVh5wwgEktDZOA69niyCd+xyEQxSqDorFG1JQGzkC
gZLbiKfoaZNc7PljX9YUXNWnWjou0OXrPkjaT/w6Ya7ybv13nGHjUpB5DTvgkGQa
ZifQkG5zV71elnaYsMIbMiXeboV4fjrPpjWQbcA+h2xobBjBut82jY73+icVvygu
Z4dgXxSsuFaRNIyw87swpFMg49xz8Ppwx7DOguMQGblUFr1rjBxfObucs0k7yJ6w
HkztEgWcogPB5EI8YJ2pzUtsL3xcUAT6LWYEA4UFM+mHaI5KI7AKLmJJeduHArb+
RPIt5+KpsuVjnMRrfP4MzJpyTv1nir1rmo9M5t/sOGfQ9lZOU/xG+XpT268AJEfS
vWBlekePV7JEWtF27EiI5pxvvS+wo+fcOL9bk3bd3ax13x1PeC+H8D95PoA6+4ng
V4upRQNwqdbPZU/RMA7e9qxSjyLzS7rRguDVu+dNvjL0LMnU7njdDXuY5aaRpAvp
T3UBb+P+QMiesOgV+xT9myUYayDgFsnHBL9C9pfQ+nHr2bM5TDX02PSh20UmOc2L
9sUTwbXxuq9QL4iaXqyeYpFO7IfBhZU9wR1CHl9gR6F5WaZ1mMOsZ1TCldGdl46v
IFNx+V73LV06zcXbM3jZ+swKSqOxNnFRpVBSklw08VHnn5BrFogTfdnt52JVPhCg
0ARDBWDzx+fQvn6RKkQfFeBRVcXNhCnUfSyrXvwAvgYCH+i4a/kvP3XCrEhRGQ78
lWHYCJVmM8nj68LA2nBICcEHLjGwirmpWzdXnF658kvG+3HEfGUmDFds9oaQxtmn
1QH95AVUlSLElmTht6pjGb2pxVLA4vR5BTQScG4I8HddTh93wtmn+bpRg8BxrgbP
v7wAAD3JwqHkfhwgMlImDDljIyBXk7n1iTq7NwBBsnK/VUNIpOiDvC1gd+jTV0eR
iJHXnt8hJXOIejZl9SkBYNB5GlNW7R4R03wadAnJcUBMC0GFLP7AiWkAbqgwZteg
FTV7bWmAJvZcC+LzIosiMVZXl1Bo+OqASj77rcZbMLW54FVEuJYU+jvYdluGOdGM
Unk+hPRby6NTSQKZpWZ5t5YfmP8Pe3al7epHQ2WFzP5WZh59suEdO6IRRSBfXYX1
3CPMsrI07ZLmj8vb0LaYFXeFowvyS5Lk1udi5mwqv+Ls4cqpvBlD28KK/PfAHCtQ
s/KbNj3i2l/5zTZZCMmkNBQB1iJ5kTwjNQgN5NpV49JjSJDaWQm/Y6OvLvbJVB17
eNLCjVf+6W1hrI850mJnY8L3BKgGDWYiFgl18LiIREpKo4DP+CSPL+3P9roP5TPG
WyZlUMGv2sgOaPpnYEnKOyeS1b/uJKMaSY4ne8DsoMiq7U2vSv7mxLy+9vDb3m2e
knDB+zy+EozdAd4cb6VlR3fLJnC69jfyv+IWDh9DYUVY1yTKoA+Z97YDZ9AOWHmb
vuCctxTd9gdsy6TNxC+GggalKgvhNvsQLNamze2a0GPiuH62wfS46BFqRPBSjr9z
yiWtUspDz76yW2Yh9blgqCV59UptuIM4DfhYr2Fv+ULHi+tmn5xp9GqLfmo2ZFuL
6ktCMsgUEnXuze1TJTsNTcxvQ/P5aWWyAKpvcqww40GpT1p7uQN+pX/me9b1iTpd
55IkID2txPeMz/3EjRUzxma4gkqKA/6hktZvv1rQFIRfDOwXWEs8KxgT/tmo/eY3
KlwYnSGCsNhd525KWEmopZ9UpVncTo3dGzQEqlDBwaFzF0+nuVGw/GfAjkB8BuQC
ZNGH3ljWAdA00rK7dzl2yzDTTKFTnaKPdO8JLIVbR++0nkrdy/9d7sIxMoe35+t7
RytLnRshddrT3zo52PiHD0OirBrYv5nYCZCiayIchj0sAgkzbTRBhx3pfemX/+mf
wXUMR9vAmD59+0tswQnxaRz9sVDLiV+29RFdrQL0rRnrZgTFbH+oKygHFlwnwcjA
INLkKHOuW9MdoRLKVzG5wUUwDqz5Viy7qHWh8E8R+QaDS1A/X+to1yLDh0Vo4Lpx
LSTIiJZ0g7cmrMjV4PNP7hwodArvJDZnMF9ejIk3tRPwd0b+Qi47x9FHD28AYuN4
tD7mOHeM2bqHmZiYJhhmx7OV7rxt5JGvMdYhAcXvYuMz83ZmubvwU74W0HkftnaP
Wa29lh0E54VnJbS+D3muV9cudsbEwRqDYRcXCgy+K1FE3nuF8lUIwfYx71tX3Do2
JBH0hjASDSiTvcO0xrjqJ6bQd8fwX+tcWRDvx/+my8EMdpK4Y6SYUf28ErusYsuF
+8mLrU7eP0vFwQbKX8WK28WlbSLBGt3x5Xfqvr1F9MhMQn2NJm0H1knUpFcT5xXE
Z1WhaZ/fWP+xKzCpjQBEP833/UjRh3Va/w/naanPbaOA+g9VciEGBBN+U66QKrXe
eBg31ji6tz5Ka8zmFk9Mjy7G7UMO8/mex7rlUmcABj0X8iQkyz5AcvUyYOU03kgW
wRX1Ex63PBIklh2/2k6+nLu5WuWYHBANWXigcHNlkIUVSGXspNtd2PLSEcsLzK3C
TtPq2AUcxvU1OSmZo45gePvHVEKEkSN6h7ppzdrqFi/Ie5CfwepLLXjXdrTyiMYK
YwfraMTjeJWOaxhTcSsuGEianLtDld4g2gSW4DJ/DwFSxa9M0s4+D1MphAZWEv/J
CceyGRfpjRKWqvmhH8iK9ydiy+RpWvUuL2g60AEYvHvxU1Ltvrr3BVG1TvKkuY0b
Ia+Ac95xbmyu2tWPk/XskFMkJI6jl9kDSw7Cv0QucP7SPKne9mKmN7X6knyLPdhn
nIgdTuZtxVCCJm6zKjHveCMr5tzM9JlWM7Q2dQGyOrUbpHNBzVAihIjloazbNGFy
ZHpZKs+m1rjZHyZy20o0wfA3IqqEfrmAPIwjWjfxhXovHEbM4FZxEQJoGrL5QdZU
Q3MAGRZjO7OZ5qgvl7gMOQgebfLzkmHmZ0dLVX3lblgqkMHToI2uhza2X4BhgcWv
B6rcZp0JFefIVtDPq60mOGHbmqbHdTQZ+SPK49TsxRIHB3CMMBFOSaXECZAIT+kg
Sw36oSvYl2PQKnuZYd7KiOTKBafcF01LdR6wMcbFZI1ndqO7N3sGDvzktEGEXkLV
uYFr7Ml54nrSOuIuxx+IX5A4mM6Oh2Fd5FZgzA0q3pVuziIDV9+Ky9O2YjfD98Zd
W3/rzrEooLMHvPUp4glQJ+/IATD0jifn2yecVKZwX/Y2CKT5HMSpiUpMtFDgfVkp
cT25uMHLlG4+lEkHSgFFPPA8foG2S150q5AAv8O0xBXNqsjxUrS+oe1HebcY9KGl
XbuTZrCaNAsPf1/8jrixXksAHl8dZp7KOF6Lvi0qWEFXAuBGYTiPY9+Jx8Yhk5TS
ahiDYDzWWWEY8igIUnRP7OhTECV5TUH6CQzEyyjvsLu+qHDHuMvKwAarRfru2K0y
KuP7EbE0+MbZiqe7gEp15FH+kLSRsouOSgXQkjgt7FWJ5PJeSPmM4qy+33ONkUcF
8DIvMiZLrGMPNOyHEv+j3NG3QF60jI/Juk0mkv8P5K6dk3bho+++AlIzYCngwr1m
/3oe1+4ngVz6Ru4JH5ZK7RVlr2GhF2QWC6GJPCUS8avS9/F7DW2AcgcCK3wMrY/9
ue4Ohs4Juvh4+HV5lyKetPLlK8HhG4PeIl08uu0AqU0eMOu3I0I9U/ID4vgUepKi
2LVYYEkCJlaBFAywsp1SROtOm+f26D4T2P7ub01eeBgX8G4N4UtZtmp5WBcdWWOM
f+o05sWGztHt5dkkgJfgmp5n94WONyeWDjoZ9PEYVX+PoBD9R2KKOniNNSxL03i4
gIDjzxI8julFcNagYJsFJyJzdl+icOfIAZd0YH294nImRbFOOO7MritrIHfBOLSa
FFUYsV6LE5x9Udglg+Y51rml/a6lus6xRn0j2QjJv/WPZcluNfD448nJ7tUHvs3M
c31h4IuKHtERjAQdVacM2g+6omEX00h3hyOa96UsSOMB+cFWLdBAWI7cfel8Vbja
f1JwQ6yk0iP2C1xcHgc4hSgVI6pz2hD8YErDRwm2RtZTuQUP4m1ewbN+HTZRF6tx
rWja99EIFMqWTeOKXWoT+gicadca5bkIX8yWT2RApPR9xcc0HrcG4AOuVMndXn8D
Q5u6pci6h/315Nba/HFDOeGad6X51jjNSJJTFPZT4EYxmqYvg+MZeL/iOD5P+W4U
nz3LCu1QfWxuSqlIOdulws6rbvTQ4WP+cTVuWs2g140V5LmN25j9IgoECajWks9E
D7/KqwXHCLxWOzbwkbmUpYwvN59mPo6NmMGhobE7TmzOriOwHU3kNjslMV4p5hXU
Tq7g+YBPYXoV5AOcUwcurl/SGHz/9HcO1mq3jboQMFRPkcd4gFtxkMOgkxSbzyAd
JoWWrJ6MsyQ7ESVoPJ4o7SgqD+74FDBsQFceD4F7TftZUOY+SyaKToYnvG/hOrQT
yia4Tof/8L64o/2KrdzgGVYuoru1ZlVjgt3yIbQIQSzcd6OWC51S7RFryAZXZdKo
ILlGnoOv6oRs4X5X+wpQTrwuHA8vlGAdFKCp9csufR46L1AQSJjTweJkn0kUloz/
c3Xx8VXI0hmZ+Lrz8fHwCtE0uF7oxCxDuzzgrNqSWVUrvZZc9H4Bca7jfMRJBhJ4
Gz8LpcLzeGkJ0Pdh4upSwnbp/fk5cr1BlxvUKpGMhr4+7einjNlz3OwhjC8I7Q1E
JNytPaLDFXD+GvP5QeKkBPZ0FDmKKq0LvMG8QUrvbZ/gcYM4kmy9wqzIsImZ+YnD
WqyOtLvD8DPmYh2CQBhOX5QLswYxbGiMBmnzwG46I/4YyeXU4aYtOrCboa4vVESK
dvMfYb1uKMvHu0QSMtpXLxU4OvKcEV3VzFN4DzLCm+kq4tn6alj5JFRNvtq9ng7f
UmXLxTHoTOfyP5vIwWn0VL2j9ui45yK9mXeCtKsgou0s+2i055Au79ImjhJIm+Ms
Tho9hIqKPB8wOgJjH/18eEfgnY22BFL8WKYEBduYLt5ONA88wS0aJuDZIqpmfclQ
22UdZT34OZOuoKor2f6f4T1eBuOkRy0odc48b2wn9r9e4KpACN+6tXhVVURdYCJo
eZJ/2e2mDlj4q6pvHUaoW46AjS4QVwammtXeX8P7bV+QEZTAdBXZga1FxwUQYBNR
3ghjLbOhNRFcYZYaM0IvBAxYd4riJZAC1JoP8TsG7pQVUMn7OLeknr/uYLRjfPZA
g3hNu+GAM7KN/5odcwSkykQY4zEMO1P8O5l1WsSARTZbwdOX8zVbHk2Mmmc5c4Yf
ZIG6LrnAYk/tLNCr4pAP+V1G/g6JWR68djnNAeQSlQptG639GeHwVG+HlhAMzYEr
uZJNWE2sY7lEuQV2fEjwrLR4EFA27eqpdYr3rSOaCZCgugelvaaTiz0ORu1wgU7i
Z1vUOdgtXEyBA1hvTjxIwmZE0kj4UHyi3c3AfmtqxHvxeFE86SyBvNLmGazJ5pfr
UAhWUp340QA4FuV3Gyw7HzkMdXklk+sE94faNXAfDOig8tJpPd1z4bpUZ//jc4hZ
a6BaE0xMBneD69caZcwrshwHqzATtO2TB0hiyldkMwNBV9HF/zw2vTXulARXx8/Z
0x3ULy7i3C6Zsw7/rKGzAJh1BdGiFKGQG2zFxxPo1IodTuCH9EszpJcbQoNorOha
61wQ1gnUp/pPM8GlzAD9Y8AVVWoYlgsZQnNe1R6nC7pp/S+3CFTSToUiQUr8Exx+
2NNWD9enJLsrAWmgFr8Ar9QgZA+drKQ6qZHn+kf8Ni9KI3tj801We22VdEhSznp7
M72wHiKBuYf0DW2RhYgwPkQ23oxVWpdihkG9a0DmpuI/mmAvXzdJAUP4SGE99UUD
O1QvyofGRv+WfV0PC7xzeYXoFCSPChHGUnNYO1wY/bs5MxruCbc5irNvtr3idoJv
5qfJD/7x43etWJ+1IBDHMa2n+n4JCXpoKF2JEt64sUn6I1ypAQ6KYYAb8ofttVPY
P99z4GplgWfGrNvNmFsS+hga7P08ga1cxAIAbvwEB4q82a//4+6hTgyavAl29gnI
33kcS/tRKLRfCAq1IJJqOsHxuytFikfuCZ/stzkQuSTANJ//gx9WZdwRLvvIfa3T
YtL2Lw2865872t+EybTXAvIyKYWrqCsJ1rvFvyj19l53dSIUXyrykc5qDOzV8sNl
67uMxDfelMU20DmVF1eH0XJ8/A2bzArHsA9/dlAMnW+CDVxm/L8OMMWhzuLvHWqE
390sJyDWkD8YmaYO3pWRFN1fFswVfscLr5yPvgH/G2rFYc3uXr+g8YI5q0H77Dzm
rt9IaYstE795MuH8ihjWNlFh1EPFzextEOJMaVNP6ry2Bx72IcDYKA/QjUomYADP
PW53yN81rGxQOTh/mUeY8cstocRjAGNxdQvSMgPCLNSuhdFxnqZH12CsHoCRloJu
4pByDdhKF0ziTS5mz9XHAEqRFD1pFbzYgA34riZIht6kjj0Bnt3o+vbyutV9vQG0
Ozprau36vLjiRyygnF2pEnMvW7re5dm5/Z6zMnjUzDvXmaaQH2PoVA7tqXdapjuG
OSjcZ2q4Xa2HGycbXa8INhRzf2uwgzOUZ71zj2pJgTTOWUfUUp9XlSRpCOUfXw1z
QFZg4Lch929EE/FvXuRFE5rAcLU3Aq1xFOovq7kQvkduXY9HXF6oL2wVB1PPnuIb
82T9/hffXTnRuSxhsVj+JHtvzj0wq8rruRFbuzrXsDIHofQQKXDPtkMrfzEVsfPV
uLqNSRAgI+efccRrbOyDcPTiMJCD+6ff6o3duxD0i2Uako5wab/xCilTvjC/Fi5X
Rex5ksZHQUnHB8jztdVZFXYc9w3wS/5CcLifRhLTru3xQGBw2jW393jsMIw9g5fM
S6/GaPnZM8se4a0FoqjfIetIbBL0/jG2E+E38tRzv/YUM+n6dBtYmNdBvPBjTLoV
UQHEe3vASKj1uRVJWRZ1Hj+pAD398vj+aXUmZ64tGgoRy0i0a7MvZIJzoojS1cXW
7bgCMfPkGoVwqLR8VQ0xEWNleClRaxLvKDb8y+WDn2lNT/FshGnlquFBwuguI2l7
3JohdOUeV4vg6vfQfyOK5i1pp8V76wR8gY2T7dWz1UIe5SBga+Dn4L/enMmjGbaz
72bMd+StUljSj+aIMFg24wy2PS6wPl/Gpu+wNzFj2DKKpz0YhdMt0KSfOPFkPvr9
287yst1XaqnKLpid9zhgVV4fwqMpMHb4HrMFCkFuXu7ckmjmFrt/sItByU1pUzJY
rbYcJPqKBCiiom33qrrMjgRmIRI0kAZBG7F2Bkc8gwHI9fiTQt9f2XhwXXw7yTWc
b7GNOlXMwlX4tDuwltBmp+LQcw+Uf9QLZKy1I3TFy2HY6QQAIEq55PgQhaPgRLBG
2WXKxBFZnJ5T+vd5WoGGGx1+H2emSGV8E38NB6w5sPGO7mRmLy+DKqTYx8wLTF2H
ub2p0xQfoWA6EYDx7H5QCLu5EdZZJlwY3vNC4PAbrxyQCEhYAfidyK3u3fZhyL5Y
Hss+oE1MJArKKIB9WqNwaysfqCmfWRAn5IC4VDK1kmPW1Bym4R7YxD43kJdlTE4h
5SKTJO6Yzq8VYy5g+4pPmVOMYsG8yUAhhO1d3WxCFqrQwTiXHaJs++WRUIPRiA91
o0OQ8regsbZU8nRJT38WZqD541Bue3cgIDYIAncUf//EIOeJj//5CjYShV/d5Bje
4Id1qCeYxqcg2mWeBWQzuFgdNAzS5WhuKZ/UVWUY88OQHSMufXzC24s7uIR2RQn3
okYvi9ec+tyre1Fj3qOZM5kfCvapgS+0qDLwWBTmwRW8AAmaSf7NGgTOEDPdNutR
ooyX0rcmOSqWz4N4E3Qin/HZ9nYG8kHahlx6THlO8mk/Pl+14bmzbWlu/Ehxgqpq
XkMuPtzlJ7PfEaZuo4o+DKLqCPaQoFTpwQ1cNANp5Nk/pW+PCZJ28tOH5+qu0I1K
lwVPyciB/hatQByz8tBDGWZCtAmPg943d4qs3oW5ID/DZmVfQvELasb2c1H9NJ6s
SciQDHPS0O67IXHqTDDMfKj4tyE021foavdNjZ6MgLHa2HZvNn9SfVuPgwlKGbMf
Lj5jCCRPiq5/d0dvK4zQlxHdAjcG2ljWiYcqy+acnwASkw5kW4ljzyj5PD9d/VkM
FN89Ru/aP/h5NgLxtPavH+ynfcvUtg5KtaEJh/NAWK1jTYMDvyYCV43zX6b8NNgh
dCYRDwOCqlqZfkTfvL1S30n/ygelFne0qoz35iGQwi0BHpZ/PGCtAKn+jpChkr/E
oPB6DXXU0ea1kmHKnxGYizeoItOARiUDNNZY7DNWAUekX/KyABTI33b+RfzY2Zhy
X6ahhcvCbvgJ1ujEJStti3cs7zDqejAwq3qYBF6iI75I3/ysAwNrFdvp5KLkFn7+
Jv1nbfpmmokw/9FOUCPCHzJgDFUiraPIaCpIUbZMzZ+AX5ELmooCR4eU+rGoNSA3
/auDxY55g9hG0wTssXmbM4E3Tqy/FpGv1kcU2/AKTPUI+Io0W00G4D4Uf6EGUB1L
0GAeJbCMNGmwHk9X8OHilkBrWxEJtH53q7G5cauKDBkPN6j9CaMHgcm/fcGj+KGO
l1bWQk0NiTFSMRDHCQu09VA22e1n1LwMyLI40+UJv0Qyv7scd7zjwMy7LCkPMYXI
PAdXpgQ3B18cUpWFWQMVz5SuIP6DGS36STfIC1dv+KOwh3ieGWR9GUE5AwDUfquZ
mQNPmWgKOMimRB3hXXBN3fv4oM/duTBEENpfh6tR/LFXEUGjlRi7uSF0I/FnbTej
hJVovZ/mCyyJ5uiWYJsKYnPdMyA8UQAFqepN5LPVoZAKx587P4bwSZ4sWcM0m2d4
vgAXsrjNgjEQWsDszGCEGA1qRHlwOepquqInFUwwnX+IbUotTNiEaj6f7BvVbPL/
P/AFC/1H1DOEwS74gVAN5MTa2koVHYI/3kC6+4cqNBxwmE5h8lJeGtmgYwnCsN8P
sY4PbjMxT152Xx3LvG+FSaYFgcBjeyIHRasJLPnonC6VuGSehZb5/waba3r33U8N
wJgf0GErPwvPuuZq+0OUBlNK1ZlPxzNAaxNaFV8F4cqw2MzWJBzttXeVQUNmHuWq
0wo5JVdaDGoWVANYR3Hex47DivLmp+Cg5UjA3hfa7cSNYDhJjQFHZX4c3/wcEZrx
ua9HJcekiCmAMSmyo3Hgmm1DLBtzQpD42hCiIPLd2f4iRfJxnVW+lY+SF8Hu66K7
ZUXXkCAaAlzud2Oqv9jp9e50/O7lZQN+CgVr+dMz/a7oFXc3X886/JNSPrOak/Km
QZosnkOMX1l0rC0AaLgsVHOWkhxF6LXWWjuh+g4SzOtZQ3jnhn7+h9VekmHKjBn9
5eoNCFMLBdFVy+yXQHqSGvNiHn47Ssl0UCzXq5Jr8RBRohhZ4gks18skGBbiJVRm
9fwkN7kIvVauPFHzTS5T/qrAXRqQV7ebQvKxo92o5X7TUjzj6jgBo2QauKkk+MQ3
aXbI7q/QKtBh/rPmjMnQneDeyvmaxFfKVk4BQKFB3W5+7HLcKYzKi7MOwLnFsQ1k
DU7dacK+lsVxyg9nLqkdobFHWtbzQVrDlQxH+l+dmkqGgSxydTUxDaynV36OeWyR
uhL88LZi7hDXbSHPgfh14tP/q7XEYeQ0xIBFlWQrRgGuOdgJQKYN8YzXHwj7Wmjj
bwqqe+vKAXrYmUhvi0XomoRPG8mp4zgWJ+7H7KPcdRLhQiLEw73S2dqbnfDwHqdM
XxNXxx1eZ276NAdWqGV9NgvUEN6jFMHP3CUVirnmrHpCCZ1WzPWAmRpiErW/Vb2z
anpH/QTpzcTqQ0GFRv8TZcGjcRN7t3LBiEC/nDRE2B9IvG0a96XhbTn6NZejBCrz
fqtOmFMPFMxDvI3EdYQUgKZj+Tmw7E0dXhznpznV3NRZY2bsprJE5UegdPKEfbzr
PNMscfftT+KZf34I+F3kd6L8HtGuS5AnFCjbOWnCjWo3lDrPtFihTKnu6gsLK71K
+uK5vf82rfzsUXxYZ1Ukh/2KJ9AjT5JXVkfIe1jBAK7/eSe1NQ+Q4/T+Qd3AGQ3x
G1ccceGgs6ERymwxRO2ChM2XPW+sl1ZyQcPZ7ULZnu+SCZriPjyD08Tz5PtFgb3N
dtEu6aFVjP6bJvfdkjAJlQ+VRf3CrySQQ+DXDiRti/iLS1teB8678WC0XpYxmvm9
hIziCYZX8BWnWv+03xon2QYnSCBtOZqW9tgeifS3+YOHbAFh1sX7UAqYUYUhUaCG
Z2c3b61sB46Kl5PI8ChzjAbYs4BDQkfqEK518oZX7rs4GNbtx54KVKR0zs1/Fw4a
qgEP7BTJb9rLWpHxzdJzoKhNl9PJCoU5q2ik3Z2XrWEX5tBXSV+dP+cZCdfUNvuH
2gsgWWuJ0WpJn/XtM3JGduZCJetvdDxhVPNjQ3BxvLuSigZaiX2GShRojHqZ75Nx
CO4oqCyAgmQcDaYCzRtmC6zQt8VepJCfee2HLVz6G3SO9Z2fApNHWHoxPUH8A8qB
3wq0okmnwRUj5VbNhXs5SOB3nwj3hL97JPjio2FlGVYEhc1IRF94U3DC1g78Mfhx
274wl5uYsxKMJkRlEBShyDF/9QEmSjqPWgWgZWxZb1a3k6zmdz7v+scTvQiSPi/L
OZ9dJx48TrxIH71F9MwEytXlsEeWHPYwatplTV3CXOiKiJDDj3Wn4AgdsZoEOIIq
5m6gm/Kgqoh+Nje/cUiAnquPbskUNAPspFD9AKL7hx1+bIWRPZzGHz67O8z4jaNX
Kyft88HvYSKMeJ0RcygO5Im8U7p8eltiieBWS6ZIha3AqenTU+68JVTw6H7+enea
M6qPiti0NuNjdHsCcLx2DtaqmBgqYB0RNDq5IGqa8oWf7N8xwAq5AQ3ksGB6GXrR
Wih1vEjzo088/BC/GyjAMXUiH9OQsORLOKFt+xU8vF6nYWG8zaLntG4oB7m2fEPm
tEm4D5JREKuLm1DChiBrhDX84xYr0beAdYiriseB8qFi6fWHOh0fXxTpIojnUQtd
a1ev18q0f41tfHC9BlMLNq2YTASJXtFtilOc7RdFA8OnpV8Q1MRn1ZY6URs7Esxj
h/BXd4+GXkjblCO+tCs2bU/Ur8rrXPzLC/mTbyx9CvQ0EFvnGlKN0N2F7/i0OJqg
3FR2Lhl13kHntHYukZNNmjVBiUyT2Le3sJ0C+ArN+z1lbogztyXux2n+t2/bieds
ZP7g0CT58jN7PQHEI0/u5tp1QTpaLLc1HBwSJ0KbrBN66okHFMFU0GlevMoDVCd5
sGKj7pmwbPCH+yfw6whgaaK6ofT4nhlDzg9NyWpq2YBrRJ31CaFJRLt73XFflgBb
CPdwwqZBtUrgtCnx/ewB9B4i8mCMAyHQKdpE41QJlIhWYmwCZF6zSskcpCDrXuKV
ML/5noZbr3bIp+9TJ65qlKUYArgo9hMNOuDwqJCvkwR/I6Ce2Wfhp0iY7WR23c28
imiDdVZ14FE09Y1cTZl/FSkLPeUMxwRPqexXcUZMyO4KW9/bpZnrPie/FB07hCEj
3vyTrDBYB131pvoQqgLFscUCGCpdpPNuwejzvvV+1+SfhXengHS4GUfHDUGiNH5x
Fa0eid9d+L/QOsRK0icytAEC6j280FjnI5kFsSW/p52yJ68DXxIXTUQL/t9CbvMM
oEnGEjbocPirf4zH8RdKOqyLykmDaaHvcj0EmMzrDmBwOgdBtzk2Of9wZMuSy7SE
KJnxnCHCgJyi23AAK18nPUX/Q125tLjkC0ZZfGEYa5b0i4WvYf9iRll00/eLHnLv
22WBlvOQNikw9MAbCh1ZVS6PFNWrfWLnxGlmv5IuFm5uFJCL2GRhAdZPWL9wpTuL
EkL54DosMMgLWsj3Jetm+1nZZ/mUkTnwVahOdlcEMDLH/ynsGTpUWNMPCi/J73Ii
OsiBJGeeQagmdCXH2Y7Ucrv+dNKYpEXE8zIaTWJhUecNoCP0nMcUYfqjiUdQ5rly
mscZLWx1j/aTiddf1WU4uCIC7QJkx9Ze5dzPXFcX1wXI3nsIFUUG/KGkiUKEWAuc
YCreZfvZMKCL39K7rQlrEzqgDCNYBgxE2iMN4hSuEDlRFb4dV1SXfLdUTrUd3dRF
jWQSD8AFvPUfw2mKhLRreidRgWtkh06Gl8yyKD1ByuVmzr35hXu1sfQktELG5ZUE
RiapNTLIrvjcVKx5ieFttuIlIkHdC51pXBLUSZO7nwHFQRoGmFt0NQS32E+uqbCM
r6UOQxdSFO1dw3wq+WwsK2UXM22QW1iTw6AEcXkMFkfZu7NMtlvVl3mTe7cyZ01K
Tf2JooGfb47p619mAOe/O6oN6mYN8JjnDa1DP01OjbkYHsZ90cu+v+bWNuCt/qho
HyOzxMY/nQdAOwxsYkJEifYiYb3CKezeHe++7StfKuesqO3ztlff2zsdDlmWTsup
KnPGBWt2gefQkCJOa4FTiIAUe78f6JqpL5wGvTT2Jz8cXVYMUL/YliFiYvcYdYjp
D9rvEMqcbTa0lj34Cv6kOufP6psMvhYNLG0gB3O8C5jD2SFwrh5Yh5oj3K+zod1h
KqmBHIQhY+2ojvxm3aC0ojwQkhDRPfybuIXSAS5gPorC1YrONgkgiraJF5t0TRPe
RgO9GsfoOfx3pGg8o4sjwFAc2IjlS5o8mL99eKYRBQPQlVF80J1QFjM0QzaX8Rt8
I2623fNoDb6s0hLaMNfLvcYPQpxN1A4I4upNj3S6P8iNfdD88/g9IZaxO7213CEF
2GYcYJed513VE6LkW8MCr5Q9mWTjVdMkW6LA3ze2inZM0W5eCIFkHJBaLimPU6Ol
Zx3TQeUSvsMczTs4Ig82KJPh8qteaOneYBYGX8+asv4N5JVUVOtc4PauB7m1Gi8L
GLt89CyvhKuMgj3mxKsihLlRFabQM4vGAf+WVw3khFsffyYcY0igg0SM1c+Y1S0w
AjIWglkD4P//sP2P37G/HS6iJWWvnkfUbGO77sVeWo4lAf64j6AXVMZSUDpjWPqN
+XppEntlXJqQy0Ao15SAvSQ8ZCh12bbb10FHS64jWU4w7jM+UXL/i4OgCb9yH78y
lcQoFyfBZyxhFUo9LhMftyGLSREt6IG3TBIaXIHvnlsrKOcSSA/cdruj9nlSA6y0
s5M6PXwJHImRuhWtR2DICoAgiekcaexR7aS2runh4SnljF/oqNo/LU1tEJmGzi8E
gGuFWdBaOaw+/TnoIvG+zQTkfbCJdPSQb2ooaLVrLy84EdY92yvhyujI8L/JI2PD
pulwQo82abm7/4Whb7qmqMTxYLOHPCst9TsmEyrGrcIAol/gjwzmaOXmWHe2gjz7
sOaXXzv50xPyDEfu/rNsoAzgOwR1O5KdMgEBwmizmLOlFsE21IinhiqyAcdKvk2H
n4EAQ8iHsOvHe2GdUeNb5QUceKe51KXkvT4dlZ7Fa542pk/TGVNzGRkys6w/qfwz
7P9A/KF8NS/zI5eWcO1Ez9HlzveacaMbx5NRy6fiDuwmnc0HMhP3NZctwZKY+ZpH
Hlv3RcoVtzLm+P0iq3O/u1v0YJ4wAdK92CjnVtiL0frSRzHB047HhFgsbbKA5Sjn
DLsJMdHgp8jXfVIkElDbvgQQ95hI241lXfiGGWm05AWAU0TmF6i5b5vs1nLf+ijB
GAITp+mFzIW6/tLgWlb4qe43hoUjpKpIonwme04q/KizwrAeqUWoSdHy0xzgWbzR
PuZ5YBXqjsTQs+g3uc3UiuxzfP3ff1N4dTjJCjyVMu6ru45/IxgYLysM14Cw+3tK
I4/9B+j5C+XVcCnKtcVwHTwYRZJG9zBjs8qvc/e9VlkgDKRNwTsF4sJPsCmJNVjN
3yVyAhkAb9Eef9lAlmQSjeGYPz94oVaNju7yzAHXszJxRcs9VgiRnSnHnrzpl58M
8cfMQryMVb8uMi74v2cFy+HCiUo9rV8GXdy1RggSUK1Tw27QCZTvRJVx3uktpEJZ
zHaXMmH6J+pXL/F0r8n2NEdkRBiCO2Tspa31GcFWDnEVpI0o/0gOAtkxM11TlgCc
P6JflwQlWxNiFo4WvpyX682Z5FCJ/X9fsXKPpzE3YAosCLkMWjhgmmnAMFSKzLu1
I04PqbSEtQRi83ua3wHlGQFw8YdJ6HTmZgO4VmhHQZGDLPkvlebnpa6YKFauZcHK
cCOZFWGCqMn1AEGl7HiU4hkNtoto2NPQ8D6J17i8u34iMgRNLNNM/t6L5zrDR1jJ
EcyZdCCqH0ptdPTGNN922a6nBUlq/SjpeI6MBquokKbaiZvS0rR9Dk3dY4J/oeFd
lvpme5QUl0fAK7d5zGPRQGnjB/n4QUF8eleDUURk54So/c77WAkLfMnSXT2zHog6
z110hEMS6575A25ubHZQFnIj7SNOlpcpLQerljODtVErPFkZ+NJPEsQge0SpxmCo
g6r3bc/x3DWIltTBcOZCBaocwd1xfpnJnUghabdU0UVPxdTKUOZv4fotv/JBG0br
VU2Vfb8o3fYiiMONfjuiVIHXpqulrtlKux6aEhsX2AI/42B9gl2Uz7vKbuK1MU84
DG+AK+/7Wa/sqVpIPGCrgWVGv9M8Lhcuk3l5nqgwLZTMGhDp8+BXjyAvAD5otGlC
0x0EjWJ21x6Whr3Fl56JIhHN6a5krz0I/L+RnI4r/MnwFQhEDGVovHR4Wuh4zJrK
7o/2o974YXVzFKxUlAJk22pCIucq4ob4BMv3oNzwtW9LEDBmOr/s2l/id6GSEf3G
3Fd7Jy6Tq+5Uk4+hjY9+PDhXXMAdq+csGASNaHuvtFpOMhUeGbHiS5+7o9MMKT5r
PBKWBiapWs7VJxOcBn9IkDFr4eVt/okeBWXUpSvk4mHrmVAzLZ2+2O3dR26pjyhX
PTZHuCl3zmTdAsQvRe2H5tWjjht/8HfBnxFk7Z3KAbiMdyfHjsSm8vuLg2cKQdER
FtWmt71V3FNanS/3l1aTpkiS2q0UpyAOQOMyj7+Ipu+p1RHBMDBiR7iup9CYbgpM
fOSkbocBhslWaW8QjJS4CeyUA8GbKgj6UL1FFENNKcJpXbKcG6aE/kTRy8vwM8+m
OHrPtMTHkrYn4lfIIs/GVBeqMCn6Mrh+fi/3LguT/eP3/WeshLWwhCjdEdzTv0VA
H8ygYxLPnLK/1+SOOONge9vRt8ptiL18ZByPB+6pW4Tub2kfKfWbBdaZlzp+fzPh
eBJBjwQMjjpDduj0LB9UK0TNtbB0SyWyb4sNQ+84PWM6r5/U+QwBUa2oOVYI8R9m
18WQcwytksa3amg2/AZLcRLK+ncoKFMmuwGo9G/JZ5ibaUOY0sQ6WAvMRc3acVPM
7CU01LKN/kHWRKS00SkRV1JHiv0ZEl1DzRxZgGoguhgazmTJGnIhn8oj+FH5uqie
27O61mayo38Odhdf4zy5mwAY3QRu2Qj8brCJOge5jjov68kV/kcgFiZXQEhWX1Je
4No4cFfdxZdguypK6uW2Y8aRXG4toMQ/Tx4oh6BsI/+uVo2snzA00rjGDHmD+8r6
Rt97sCX+GQlaoJqNjeS0IMRouazcEudEV7TgH0SeogbAqkAEiG2FLVHYBpnqFeEy
d2byebqLP+hsauohqEdrKR+7LMYE6nfWd5zpaHyPHAzmRMATd54nw2uZMlpOboF6
3Tpcs1I4eTLBs6w53gHDsnLqijcL3ynJLYm04ExQ7wgo8l+v8jvbAMk6Ddc3f/rg
LATbHgbccXBCCQY52iRl8Msf+vLj9s/NkNt3EQwAtcHxxTuCtar86q6fQeYGqIpL
mD2cj/NCqcCuLzUTND3LtLTzsrr6hsHerBg+LtdA2rpI2K/G81GzDgh3CCoZqss9
Z+zNGwNQ+Vi3e8pAT9vyI0r/7Lxrs/TGIw3L6uKX8tdqx6Q+JCX15y1iiCliMlIm
h2PLOyAILlyATr5MdS7hoBZ9whaaD12Zjl9VRXZ4DdZ9oO4Jin7tW6N5Z1oHCmYz
QBTE6+t7vQelvPwt1xTnjEE7fvlspYzvUbFdN/VZ60EscgFqkUzLmknng35i31xa
ELqL7IZGasXpDzxR06UWopqw9rmbV5cKG0GPZbzT70jwpDBI85fqy9WbWNCRA15J
7WJZFSfaRYmLhYufrbz4bAPnwgb9FJ4XY4IYL74skUu0AqoeX+IvofMTAvum6GCi
t/x7EliHkaXDpUJhHo7SrwoWsh/DOfvRvea1cPwNK+y/l2hE6QqznLUwunUqk1uW
of3J7I/04hy/scPmcrVbjzXvYkPfj1GnMgkJc0HbNqMCsKVYoi7yuKqyklhLiuEy
TctCVxgoBfvEgUpErUjAlGWAJse98faSyszDvoRqhgg+vT5Lu7QCGjhqztSapwFR
gyS3UEk/PQcza1nLjhZMeInGTeVrLC8eqAW1ISi1ay0G8Z+J+1BGlVs6V527D+YR
jz4ztAomeW3NBsk7d7sIpUGX+tuyliPftu4xCOUkmUEbxBeCEuEv+difHbRrQnXH
UfZBTBKEUUdxVngVVjz2qnabnvDDopx3teA1Us+rXuKYYgLYjvvXnxkpvwy+Ft8l
dcCE5hxLxA7sdNiMorctu5mJfERD9yzg6PQIyH2Hdx/yxyXjBF1T04UDtjQBC7ok
bWBQ6w6Qs+Dn7hn5BPcFf5Dolx+BmOp8qhdf9gZmJxDo9HGUeE6DcVufHZLP9aWb
dFvQuuR0Nwu5Xmv1AeiHJ9W31IG01k2mGn7XA0uCaEp4wOLctYMN8AsEVI+xF31G
J53JLjDYYWyUCBdR6p/3jq8CQqe6/eGSapt5xZ1L2b83Pn2a/f1UMcUCZS9/YjV/
8zEDfOYV/uSLsNiT8mv74sslxVUGgtzcIpqgE08k0bx6mkbX6/TcfzpmLbkCqJgh
mlmZkqFOHdEyEPsHfkkVSxmfUtsP7VB7+ajrB+gu8Q9mL2MUVa6jjXnZ+zNfHBkN
9FK1V/2HdUBwtf9JynX0cDlXQPWIGuLfdD48hWxLRknImIVoDaV5IdsPpdyImp8q
lWp1aht3LP8SQn0Dg3QpO/fGB0akM064EkrdNH+nC7GOaLZxent8eFUaMGQOsTPL
RabQtT/DQN8iGqRHfZZ3a9sys60iq2qyTzIhoVZ1B0x7q3Ku8Vpj6X6fPPjgJtxe
5S5aABpyrUhqSqkrEgqOyvRH2EE/tYXo/YfhMqdPqgoZwvvsDkpZx+VboVQI1mqx
vdNgp5dqEDqY90s0yKrtblczh1cUFQ3emS22RakbgxFoq0lq9/E5Ige76oGX3YKt
3vic8IJyD4xWWfuP/QUK47q+AdB88D5ucmzf1k0s1NBZ/onBBO8lCMpY6ApHiqyg
HcLecRTelKV2Rgw7vHwBIowRig5E1A/9CtYbQtlmS+F6SH5+0xhisLI2kGOoGRRK
Ca5AE1DEyl53qT1vs0Ux4OmCqjo5uG8Nkhuwa5/PSkiSPx2W0pJVwNT2dOUAKLaI
jEbNindRHhYhJBuMtfrhQXfXjBSR3v0FTyDVoB5WCHSxGF6TLUWGyhoCPowb5Y6w
Xpuo2DeczncUdi+8J9p5gEjUDpaKkn/J4CoS2o2Akzr+MWnYOSHmD3nupzkGuMMT
iriBQ09xTF89CAOusOI102NYK8RSJP+a2kq0Uaczx7QNmPlgVAiYmSb7EckEZiPw
vrdf70OoNbaQ8IWw1kk/AwXuHZO3vHQDW+XIfI0CbEuhV+ZhEfjuJVBxbTqzjZEn
9uSoj46xpmYwZdcMLlNqE9jWh4QdaJxRCtWCiPwWsBuDR8n8eNa+zUhXo50YCfOk
0MWPy9DI8VqL8oVmP1SGD1vKlQ9LQ3GdxhiBupPR4MNO1YZvo/ybtKoERhE5+7Xs
Ew32uzW4DecqF29RMIdQgdqItrTn5/nR2jxdxUEaOBVQZOvjrkVTGz/rJMeSqn1P
VC8iI8J7yIbpPJVQdi1HwIZT1lTRvhszgXDY08S/cK4PCsplMIZC+Ssw/Qlwtfkz
sXwJjk5q3QnZMp2tdApmoZ128TEdrvs4XkBZcDUnZpIdAn9e2h4PS/19Z2HWTI0Q
+j1qO+TOGOmX8slOGnW/rw9jouebb3CfwblmgjEGbHL5jaSc4U0TjAhiXpDpbUxa
xNA2l6/7M7dOY7cTgaPLMwTzTa02rl2tIpheKclTPmjACOczOMVHQTMFBLNaZHLJ
BMkh5nn2clvTAbAZoZpKAQEKy8Wa8QAJecDTYJLI1uDGMlKf1La5JwQQfvmo/TIo
RS1WCEtUdK0HrGZuOGf9yHieyUQbNoXDNCRjdCS/aS6J/7A764ccBcNJpjXe4kic
R9l0Rgy/vdchOJisaeowlq96+WBKx9ldR2wDFPtDXL9KYmEZD9CrDH4/kpAUyG79
fFcLx3P//h5Tus9qm6U6Zz9hPWg28P6USCACDEi3abK/RK8+U1sxuls4KKS2f8oT
ju2pl5rEqJZCEOTQEiBaAIk4v5pTFLuxhobWcyXdW6+a7XF5w8Bp3gNLlGT+nazl
N+3R7tl9TwNhMg5/WzwUs847+Bqn8rI6iB52hznIqd3pxChrtvUFA0scRRfkmYF4
JqsB71jCfFSAhilk8j7dTxdDima8+X9LWeRpxJEnrfbVlFDI7hovSXAwqcuSwyy5
noUS1C/NbkORNK5ObJrgIFVncauFaWsYURZYfInTs94/NjIPtN/dV20KzvoLoPhe
U+Kze0kF2IdVQAGnKFwm1Q30nxVqRE0gtSjKJCgyd51aE0UwGUcFoIXiCtITlyaZ
AaZlgebkPE977+r1Tk6R3YihGWDmW/KeL8ZivIZBHwQ4r3QfE/F9By8Jo6jlpNjT
disVbvsiYRLj2P+lR0c/1ZTxtXvdrUWJhEZdl7WLqNyhLWmhoTV02IrfhtRdJfkI
rzNafAT0/QhvEbDm+UFRpo87p0G/ETjQ/j+5+WzhF+2mx78w7upvAKAheRglwQ11
ktebhLweMZ9ktoiIKJPUTUstQ+YD9/Ljs1uKZ1nN5eQ3JWO9k5rkqhEzwRWdWwUE
eJbssn/kSmEsjGU5FCIJ+u/oGZO0tV+RiC+T6SV/+d4xTeIA1i/2zniP2TFCgWSR
S7eGOgEDaCP0ThYS9fDN5C1M33iPfAyE/TCCjDUXPEumV1fMYqhEgU9BxbwKWIb8
lmbsMZYLBmnG0xAe7Zhlp10H9XA8xsKBk0MSJUPtQklcCcLMacPuouCjyVijiFed
vcy5ohrWrJDMpX5DPJ/8oM9SGJw/HgVj8cvfNUrBXZCTQLdAcEaM6OO++Q5ZrWTl
4Cq1FrG7apPy8pO9ePaW/mfeu+Z8XSS6M0paq6chSkUwdhBDTV+Aks8+v2F6QpjX
2fc+5s7cHVus26FhK+hkII7V8AjBH0Qo9XHDvyuyxI71xtdjiFRKeI6r5gTk8egZ
WJWDuh/0FI0qlKaGU0w79AZf9ragfkGCDzmWwAVdygisxJAFZqyLKanbH38/Ox5r
3UryFzAOlgBCB0ND1Wr4m6QvOA3fQlKEVDwzFuHHjy7gtd9oCTZEIvo8VRbILsEG
A0sJwrsi1KPkhaQwcgVxH2mYfzWTKBCDy4iVL+11LM2uV3U3wr+qyx3wMF8UzV5i
Wjg/eYQa0Zxh0jaZ3k6DYtWmoz++uWy8SJSlNA0eibplBbmmhg4d3Pku2+3+Y7T2
g/MSKfRJCHa+EvGf0SYma7XU2l8hfacfHqtO+CPOGHIyWmv0Tb8p6i1ekscD3Uwt
tAVdAHULQqA7m6WpSTbOEAeJorR4RfNApOt3jjobqQDCXywYLYmi7cO+XBnKgEi5
eOspIZo5sYeMiOZ9+yS7TyZOUQKf5TUulSKXBLQockDs58G0NjL8Zx4IobbJ3g9Q
aQWc4cNGHedPhDWQSW0f8lFEZxJ8KVTyzQXvMJbkbjSHlMw3k4VZdzXwneUsMOE+
PF8QYV9/YseNDbAn6dXwNthybjkhwKEaKSaOy50R2Rd/4xCZsD1i3I8/vAIgOKiS
6pij1QRj5/ObD1CKsFuFOefoX/ktJdOZihCF2Gk3M5wdxBXh4q/zwTH24q4votCV
dXURgatVj2aHSYq2Grk/DjzuyZeCC7Huiw/AHX+vCUwVVf4VslG65cQ9wlaY8QD1
FQnacZeftwzlmtgyqZHwnKbPlsLJ/HAAHUollNECj/1aUzprHp5MECehzamLr5+7
GwyaTEtxnWVuP7k1iPmzyL/kQzI1bTOSg3gep270EfepOTF/vChPsHhljr6ae9la
GP8CiKlnAe8Y1rCSCwVx54S6pD8tw7fNYu21K1WBQTrHzp/ejjMCGnpbKWGxEAd0
Y16XlkJxK8ysnm84b4HmUaVYSQ8ikIhW+I/0WpNy5v2220EOwKWqCQ4t48OXsaAl
42SvEDIR6ry7wQyvqrHnCXOjVjf2aA894Flbr4hfYPTCErhfudgZ1qG1ECmtV9Ax
Ej6yrPvs3uQTxXyj23Pg2eiT14LN/QWTDRGQmBXIQ/ko5lo392jAXRyO8KIvbmRt
x4XxqDnTJbLCuUF2Y3op2A+rLblbXRVUTgZgp/9vapYbv7+0gfdkjJ8oNqkSLBoB
Wt35++awpmliksgt3bJ9xsEQVAiYmMkDBDIvacghUBoBPLrqiAmy0CRFpqomE6s4
Faw68+teAH6yFoxu9eKt85P5ZtCQkMj8ETjvTM6OKAUuJlVFp62kh9HpK7GHv4SJ
ovoqPFR98kcW24CRdUaA5RK5z87KRrxTSgrMFNSOhc9XFLKFImSYGMadpHzq1p7/
Xm9jVP8VsY4QexhjQj6RY2lCRwhGH+aOIkcqtYMJJaZJ/PLNob85rVp91A2Vxjrq
h/gVLL6pPqUtayT5Fc3auRk79JlqXtxbKbrIQwxI6fkm4x5+8iFFi+Jl54w+rRkb
RiKdGzWX0dZKPL+GrIyn0OjOKA+dEso5ldOTvO+jUDoo6Mmnz001sFZ+pT7rUFRb
PgfXtL2HcIq257JEtksMeBDrFUWSoE0Q3n1JPYtQGNmt2kPFioHzRHavcx0tjgTC
XDpVyAVy6LanRz1NB2fuadD+Opp+RnoP3S15ztqX8hXmG+5v8A6kWMgsuedSPUaO
Xl+NAXGpIAyScVZuk75cY51CE6AQ9yCxkAPje3jBWZljE08+Ba1LiDNPPwdETXvj
n4JWtyXORRofg1c2wiAx/IDJ4klJnn2Da35EHhuBbX7YAIEnv1l/mgN5jJeW4iyh
hVE1evoNTSwVqjy1ZChyZc5y05xzpoC4wEePu8W+SSXB5aCTlya8Jlh0deAc9w/J
oyX3+FUxFzpYNJDT0ByUT2a0ATtKxokdMqCWdvu0rj1CVyjaAdGFiTnOTcos1Xqe
lW94rcPFKIUZt2n10sghbpeg6oi2rJEBecz+UBb8ZwDXwuoStb7CXHUQxEsGhNrB
XRQFQgIg9uocwWvqV9ob+9nkqkCmBlWtcYUVTnMXafYKJOXHNQr+zhB7ffXBOwfG
pHhmlGEPwxdIVUNGq5nmcCMa6JfFBabQPnxk4SHY6SB7C347XQLRG8fNz2kFqox+
UJOAH33D7J79KNAWDQDnEXR0o3bJ8taJZGdw0G7rXxpq65B7Id5I044fXJd11Js6
gpFTXiGfLzXfyznZJZ8GTF2vknOJTeWLuuBWgFa5oWtB6EJosm+489QILAFVDbKA
UbOKQQOpGwWDfKNQrmx2bKCfyap2CN5+/ZCq05L+owpWoesgIIMzXn3QM9H4GlJU
5R7fCe+O0r8wJva2h/wqS1r5pQybzesPKrB/GhMoEJaZSHoZvIH8Hx05dHr5DAKD
Vp9pEjJJixvkk2DdAqzavkKbsLYj+pRED422VIBDElYERais9rQKWuWVKv5q6KBA
EYXT40BZonGppjuWk2CKbY2VpUJqrvsW2Q0qyGPL5HZlDUN4OxjjGkLGh9K/vxcN
iI4wZ3x+moPk/cvs6kr9n71Sxg30lxY0j5s96VHzmA34fMudnSqY916bwhaY2jzY
8y8EXAtyFK+CA1uvuSFhedlOOgtUFGZuZNoFiymAc/NVg+wc2rfmzBldWHUCw/fw
7KHJcby5FHsdm+4TDGfk7onEvLZAMQhHhxXt9m+tdqHHC3o7aTGmEtK4OGHP6bKz
SDCdy/CMIVSH1+XS3ayQ5+VT8l3C0sYuHZrZ+koCn/YgNCqobDn2HhyiifBSgj/e
YMZM7pDE5wmcb5gA5D9OItTHY6Lv3CVj1BjE9x4NQwsCAP0tuMr2xam82XxxIrpn
LRztjkeRqR9/DFy04Z4QHQ4faNJ+geKYbUT1ADXzR7VvuDgcXNMv+h5hTQkCRUfc
dIiT7WrKxxWlJ+j0yFs2nJ7XmDEU3A84QnXvlyDdD7LWN+3Yt1d3krXJD8Aq3lLl
6Z8VAumHqDRwILqFKH95lgUTIgguXdKRWLioLky8k7NHQX/dPkhhFktGZnq/V+0F
GyfiSv3rLjxqV3E2HXGYbbLNtuAUBna7RILozHYzmDBYnIlcbiJmvuGK/Rhgc1hV
SaQZ+qyEFqDzBvFtfdSJQiHGm1PN0h1QXJfItXHcGhH1O6QHkJeQYiEu8yyRxkJ5
ms5SHTZeelp59hJ3KTB8fg9PtqCHgo3eEWw0nulSHAxzqX7gPPNzP66+Hx/ZIdK+
3L34VjkGprs8iq9sHKrTmSGzeyyOweyQOZ5Ei7AyDa2sgyEYQXZalym7pWwWNeyg
dT8j+n1yNg5W4jMTQnCYE5vRQGWmLHdcUltlbAYb7U+ibfWmtN4Fs0jmxmrDQ6hq
r3yac/uS0D6VJmtJdT2+js2bLqxm7vRCsrdEWNha4RduNte5/ZHNiJpFk8Vd0z2W
ctWTBQ1Pq0mPl1OJf56s6LOAFKU24UQw0fEH+YwawXESzMfnM0Jz397b6Vvi0a6m
O5VLTSuMsxTWPWOKgKI/Xas5BA1nu8XMEARIDK82mfAPDmqi9+jVIWDinJH7YAzl
FYUZsynZgyfBvSfTnU3qFnNOn9ONqn2q9FequAeTUcA1+41kNP/hUUhKMQwDSG8B
7BCjBb/ypFUB7HkQ2kvu+2GRN6NPoLx3zmaJbLk+Tx5+bKqIziZxfFx86sNqFmv/
KgWL9yO/35w8QEkkogzccZj20IiFsMtCAUN7B0tKOfnnOJko2Pmuid06HL8Mycym
vxwmuEPnFPynZvuotlVF5D71slgm2Azd0m4PJpYgz0MVyAbEN7Pj/e3T2hMbVGF/
FSxpQ19AeNEwAlfGFtEWxUJl11lP7Xz8Er/sNNy4d1cZLY3xJjcWk6tUCvyPXtZ/
h6GBEB/+s9kZEKlRawbVUnPCBeJ83aSrBJE09tTsJ4Jn7sEnTnqee8CGTK8mtFQV
PS1t80iuwTHrqXgPRS/ydkNE94wjvZk7SPLEhVEncxsfhZ68O+OarnjyR/2bmVwj
VpLAzzpWcQgRR5o+bshptr0oPYLssX2Cx7Ah6RHwO+CRx8tM+L/oQJ8q7D0BZNg2
xJWF/Z2zuyLEEVZ1byW8VRFBtosAdOXVt1+sLdsA18mBi30RaBWYprf3CUeZJtbr
rOlIndj5AtEsIaP9XFhYee+UDj+2r+dja1BIFJZfaNN2adVOtI7mXs5W/GbSEJtU
yCXLCUP8acRbCh1m85de6HfKWkucUS50mceyfhrxyzcSixa9FbXhcLAq4G1YNIB3
hSoB5aND+h9wFd2+WxJvW1Ow53Sid2rNq0oSJfM2yfhLnC0hsGqc5lSVG/CWACIB
WMQIEMkx21pOKPoE65uE21JASwWtvrxtQNNQ+rZb/FfdE64YYV04C2KVuhLlwg3I
gLl8kLqdmeZZZQhvBrFA7B7bP4nIcfIEdWqB8L/+qy9N8biYfArdMus3IpOAWX8l
gazchJzIWqMfZ/odRlZot0loolthfLV4FPIznVYmCjCu1//YRPsQgFHgY6pcDQA3
knNjTO713nfI4+QbdHIlDsHyqs5K0b7sDnrD2yx2o4dHB4F5pIK8hX7OZG2MhLd9
sC4IBy2H87ty8UEqeMccSf23KQnkAixQmxB/oRs2c0G5nLsDuDHwjLl/Lxpg6u58
XiN5koC3Q/VGloq35LBdE4CHxP+daU86Nk/eJF60MAH1njjfwEE9s11ypDwc0hfQ
kOMKsAxnzvqUkv+gmJ1X15hMNnBhfD6VUrKPu5CU2JtIMDySyOMNc2ZZVG+PHZtK
Kkhcb9bFoHu5ZzpQGY2Uky1mmpZFef3PlSyUUyPNoNaXG0y8RLH6NkvCBQbcKK4N
R01uHu1CXxMOhseZeh/HadhyofLbR9EKoNvKokJnm0oXAlHaAJmAixC5AIJLLV7n
/oAXk0Rfos9gxPKf03ivB51CWanN30lFJ4l+eHZKvY4YZo0ZBnEP6NmQtcmJFADT
R/giwTCxjgltbde0RNgVOBOkqbAXPZ43IPxhIl2nikqFgSzUzjS+2Y1vSFpJiXAk
/8g7r+Qm+TQUFxZa6ooycEX7mZEJX5IYBHGBvQxC0lonqGqlTDDXZO3crgPrIonp
Mfi1St9YM38fj+U7Ba0twy9DWquvUJ9glejHw9gXn0L0vUkKJO1lBGI037FUcHF6
jRiJw6lsQkfP4sTGVvrWZuVr5s+OJNrZLC42CgJtxuluibi1usv+00rzY3ddCW4W
D5Ncq0sC8aoWDItTuBlGrsP9hzt+6NcjEAb1TQa0ZSNuvI7D/ycILazqqzHtCPMD
KhdDjAt3RtYSihWyZvHn8HEylikeYCA2+mOsrSNnK/BIhi7AOQXhesgTUOs5IOaK
AWrSVoH/vcu7PTOi5pWLHAUwhfwHbR4bYqA6UsL7dhs7+cm52tQOyh0I1HUdnhfK
rQgn9WujJHW9qAOTF83Njk6JAJEvWqu7ELSBg/72D65Lfp1Wxm1Px9bkC+KXNFFW
bgo8O1AQYGx0wV3DRu/CQxhPEtX6g+3MZiSWKzmlFg1hubac3zmEAJEo1KIdjLs0
5o3F68ZCtb+YMpFOO8/tMIGaAMPmFj6jILVGiqcHT8gbo0vDq23xCql35H3uC6zp
PmnleDbMh58ub7aSwUj/ajvUiVrVScC3zIclHmslycBC+9D80+zK4188jGFuFa5D
zHRel+wMotePobSOuaIGrt7AzSVU5rLxgxYjOZOiw/osxFndMTVjiPKQzNXv0Uld
w0EJMA2T8Gfoptx2kOGCEHO6/2gt7d08hmzIUfmUDuwwHf+PSDegNhhMjKKOTn9i
b0r1dxKwu/OrDdgSeKMyYUUFiaM2WZHKgkbaUVkbX7013y6GfYRGkJyVSBbynahV
eZWzIbtTLzXLE2l9Xs1LL5Y/hN1pTwRP3PmHc92qyLJP06TP+CVvxPUwkqdG6ikS
6Po4DnyZkUrJRwA53DEEC1K7w/d7ywxeSxmYBC3Xxa8PTy+OyV7o11QZ0Nt87Tuc
MltowPd28HZ6GAHwVv9tRiUiHPMZlI0BHj/loxqLrJI2eRWqIji2Nrp4A7XSARDl
LcD1jhmk8wp3sV/wCa/+PrapvLXcqDXHjkhtc+SrJMz0+X6tpZNzoGcQ4K6k5SOn
LKVk4iZvnDpaff+/Y7XD9faZqmKmelaqxR33Wjg07gonX5caeZzOuRR2btj+dwO0
9GZgMXkDk0U0hacxIkBO/QpDsNXCPfoydQCP2SSwqCBVf3sor4dxXFnXDWQFvXZS
vTaz38H9p1tBy7i2ngJJymH6w4ooNJzo87CFdjNfVpsP1sXmT7QXJvoWnS9DDu/M
ybZ+BlpRwtKXgnAIz7Wl4Pqp65S6QatME0Qs95Vedk5mXVPNQoAXIpB7cVYEIBn+
ye1Fsvx0vknd3yBYmjQcX6JPxPRaxPHUubpun6fdZQxYpGDtta/TKB6FUbhaXame
g2f60X9LvrjaQM53DYdcj2fgm8s6rCfktGodMZUtHDQMsiirw/cmdhT0vZmvPCBp
`pragma protect end_protected
