// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:45:22 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hA0X8hJPZnGRrjTFPvNDh40I57t4oThJAzP+iFsZ42WKgB/kNgU2ARSQJ0HJHrK9
g0IsTs90NF2coALTU1GZVmuIBSAcblMW0+1cAMvxmYdv7pvow+T7XVCsUDtCWYM/
Nd1iU3x7m2r4p8071AQPKbqjcn5uK9YRcPEMw5y/Uzs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28384)
OBuYd8BC039TBV/gADnqG9MXDa2DB03XVDMywGSrHQYDeNVKm9+H6HNQiY25jqy8
yaj3IiQLKAp7nykj56enKFqeFXXwGfaZkkrZGi87L4gMqpeEcRSWf9ZrEgJ7DrbB
QtM2EiVp7+IvfYGsPxyGDGx725qtnw6WR0gJ2Nop9wnn0wbV6XfvIaWSZLlrZ0vq
aLsBfx24SCqsQcAaSf17lDfOR2+JX68OswumINMGyclWYo0/50XWGSEr2jCyViqt
viJ5uHClIYBHkmLOMqPUuhD/EHF2aaM6atlz+azGnmYmNkNz6HkA+RbG99OGibxn
buYge0YaeuK6Zqq4p0LDo2ZSYrTcGeSFpTCLG3i7s8CDPHHt7XYnYQY1t3Nxz8EJ
GO7Mpu50FwKfXUtorwzb68ySP2pWv5bVU6+1upJbefOReEHVBMoxtC4vShKUjAji
bxJsE5Fi0R++ev3aG0zCM/Q9M1fjeTf2/EH+MaY5+k9YH5OyChYx+MLC5syEV3kl
d222TMubTu4mr+ooFEIyxVjam5hivRi+gYQD+2oHMyPFBTAWfdL7xvtkiVM9FHS0
3yDBnBKXJUkqTdNAswk0lKsV41EmieqVtb9nSkhp5K8542yrG4LBeT37A15BNS98
AWLfRZ71pou/BCvKZngSXI8QK8VaSowZjVCB0JTStnWMYBraBksrN0LgWnDjOnTz
6+VPV6bExixJ3rWphJYe9euPSi61owlbplY9EM4Ci68h5MhItO72Ouuxzld3Ua1g
ZNEF8orgFiMzPL/BsgyDVTqlq8uC9rj6uBjm2AEhLsRdKnO8nO7EQ5THNiRXQcpM
aW8IDdQd2DxwE7198guBWlSO4rIkCydiWJIR8nmd0P5hZcvaL17NwmIul9U/HuXO
4q7mEk/nXjzMATnBFE5RPj6Ymsd5dSDOmIgWUK54M5RYQpejc74cCaGjyN+F+kto
esBS96tpGIIuCwXU7GfmkFwTtt+4gEMbfaIxxMWuidItCdpD3pOmakij0CCWQjWE
X4DIMsMSRg8v2NZymkw5KwPMbAecXEGXwr/5mcX2xJ1CJYRX4eb6BYhDfU4vcop7
iSOwv20C2yX69fM/e1ie9/tqrnERNuiA3CNJZsaiL9nRoWjFBfbiBhcvRsPLtiZv
NG37YPLm88c7paYVnmeQOTXqc/iN6AEC2axDEJWzic3/Uesci8Sw7xYaUPP+HUq1
v+mWiXAXX4FpkXj90yX1MG6C8ngQF9abrA04x0Zbtsw+Iott/RkivVUB1cOgNyWF
5/aGFSQQzLJoTCWXGW3Zs3thJlIr1Mt9iWgEdE97AQeFG/rJEuGxsRoYPa/nm6pZ
e3HHQcN3lJijN4CfGx1lCR2p836+cIw9M2xVJTdHe+nhQJ7yx/uYlYGeDRaijsKa
uOEj1a5h/L/YbkFYjwyI6inoqd5LXhjvoo0lIK0V/gGv8t4STNY6dBn2C9lNVeTN
Yw2WnzBL8oBKO3IwyKJnbMmON1/FpVCUTdrFaSvQHBZeE1E1NnMqImQ5DhwH0Gi0
1goTNv85EMbJd0+gy4G46ScNssvuyKKTqVAc2GkQkkuLNOPxPU/NS0dw2Pp/a3de
YluH19a2E9vSi031VDET/u7k+GCOEzkF4gWSVGe6u3DR0RcuO0D2wK0C6G4bZsyl
1jQX28ykbVIIrdZ4hbt9pph8lSO6swZFtAl74EgHejtKUWf0XU0+AmgPJfZ9AmhS
ozvyssqnUsJQ7gBOa7m/pNt5OAS1Oop2I0KI6LIRZs4t3pVA1JWQbp/P/+rZHx9z
RvquP/Czk3Dqfzmt8yKhJK9ESyfgRFqwtQVmrneukctSxk750CN5gE4WE1MCzzYC
T6OaGqoyprQZwuhr8Z8+B7/G+ZQcI9j0mc4hQvzZW+rmv5x+b+M3soRIlmvdqzIU
6qzgWVRIzZW2A2C+M9BDaKECxnbeZ0B5KtiEQjcZDDW5kXgG/fFOhe1xJPzphoV8
P4PiemCOrfihvwy/sznvp3teNE9QzNL64ZTi5emIiyVoQlb/36TR940F+kyBBB6S
bt7/ogOEzljnx1aIhT0Dxl4eCYVOD8tfN5LSWwjr0ZpL9+kRv4vmdTxKDiKMnoJx
gZL+7Uw4vKyDrKu7mefQt0KipFRFOtYW37FSwHB8d1jwlTmza0nJvqTtKAaQv924
Inymg7+na3IdM+tfQDK4DF2f1Qs8LctF/mSFcPzepE10pxoL72oeC6sa9/qh4bWx
Cydp5Vn8VStuwXrBc6Bm4e+xLcRU3fDSNZzBnsTT4lxj1DIYrK7W+vtPxyXu8VLs
rFIPieUugsls0onfMThUOVv5W8EQmNLLDfrdAVY7zfqcDMwrcsD4iCwalSDjga+u
jSJtJXCZjZhZuVMJPhPizSbdqGodOn+6thzK5jMc+mwruuPTZwrR9/asGArtpOvH
3y9MRmTExMXXLovrtj0RLFaCHylVao0ellzd5f5QrGRe+h9YXkEcXEmbhvjL4U0x
c1Tog8cCOuB+08inxSfdTmb3L4Hh9+kPCqMnRQdlDv5RVbX4USuUPQETjOxCwRcP
Og/k09cdzuhxwPd5F1w11PciF+McKh0xHW4FD4FnfJ40c5l8G6wE7yILvIqeJV17
MLAUVOqhhLpxOkU6Qqx0WVyQjWX0V0O2HTKE3q/JCWAVt268LkwIzYS0YjBl8/dN
iCU6hHuSOLR6Y0paCt1gjy9UFjSv2SzCJO4aab55VvR5QWB7kZMR94K+2T05CD7m
a89RdQrc7q5C/ubf6oMwdA+rNgzgy+aDMjsnXKcruEkJLPnjUkMW++TC656jq/CX
SZGfnqAOoKtTsh064aWRMhl+PgFlnDieQAsiDY3fDvLyhJpI0F0wWBsWvSZSogiq
qgmjRqbFvT+kHuTZ2JSqNzPsadHv1DV3ThxpL0WbBU5He6Yveixq7qUvEcUTRFjI
UJU5FpZwpPftiOvqo7No5MMTsn/SEufwd9b1hfD2g7W193AMq/KfynF5FH3k9gkW
aF9hFy0aktmhLCvU/cgHelAp9tpuo2lMFjGTqySofHdRJfEzGki+3141uFXbPGjD
wZm67hnv2bLT0y0ksKkCSe8hmpog+EOmztpxEPuS2eVZNCeMYH2mkWCFD6QWyiig
mu9mVSuNkWmQbCD9FvGwE2ncUcPTsBsA8ZFYk2CX7Pz7oNNqttXIFTEhcOkQFR1x
jzJv83BWIQhdUDWTEssaqSKrOPXBcVfk5JMCtEun4ZxCcHlMLorNnhKmnQCVe1An
mrGB9Q+zEADyHAaQ1VYp1wj+9WGQd/a2cF9Wi+I69JYXwkRI5unMNS6lDMJNNawW
sCHFS56bm7huZAfQaRmdFT1+mf4sSx+kJkFKbAUDrC3X1fkubZcO+d3TbW89kq5N
reM8ZsZ0rgsqLwvBk6feRdhwVQX7GyanUHYAGNf3OrxmP0sHBJ++i3HhxUSTV9dw
PWDHWfk4twHUJIg0PTLyQRs1NZzDx5jxNrkVjGmxW7JmXYpXWvQAcaacdPhIgxh2
kM5JS/vcrbOISaHgO671Fpv2tifFmMtN6WnDvYrKQsmFfe56OAEW6IFKbWdyd9Ut
xNMiHctHVK1uS8SGqpLtkae3+xlWXoC6ekX+OysYjX6nbNKD/7bvEWVVLxvr7dqv
3vN6qebcvZhevmefjSWtf+95Q2rgwdlYHNY3n72ucbhRBps0mrEGAwcL/qsQ1Mms
LCTWdXy/b4F6N/hg7WcIHciqilZ2VP3o5F4WYQgPIeALGj9PKUDQ2NcBmod0OwCt
hVM8S0Z3Iy8IKcdxGOaSjz8lEZiVsEbo8EdwyZ3BKWqIub4QqpKqFTwgt8WrKc+R
rkOLlGDBgUu/dq9iLUCxirhvGlqiQa7ESoYXK5j1tzDOIP/PZN0Im3aWpYzBt6xK
KpuT/DApWOkE5WIyIKLVPUUmis7S9I271d2MJu4Ie6D71p/Zq1gVdKFjHcMcz3YO
Bredqd0QNDvynbaWv8xTxB13HydsJE0oc1sT14rDb2FygEHELqDlADTQjaHEek/r
puIaVhAi7DxLCwkFj3vQM+wRPrrPuNLvr/MkoB/wiW40TWY0QRwjexbX7bYYy9Bz
OPl2RqUYe30vCrG2+2j45SIzLNvl7GgblO+FYJvIXrau+FgWwoHCtzzP0E0N21Jc
c8Gz2tGrT43qfaM7RtCM4/OIM7Yu/RCOqBTktsBCVxgvp2PzqR7ffjh+qljvrEzl
TvLb3CjFNKaDKGDZhHMfDuA+5WDo8QR6qBjfmVd0hxdfzLSKFmjzUzpqqb7CMiAL
gAMwKyvZuxFP82vgauF54HuCFXQEiMMl+pc6ePbHDWMwVtXyXxw/VIKaLdFigAmb
CeRHNZzPHtskosmjvyJQxafQQ0v9o7Gp92d5v3bHE25voJs6pscDeeTWtjrrOwun
cCe0+f1/SUGAGcuf3JYuya7fAVOfyX78EISZsg5Q0AhDmNs/dsC6PFUNv5Y6kKlU
6GZD4wGmK/cgAa5af3e78aNCgIwOMFvu6so2x5mTA7PXUocr3yj54LPvZiJ3CHfS
KU/PTdyJusiESqM3vf8oTThYnLPAAHYR0XlqOfR936b7I9gQ55inxogfpsmSVleU
endGL01MDdVmn0R8+Xgn0oPKWpN6jN2mwYAr/IOSEjivxcjqmZJhoXepAkvDJUtb
Lc4JgK2LJHNRb3lE9U5KnvdxNPvGe8xhPEIhC/oyYqDT70i2yxMkttxsJIPx71ud
IoH1v6WFxboHO33+K1fWsmRjvsKJSmR/gSOxmVDXvOsiZdaOgz/Y7ymjwv32uf9q
BSk2ZjimdsGvU33N7QviWh6dPRVQN0a+9haob+8D1eB73x/ocmQ97QEXLGc2F0ES
C1HZbswFyliX31bVNKmHPKCoViLEt2RHW2dq1RtuEC7RNe71Rij7KY4l2KymoxOg
bVr4XPZ9fYZa2jzgFWC4CMFQTczahf+l9QrIEDpWWFI69aChEmFPIq2eNyKobMEU
4z2MXCP1AkMfg4G8M5toxYKxEuvXESA4kIUxq6gYolMhBWQDWhyFRyYk54bUhPJm
LJmJKmvvWiOdojexsw6+6Wv18Y8G0I/vWl1x6n/66zOaVAzkRXn2M2xx43z9cLYD
D75LL4S/XQHPQWHUKgcAw/ZPBG5A7ECH2IIlle2qlnk/vtA0gBv14rI5+GzC6l+Y
T8BB8K2L+ZSBim/7r2U3TVbo+7OgB7MiMTqRvEv1Ti0XG5oTGf5ugworI5CFxaK7
/vibK01aSEpORTSSbE09sWxQTSVDq2S2MeYmBR+1GiOKpvmuHzSMSiMBN2e1DBR3
A3AJlp3vvW9WNEKnfxVmFckP3rjcPQid5Mu6+aMt1dpEZcXS6XJ9DvEGo6CldiyL
PULSs3rAbgzJ1/195Jc3lZyasFa932Mw+yw/qMbvDIUpGdOPGR3xTvDMRi8yKlud
OYUQfKneXcpO13Z/Y5sWAa/mXC/Zp6LKoB/CFhXLsVyIVxMvqZxWyPFDmZHlfD0G
WIyr2+2EWPllMlIKJxZx5W5cEFKgEp0p9Gn7POKYww4oNTBx/ru0Pob8DVXZvXqv
EBmoocQnUGZ9OeXlqlHNROg3yAcJaKQtGj93KbEEU22njfCqqTKOJYoctjNIlOEr
uH/+1jjVdl5LojzITFKquTjYyIhrN9TqvuYjGcvJXn2ZxkG8v1mBExLtDpwtJJgS
L1JCQYoy/2FVglTwjto+/KZcqosWt6EIXNZ50AYdAnZ5nWosRxYBRaJ8Yul19tNu
rBvSjwfQgK8saarLQHv4rUDpacgCHniruvOELJvvUNzd1g4EQH5jCuOh5T5EFo5K
4dFWPr5dGEXsnvDkdtrnXYWXKPI/ldEqIQo0K2iYphEwuvxDUrmub+Ru58dLnQzY
cRF2Bv6YNI/IneUkpYjkZU3et8hF4LN49dAwfwqwexZBp/hFqcbdlf7IBQSViAK0
5eRYEBcPbyJunVKEaNn0JISoUrXl7rZWYhOQmZyfvBrXw2u9YizGRfst4FbFUJYk
arE6S9ycvYuAqoVKn1S1ZUX6WTSvqvPRR5ke/HNfoqHR0PUhWxc1it2M/VMtRV6v
qJEflV5k7VTqwShlpfF2DBJcOSAL4uZAfFoTfeXZTlwJvCDxZbfRjAmsmKnthdvB
PTt8DYCUQmB/Wue55NO7Khlcdl58mxpV4vB56U6k5kMGv4k/qyprl2DP/4SB/wuN
D1b+thDW0ZlI3S7MXG5Ita2FSgkPuHDg1LFPdPvBdZKrGQx+PA899VyOCkqGGqTv
QfeMXGgCN3x2UJvGwmeC1c7BAuSWgOqUeuYDd7h98IQ6knvfzIcb+7rc7NFf4qDf
ID/UkCTbTWI8+pskGg49Df54KPtiKTG8a7KniCEOwhM+0vZcwcH+8b9VMgrjTgaD
Q3eacCWLjyOFm1vwy07Ch48/INoJSc1rVhag1eid9tZPXbf6UD2CtU0+pOOKdXn0
VT1ztyIhjSXkFVaIFWQKZ1UcEfh5l8tvudD0UOetr6nkQCdcHb4NqXTF0eEKPFFp
VeoU6WhViB6j3OYNShq15GkynB6l6+Ur5wUplxRZqHUYC/0TI4QMwe286Edrm3c9
WL8lEGVcYJ3EhW6Y3sg3gSPz31sdSnw0dTkgjIdRhqTxqr/IYWVfAYHpzucUbahe
alyTVKtKQKEiyuGCyo9LewNUYi94a2t22tR4l7fvZH9/XQao9Aubm+kHL2LZDDAO
06nqNLrE5zRckT6Z9lVpbl3D7URnr3lMVCpLMiBVl0/mq9pDTCKNa1aeQy6t5+Km
l7FVtckbqONPY5ufXWjdtK7Vq/DUDlVoSsNUSwyOf47spmYmB2aPq82Jz8qYUR8q
onmjt5ctgjsS+nA+sgCh6JPIkmr9RbKSLlrwYISa7zmZKgU46PYG2l6nFuToWEtL
XPPWDFXePo62tQdIpwu9QWlfQJ0poB3q6i6i/LF3StKuqVRkXeCGAWiyMoXT0nN8
+4o1+YTBs3ktZ+dTWhMepe++9LGQV2QazyHcyZ0PTX7Qpju1/c0Ri5lsMEEcn+C9
CAiRcoV5KBPPGYPhGc7lvc0MAzt1fzKF7WS8K3psywNPWFOxjk4Ci4EtzeNBHKKP
6ISZLa6FHFBcIlVh1AX7MRTYjL7edMs7WqC9JC/xyb+pOFzamwkPPXOs6wqUVBoq
6huPj0zTlj3aaINcFSsLsJhiAfP6fz5aruvTIsiw6Pn3BxtYJtnhYjs+AZ2Dd3pq
ZsR98j1m/i/AH+Th+2TPpJ3mBAvB7CIePtYr5MBXOgZNIHCMP3V6LUeXfz6LowjT
Ocx9En4VCj/PnEqQKDH0Zuq0HfRpw8pGBKv6RbbXOAHZb3nsgFrMUhorbXtryRea
A0uH48s43bmliCEpq1O6Ybk6vajruGUIy6eodMHNZF616gai6uMzown1+y3VPv8e
DIsdZ3LZtrSixqTloBbub7alU31LfgYf/pwpcMaOFNNA71+uNLR1NhKJvIpWoI8Q
ezQVuHTlcbDAQDR4/gEwPALfnZIKAVU27IGON7FtOP7gtp26YTPrj6/IgDa1EtLy
7eUylfnj73B0Fia84PpyErrERYgO1WkNdcOREvZw+Ia4m+59wKyYupJR9now91of
LFttqHPiRTy6JE2TP6EkR2IEYOEvMNVsgAumZ6miB2XVhTSroGhmB7o1l7+bumIa
BTaV2vIU4SC4cJOWw8a/Gmc3ntdpc1WWQWMqc/VzLW30OaAI6FM/feCtCisjuDLx
9GF5YIrq+BtA/Plv4lhao8I0fRdwBzZz6052i2c1H1T7dZep5Q6aPLSJ1w5X33CM
X7UzoP9eT2sx72ZMuIRKWUJSr/h8urJSL22W1EH3Yg5f3jW2Wxb8LrrywI4hyGbn
ve2KCk0JrMBFxuoY8vGSxqxLI0gGGMGEKjawZAiwWswwnLa/0SygHauRrGN1XstS
PLIfp9ooMbUVIaNLEjc1eFdVeK/+5PFhVzrZwNHtgHpovNTdVUXSbUTkz2KERrbF
dcTkMKE+5dw8RIdD9Csn038kMPWjfUGwxqwvd3emalqgII2QAjBhXlzjr36LDRXK
ctrnqT3UNFPpHb53IZ9D/zoWdHp4ZGHiv4+bttm/NzpO4hwmD2qrCYSfehH973De
VWN4zp4zf5b7XYlZqTANIWr9kmwyxxbLqDSxByH+8w3kZYh1QCBC6IRAZa9+Eqcb
VwfveV06MsU+8dbJOKbIR7n/MjkRCl4akueklCQOLZHlfQ+0Syi3veE/nCCTrf7k
3wYl2M7zgccBEIss7SAPflRkQWmhCAiUIpOmdf3aNr7hPvTa1rQzKSBI3/AdupFM
Sa4lj/5WqpaCxwywc7Wp5KufNBpLQCM0vk1D9gbHwXtPxhgXNlcQnPDTcaPUw9lW
6hIH+t47F5gJ59qqKa/b7D+KnkJSRYso38g+yK33bmYq5C/YJDbH94f2Tx6RzOM+
WNCqfl8u+t3DHqMSXgUP8F6T+8HxAc+mix5If7jlhhfJBZ0wM7f5cDWQXS4DDLdR
LB+aAUDsKRwD4o/WUNVT6gUIw7EoF8NmZ8ZRrws//+8UJl28+xELStpWZOW7JbFQ
BJwedWhoD6NC1Mpwf7716faq2wuKUKKlGUrtPflseV9+94gfl4HEfRhlncvr/zxF
X3GNsxdb9XNUIddS3cmhxZ91hmh3PJPkeGDHhDUImlSwC/3PY0/3+SF5iiyHMjpU
l7B9zo2KcskaqnmhVK9jq+d8rcOccyJBAop3xxP0QC/2EYvyXTKKrXzMia9oXSlx
zhv93UBQh0spNFA2+3UVMS/XhDc/7olVqmNAgT1GkDX3j/kWr80tGnZh/7IrGtMy
PbF7BfX1W5SYrZpJGsL57k3HRWqHV5dBsnBJMNl5so9PRSMX1QZ+ovCz08anT8jv
kzFR253SrVvmgbPDT/lYJBWBK67SEDdjFR8fztLY44Iz/PQ3NO2NhECpWxoH+bdA
2M7Vewb6F7aKVpbbQNEykam37zn9AjR6qgtky7vciZIQ6Gn96txqWBhYGdu+03Ws
bMH6b89BgS3VIVilUbE8RvVdTVxKvsI08lkY5BL7Rl1/qR6i1NpBAUjJAjUW5Ski
nBtqJUgtenZXbEDqJ6nF8yKarWYogvOnil7gvUcbknWIc1b1RT8VGh1pRrMBN6sm
4P4dg/Ay68+B4qUPHIMwdDfrc0m7c6U9PtF3m01D46On39XgkDv7z47hd3Rca5S7
2+VmJ/KBgdiU0yBtcn0/T1s7Z736z42rpnWrbp2JWdc8g0ckFuhMk11vA3eQEP2F
B7ORDlX8tJ48xF45qGsYHr0AsVelEU3QeHDvEtFU3jgV5Nkc/NgN6Q/HpgSV/czY
WCpB4dZqhNMFLLCjPZUqH6UyYKxw1wQJ/Zt2RQXIb/w3k/yfxY6kvkEBAk4o9UM+
eC5VWbN9B3PXUuBrfNd+cmNdINtIC8oobT5Wc0r60JhGrKaUKcTgLub7FGitgdPW
/+9GyvsfNeY4PCnovMwwi1XO27oG5E90XAUYaj2/9BUk1sGqi6mjmxfP6aTcAuR/
XTtaOI2mGH+liN8LSpvCbo18ZLd1uFvlkbLyRU9NBSZ2aNbeidrSwhEQvrihW9hf
0f9LYD6Cc8tL6g+AFtslbFk6MQwdnFKoVXYTlD4m5s86RJMeM2/e6ZsosojD65K9
et0KssIW91s444DMBrAYQkEJndXNJb3GjKAE64Dh/ABmLkycVnVD3s7NL0aB7gID
2GjlVCm5hl660eEFtdflwuK+hwbZuQQeF/GV1zM+n+3VS5bHD4WK2ZfB6VZWr1mK
K1ZgSX+KH//rx/kWtnmz2LDjciP0Sx0C+lLkdtztv9fRc41olMsz0sLRW6y2uQ8s
SRCGDP3nF/W3LgHIjUMntq1e6EqAmx7T4Ec0qnV+LpLYd9PlMFzoWPca144bjzyE
72KwV2RhX4L6MGLcg2BrG2AYQJTGWw/aLg+ix0S5IoJT6aBgFmeigm6Mad+x5Gxf
/AL1ahycQVaXbQFF6r8mgEEa+ysKKaz4zT1iKzgynufOZWd4HJhrScdiCEsvL7cQ
1BVVE2ZGtFPXivGnr0zysJv9CTu+I3v+04XDCJ5RhH+0RHCFjwr1VeAoc2604GTn
f3mu5AiqrFAFxCKLB4o6NAtJqFAPkzT0cAqULkGbYW/lt3iO7jiPqOmv6mgS6Wvi
qTaHCjFlWFPvOznSOGQfeK2Gvr50hAASpMWd2jNFWCXkc0xBykwnDgoDJGTp0SvF
8pOMGgTbX8wNCLl60HKSDMqeYrPGw8CZOKfDNaEsLRNSh2nteNNUtjE7f+vVoaS+
usADJ50jLIW2D8073T7E9L5f7biDg6YYwUAjxakEe+IrKBBu5jWKztsYuRQKJCbM
68nFXvgPBu+NNMy7Ci1xPro9AO7SUa0p/7tmWgxqKKxYq61tPcYjVxlAStZoy9R5
E8ayLeyy2j74QbEYVaj92GfwFwhgof5dNUxcRlhxySYmBkJ4BhTUnZJTyV+sPxAH
JxU6DHnOW6HKuvuai1kIhIiN3yory8Ms7XoQY/QumCsf5bRRNNYgMXbA3UvgZ1pI
f7fhkLWOrEKCckMXX7nG9RGd4zwkzfGgW8XmJdKwpIzNDN3TDTyh14IMLKYh2qvH
9yfJFKO9HZc9jrQYx9n3nwi60vHoaWEtg0oKJCBwGWEyXJZY57j0CA31EK7ODZME
M3h8ycMOZWLQc3kBivfoACaBap9ZEE9uySoN01i+Frk2g5SkmmfraCYsj/9otPJQ
sXYVOz226soPSgiTMJUt9YUhrn6u8UZgOhRW8iC4+kLa79nrp1wta+65951a2c7c
5L3nbSwaPofeq7+nj9Rcd0Tbp4+Bz+E3+PydePoWBjlpZgTc4sRRbwWO+cIo++9O
LvEw2BFIehpDZP9iUPccps45ZBRd9sT1PMGImi+w4c0ZI4sWAuy70a802eANzYS7
jdAjNM16PUBNc2UvCY+dCExWlIGgZpcEUVIFmPcPwZPCr/5hxc0alAjSuvRiBofB
7/XuJK8H0wtvG7xXoKs1HwWLoGkMkdoCzqe6z2fZtVxwCLrjMqv/A1ctdFFR3TT9
tlkSk1Go0fYMtsGFzhvSKmxM7LXeEBdfgulsKJ5mqgEqeok8EuYVldiNLuHoLAoR
ryS+JmFPNqA0qVpaJqJzOZmMhA6/BGie1X37VJ+/7dB6iY93rb8IZKm95GTBPAM+
/qZJm0JTx5Uw3FEXO/GKjuWET07kBdo1PKo0CrNYcH0BmBteL1Qu0J6lNyPs6zhN
9R7ij5jsuUZxHS9xMhI3qm0j59mdFaUZitty6OGA5TnwQfx47BZztTKlPUiYssyU
vuFMDvJJN1oLuslBgi9OCIsLpt/CgdQULxqHS7LkZmgULNF15xIyYyibAALoO1Fm
RsfRUajPK66G240W/ryQz8xO40QhNN09Mlw24UA/l4imkW68KuyoJK6j3bQIw7ji
1YphqtdJEiFoH2lUUmIY0humVpvJSTJxftUSyieNtw6dGjCsELg2BZLt11yP0muf
16dWSLGp9QYven0Dfh5+rH+1qve7HacDenmloHwPxnD1NMaiEMftrTJC72g6dOxo
LSDZwDmshAogOQ0BbtlW9HFTa+vN38OlVflVVN02iLymxbu2NCUd9m+O7pNoKvi3
PdmFTUtqa22fkbJCOiuvS41IFZvYVX5PbCQ74czJYLKh5aFCf3o8N8+PTOGYSz1t
WBE7602MB9zK58MAVv7jXEqkGtACGQJJlgOEolleCIZ9lIAtq10HtqQIefPVf4VL
GvqCviwQqtmZctXFy3U+fKeZV+B9SApxDhdtDqtBXPUiaow1RZMUEVT9oYuJUsev
krqFb+6hu0LrgDNuwXS/U4I19PbcHdGtgeZKxan2VNpoB5rt9mj8KF50ftnSXd6j
tgy0vMoYpsA1BU64oDMVjXMjTAQCHdEm4uOEkxG14pDWfe1B2uI4Bb92PrUOvRBw
CQdGiLQQhN4H4h+1OQba1SEwbWNf9OcGeCJ4bb7v5JQuLP0GDVCuuMayByw7FmMw
CEmBn3aeqbfHUflkSmNeJS0QNRpBagKGNFXygR8k9K7PB7eAxm6tNmdjmRYC+v6h
hvmhH3XwW83Xly3AQj5Tky3mNp6EFKH8EYBvFgN1stciHADXV7kG9vgyCNtIsk1u
e96S6kG3lUCIy9ivSXJiM10Ubue/GT6A/orTSiZPKYn8ddNj+VGgbmnP1nv6APCi
aIYOQiyESWdw7YFb71qayj46G4YUokK3PvjM0aHNCabZL0cq1qkIOj/WUolyOnLH
ld3vTq5iiSso3Yoq3ocgC/b29ojdnk8yZDIdWWWAIezI0Vw4lYB5MS+iynKr7Lek
WnPfv0N0j4TsQIj+GzcBiEkkjYPY0TkSzu7CSzncYSk8AasjeZ9JD+so+sSuyznQ
gpBzbRmiF6QD+PXjFk3PmSHok2Mliz+Zi9/OUEFF7ZeRSrMsz0wkvX0ioJesPnpU
vvup130RYBpx87UA9TjfNbzEbjxPvLjuIc96FTZwzvYyRRCdK4b7h0ddIOI7FhnO
AWduG+ZwTjZ7ByyPRI6+zB5MgDq3dihsZjcCxwRaednCs72uAz9ttKUo2wt9+c7g
x2kQLxzCD8b4FozRyXeZTik6huO/M5zixuf8SpKYTp4WDJglzHXU+u4QO8wW7fuV
AXY4bROyurHaGhZjqfH3dxihsOIBcvACst3O1Onvj7aMmR+rH+jowGXqlDpwe5fY
sNk1rPDTjfSd2+Y9yVaJe1AC7vliv4fGR1rzjQoBS52KtfYiY2ryMGrwW3oSSlCo
BqXHgDbwIv768KhwMxhb666wg/JR7qZZWupM4HZ4xiJ9DmHuupPvnJmIJiZWUrqa
z3CV+TgoygktoGvabKhIt7e4NJltxkmcYr3zRb2ynuc7I9uqsu1xpKoVqO+vCDt5
zIggd8Qus99Asa/28/J5o2EvDq881+Cwn6G2xs7r7R69/xkq+n9xY981VvUsCko9
pM+uQdd4V3gJol5iZFAz9yxw6DYvV2RNw5Z9NFbbOoL7T2TttL4AwvGtxOS9zeoc
Gw+EUboWPBLNxG/pMVpEj8fJ3M8XY6lICzfKYST2yn1UrjMh9qfgH0ckZ5TsiT5J
K2NDql+BtIm9yE9U2AvzfBUSNW9U+Bri6voHSPMm/el7vDVy3nX4UWhgB8UAwB6F
A0UZh8g5JE2yWCRpzbELSFm2rPLG3MSVDB0ZgPENSy4wzdn0H8FQu7gFTIfJ8myP
9zWJjcqnjvZ416MhkaE0P87O1nAJ2lJy3VNS739bbkwsxEv7SJC4yjzmK07S+36o
/ijur8tEZU+d7UNPojERBxP4uHaaRGeBeBGYaVqovEXCfJaOuwPlvB9b8mS9YYLa
YO7d99UDvwDKTyKEn2iU/wqPdyc1k1wKBN4MZbuhxCxzm+8MSEHZSpct+4x/C1y5
8sIA9imjMdB1v19sADUzOyfw8IoeuUL6I0dCik0LRxaidNppDkmlgeNEcktFgbY9
rbc/AqEHJf6cTNnYtzr90/NFeEgMOkV5qeDeS0p48xwHi9D1l/GiPpSNP9TpdBvU
6n2WVB/mUKHJG6SYpFJUcRDpTDO5XNOBbjHGJhNSixy6I2E7puUSfKVGnUB/NzZP
X2+sVq0dJ/k88j+YNU5vcOqUHflknpdf6uQ57bepKNZEteaopfJgRgyprAvpI5+L
ZZVUqZRqRqvI3KtJJt3fRvvAw7SieELkJE/9VK8U2KepxkI4ZVcwqiygkgmVlmEb
tHhd5EmQdfIVHkqcpEY1uKjf9mTRJZXYQewj6ABsUbQqAcny4NMLRZgARqYW225E
pU3/L1F2+hOxl0Y54QTmiOy0Tqjudp2COAggoYpI/OdmTE0nJlza1R6UJqmErtXG
5A8h0OKe8pBtzfN8iIKjBFegY7w6lLZuwhXccwejTzKucK9qh/sJf4OCd+Gvmfil
/N9alSzOhdwsg5uO2aorBpmBkLPXxWhb5bLspltEyn+poePu/mW6KQbHuYd++hiO
nnzTeysyyLXvA0Wix7hBMvQ9KYqhsCP8ldYUMP4E9DzvSWyUCfpcvRfeF5/jreu+
cSznTVARwGx8UD0IuaG4qot4jTkw0swYMF85KuE7gaBqkow3dcDNyf8y60cCICrT
B3C2myfXwoWvhnMyCLqZJCL2RvMGQ0X32FrfTJ+0Ap9eKhRasx0zP8Xxo8awpCeZ
HsIV8Py9aIJ9/1nOI6XjOLyUQL+SOMywgYpt4LIdGDrdKaTm88hNZdrMr/EP75z0
BkQF+UKq8qzDzR4+pUW/D7ZWEphDVV4OIaIvuC7Q0YiyG5rFlqZY7bgEce9CJCvB
henCcIMGS6IdnLW5pcnF6MDjU3npSdM44Iv3hxmtBhUBB8fsOAkYroX6pWYsTdLD
M5C7opwi8vLFDLLyygFKPDf7YItD75BUf/j4mcUcUJDz7RaBG+EUKAd/XUVQhfg9
8PB6MAlkpzET/p8D8nkwRhAzihReRVPZzekpgVj4vNdRrJG30QA7XryEP7M19N7J
0BfQduJwZCq56nc6zZ9leyK04tGAy02fvzgWmeTH/xkZJa9rw0RgzYki8KFu176I
ZyvK8pCXLfo4i6grsdxmqsNrUFF9n9DlKYeyCb3kxN4SOcddojZDqOPZiBENjBXy
JoSzVzEtqMHxMQ640TZecYT6K7Q4TbrMlBeaw+rWjMlX18jhvzs6JKmRXbdkukN8
WBGEPvQLSv3uWzV3IZ8VTUaVug72FkOTFKUyBZnh7qWhtFWjdwHEoBlpZTSCJRks
72hNxfwjP8MAxL87UUjdO1P4c25xV2ZD8JagnOiTSlA7y/qKLDM4ehSiBd+dCv4p
kJMb6AdFmGsDfFnprZIHqb2Rk2J1IY12jEJIR/LCtGH37Bv35Aaes2h4omCEGnXM
KacahK4QFIukGI1hvVNjvX5+UFCEMisw4h/y7tov9ngK/EYH+NFiyt8pbLWg4jhE
lx5RIpPlqahA84c2EpfO5z/+oZilnR6J3As5BP8SeOTLLtzFyDp9MRVrEbz2HQnb
u2rw+0eBTnnhRqBlx5kx5a5rZkUfI80lteYFqchKzJohe8lldSsaF1xwXR3ganuF
ohVnZLRFlyvNMKJtgzfn7CVM/IwF9Ki+/mFxssOxKa/cGFLYb8VOHHMND1mas7aO
HhNB7dzVqsNfHWNVKFVN7kUOtIaJIHZbtp6oMFtddIKc4vT+ILwt4qUFldjjZaGc
G8VCNiMefSxoKBGAXMJPt1yGsSpDic4+dlhfJQzVZx3fIGZK0xDUj3ArabCdGztG
BcIQ+Q8TtB1ynKafNnJNlHzK6LJNeH5PQoZOCajkQKSjFT8hqY8njEq+Zx9QPjgb
UIW4fUMWTwSmo7njoearS0YrDwzvKGzknNiNu2lN6+jPvCmTDiqW6coM1KO0baG6
SpQmxAQD20P7ihGlb/GJtzfM3f0nv53mXetpFMuTXi7BdbjGRE5al4c/CiMMCBTG
HsT+BNdgMALdThuZB2tfmLoA48c2grCGUX7X9GyFYsbfGfo4w6E0/qSorr6YCXZ6
yU1m7bAJL4gaphbvD6kNpJjSKeIzOrvMZj/9NLvWQ1TD42nHfS3GJoqGJB69jF+b
D4lujHIguOaC2dLl+VGPzdnw/rW046SB36C7aCw923BO88KyDww1G1ubFi5VNn2a
98DTgHKvc5kOWC7RByq2GMCRiMlc5++5uHdaAyA52bzLZJkptZm8aul7Cnjq7TJO
sPuGmoKr+SBDDVjSpe9Cz9ykchP+KEo/SCRprENDyLIkcipivQU5MSSxB/PwKTPQ
CYHiwIKppc/6P6n244sGmTCpYhEcP7KdzOUrTawQxP1mIaIVs2mE0OZEXFvBJ3Q5
UrTSA1L7A/4TdV0XpGJXyRexWX5kgPE3Ze44bnoEmV/wJx9JbdVIDs7KZ7u/SLvz
r0jsLhElhiNyknyyj3vGkELdlIBurDyNF84jvL/gB98hME8Erk0DnHWXhwtbvair
Q2zAshJhW0RKC9oXeilR+xwtNdsluKUwXHnvUiui+NO8tBdZwApU5HDmv3l9If9J
q3zb/sMosfyQLNBCq6WoOlU/4vkusVONgoBP8ymOAh47p48S4JW8ZfR4khBQiGZx
KDfG0vxobQhfilViMyoHfgJ3tfbvAbNDp26HHyqGACN7COG4jSj5e6YLOX54CFuz
AJlOmIeI2su1QVp0yLxOEZ13qVLhM1/LfEPSlY38zVTQWE5x3yKNZXWhvqoYYqdz
E8+cYPae84XGmzI8j6XMsYsZuveqoYOzcvb0VWHxzE+Di0M4janj73E8PGiEAM6f
zYxGOSrMGDshwumZtsEF25j+T3yBOVbwn6+LBaopdL224h0CDhozUPqALyj8mwAl
pHCHsziwi+yEk7MgcsWiVQUXhs0EUnTgEowswCU7mz8Pa8Q+nV1uS+dv35Q40vBn
LaCS2QHzbeUWqJ9jRnsmPsMDVZLTAdWPaCiqZDjofLLLwINUILJBRdXbHo72Av2I
bQA/GEH4C1I1oqHPnILtyQEj2AHxxaIEgG6cnf+y6uKRykE1cP6YA/oggSc+2xGF
iaUYPHwIHzbzWflt3RLxgrgKJCgt8GZV0XTRJtVpluWbsA5iNl/IZKSTau1PTA9k
f4CYuYHkobx49ZBUzanhpLLOPQgMXNc8L41LReliEUOzPOdK4IdS18Kmg9KxOqyS
QGNCeswCE3NsA+a/hALItVteP+G/EJ1dRkBbwXJ+6fVVBOTcuMRYgai4Bqe5Eug2
rquM6c0h8Dv2xEsWbqb8kSXqIN5nVa1TI8e7rnQNgDVLKmgmjuIDvSLH52iP5ZVd
Su6jtq4P860qDixcFxeMGeCRPJYaj/IY+SmOfxqXdEZ3TDCFhAvMZDWqzV2OZRsT
DeysDAbpTh9Q2ymcv1YCXxBzOcJ/Kg+nCrKROMHeCQbYOAoOLGrV+HdvtAScCy+K
5e5oNh2sUZCyADEPRSZgzRRDK6MfmxTkbcDGyz9UxsQx6Z7m3tMG6GQoDgLZsB+E
cUeNeabWIdSVbcRwkAwadx4XAN2UDi57AwT/XgB3Itpftrijob/wUNtngMM5r5k0
3VQVO5u2OPeNIgIVd6tp/Iy3DtYWMqnt/CvyB4b/VfosaK1gngIenoB6B6EkdLyw
Szl46OgGKKxxV01TCFZpYhFiR/x4WKVE/yQZJI6QUNVXm0ja/sL5RZEL6FqC9Lq4
fJ9fjZW9cVQC/8qdNa2UoItl93iqzNgPB161UL40X7d3vmASdFOFXgmmKSQPRQOj
Kez1tJthFTeyVk4JOCMtg4l4BNP1WJ/GBxea9jPGmYRgOc0yy2u4SkgnODrqJZLo
XGl9dj6MfDnxnqflfAgP4Ry0tzjCpe4iR2ZXwOiAKIgj5W8sHA6ZRkmAZL5ke4wF
bI4xOP58ZarC4pm0T07MN/EtkQw+0ujehoYSjZ8ONmpF/JiOL9kz7EKGI15Cj+Pu
JcTQtY4YB4WgU/IPvhtj7zreEWR3fY//ccYL2L0kZG3znHwaxBPGdamnT82MuiOk
baGVAGTfM4ejY4LZJpG484y4g5SMnle2gSsktm5oEgxF2O47p12tsGoUO6eiXzJc
tqaqGpidhLh0CwLv2qjo/qM+F5+4WurhGgl73hSaXGJQkDXius2FEzENOl5Vbvx9
zEOF/6LCxPoGNs07eFXPQ+/274iPkSOjxLia0Uj1FfaRomSm4VCqPj3kQ/3JC6Rv
QjR9nAZ828B5FJk0iDduHv+tSWMdz4OYnyAsqJx8fZiMPYqrw9ZySYjx/V7t8vqY
eSL5ZDNxt7AQkRX+KA0WCHARsOHHgRD1eCiuovHm4IqNTq257brZn56zDyjEshK2
Z72pNJOIs5WB7jaSVTn+15cc2vWE9A2boYtiVidy82ymwV8VIGwxZwvDe+5tMQS3
VfXH63uTKsWfAM7AzgOIznyfXq9DbKxYI4pM1bHqtNKdiOAls77IndyB+CxEI8JC
BkjEdEZsZK/easuc7NuBqzYP/q+DvQk+BwbU6CZp6UMyaCJJz2oSWuBwsDOc9rZs
+pD5QIcgoDx5gFzqNPbzWNcZBZ4zS94yP3tSqLzUbqxOlPAeN3XYZ93umRA9/Z4C
QAF3ei8/StIli/5wsWIoswTz4UwsQLpcG5akJFsyu1GXihTnRGOmBb/pA3OLVhjH
nCW9VOC+ezQjCpRxv8jGWwLIEKth329uD0a1Z7yJgkchCdLRmjmYmbos8khYljEw
sRGMPfyz+rkxfk9SFvUTlj+so1fo8JZD2aOBiKhc/9k2GkzAmOFHXBmGnFqacwLL
eNlFYXaMkZTa2wDWUDyZGXFk9Ky08BN1Xm1gVwMFDKwysGyQ/Ftt6lfw4PCs5yLk
YvnLLWa387XXw7hjjXeVYWbQEv0O+zsW9c/CBDJ9ohCmDbKwTobwxKf/Jyl0n3Of
9iwaClVY64F8gUHcUCJmNSB5NGH/hTzwXc/3dXxwOehTHuiVnZbCI7TeQ+j44/j/
CHBIUOYf6IcdRUaYgMbaYn7J+xbicdV+zFgMyCJXTYOEaqpXt4nNasUNmxMzN7NG
QgaHbG9vjxawOtlqAw4CukpDF3dZYSeUbbu6tTDVIyVVqNNf9IlPPKrb3eosMIu7
CFCc/OKNdmwhDhWblDTdcLkGcfXBctEqYeHw3lHaLg33hYPgcmXPt61NHKH3TdH5
bV+lQiGh6GOKtDBsVAxygrUZJ+GcCHwhDqEsXcrizF1x8urHI1SbRAJ++eA8RWHR
qDeb3T4NC7Bs8vGNVnnhJcDDg1MalOmP5cnxSgd7Z9f7vWmODczVtnR3DmhkFb8A
GCaVFDfOalRHLPT0ORhnbncMZ+6m7K/RYfWlzemibvnHCN3ZSlBoWxZI9+Q63VA9
r2E/0NruFUr/xpmTPeV6jOZ5zNudWP1HT2QQpPPLxCE7ASJL5AVMKiHthy1sBRWh
r5X8UERy4aeEUgMFGJkhLSFVhJOjCtKUx6T63LArhgiAXSAUTn06n78/xpamdVYw
7+Ut5XDpKMaUjAqEdO+1MLOPmXr7iLnljQCe5QBMDUpJFdK1Il2Vht2YdLNhpjFL
ShYUNnOt2Ly+s3Qv4d6sgNTYYbSHN7Z5B8GGH0d4Qrx2y7Fn0CD4sGAZxPgEmH3n
r6vo+sCpZkiZ7yzsa+hmEFcx6Fq3bII0yr5Eqc4wSbuppVMmzKTuVCr245zFGETw
D/45khaMr1MsaZfjCA6/igt9fTTNQCGET88tK7oejg8OzZIiglZDxFPmA6RCH++r
SQeCkZtbig0WE13npW3I7EbTSL8KTjYXcTCiTDeGXzlcHy1pd0I1hE9Pus88RG0O
qZNhmfNH8Eua4yKDyAMkIdIjPXC+utCckoaU9IU0vkNSW3WZylZiVrguQBjN7J9O
K0NNa9EibjT0UFr41KsYKN1CY4rtwKXyV6FGz+4g29TSFBKlDIkGIyAxp9pcweyh
IxGo5zkPJV/nyU5j7p9w1tjTfzQ61sCi0j5Pm4EbJ849RKL8W7hkGJBMbXVviqXQ
R7VxJM6M0NxuOhpy02lzJTuOzR9vILUDymNP3RF4Q2j4S+5jmbvNS2EiY8GbK0T/
2M3JcVtpBjzkSmxNV6Cc4Pt6KXo8ODr1lRiMd5BLQ3QyBeFVnNcOzmTBN8l0L9TN
hqQLOHu9grS2Xz3t54Bzo/W8+kWR8Odi4DGJV2q0eZf59tRa+eC2EsXU2QnL2j2z
YpyksMgmBWvE6LNHT5csRhTAoOUgWk8aObexW/wdYx4KEXrGNK2+aaFsYKu6JJuN
Pl0EVtA/ZbAGOtjZURsYdGfUcNY/ir95zzR09VjvWFeCioLfTniTp85OW0W6JWFo
XHBFe5D1g4q9TeidZw3pZJoEfEyDi+n9PMhTYmth8Uc9vYlVEo80ulAhUdoMwHMK
XSjd/+tTW3m9jC774+ndj+LBBw9ILrhCwdp3XIZIlPQ0dTXR5Anl2es/qpqsqVZq
q5Mmc31evh6HiCOn0AHtz8ZhzurEgxoRXXWKpBVPbeRWKSEopNyG/o0gWoGTnvjM
3OYnAqEnuefm1ILW88er0KzE3vvMKWAwxh8r9wd91YmIfCtOczFeGZijlu+5mRzA
/L4OqNTzIyXMmJceyJu7R5j/eUf7+3nVoebokChKA4B0+CjFbhK9h7xT6iP/B7/q
bnjW8pnFrHmxFrO+aop4GivhQjzv8rgGNAYgLm2i+oPQp4OBKxVjOsJqiQsPZ/Ix
2mgwOLlLtnCn9hrYuhMytY1881IiWZfd8ITXo8HC/Nld6OzGMej2NbH7EoHArJEd
PfIqU5Q84w4anXyAQm3yroQCTc//Of9U4R5QmDjOWI2DoEjw8S+dMQ2trC0ZNElc
FS9s/U1f+hFVd36Fq0dbRsZtSMvZgtzWXFq5nLKmBRTibNyXXq6bS6JNAvF4Mcv9
VWBpobm1NksdJOCotSSjfJGdYJ7pLrKWzCvLJ2JCGGYINDu3/jJyJj/0VBgXxS7M
I88CzCUSCfOnuLV2aAbCXlj8e8Y+jJMQtoGJziVXv7Pes7OZF62hHvWEDwesbhqj
OV8W73FI7L44p+j4a2+SGOt/7B9lgRt1nmjwlk4Id4bxcLEqrCZBZf/sKeJB+qJd
LTAVIK3GvRHuwSiB3JppgqlfTeB8vdqVA5KhDDy45PJxwgjAJveVRwrnR4EQPqTU
zjupDdhbwvKy7uA0VO2W5WnQDPtPLAbLNcVSLy1lOBdYG/o9vF6ij+qnkt5HXPXW
Lv31ptjIaAkfcwJWbLWwRJtlfQmJM1oSfqOR25/sUhh4El13z5nmJSpExM0xOmDV
YYrYJe/CIB/VIJtXo1TNRroRpLd0CJDEFmI0yoWqs6QqokbNOCCMGVWrhmWtbWMj
2oq2Rc1YfuaT4zuD5FRyxeDayi2q2iVIk6Le+3sieaFla0k2x2XF7KlI4Fv/wkRh
56kv2h8cp9Gr5Z5Kvcg8WS5bf6A7Y7HqqV6PgarFdAq0sOYFPaYMfACfhoYMyZso
dMFrrKQwsDFittCtGw+/Yx++X/PqGg6MAkPkDMbE3NqYONQzIQCxy0zYIKtvBJE6
1JuwwwuTQEDYqg/Cl1FenQV1G34IUqpSYjej4WWk/LcGQfD2PcBxZOUDkVlFYLqP
JNHkVfF7Q1IZXEL9eL+lLif3Bd7APtgfv8Mm01sZsZDsdvXGyiYG6JW9c+9TI+sU
qUY3vgVAYcZpFq+Eae3G9PQQ6qTQRVYK+z1l5Jx2TIHzlAv49GT6atO1aM8RmFga
2wEhi3VMU/+mkl408cfGqknaqnp+KPvi5Yo64w8WPj02YFggvP5bORnXVTeoAbcR
CwKOrkNNp6ObxHWv7eh76WtcjjLx+CBwCNXnmrLYV7tjxVz6UlYnzDg4KjoTalib
PDIX+iSzXnLh8nJS2n8yYSyzaNpnfj2D5ck7mpGw8bRIqfvd9DrB8q+fVe1gteRW
Sz1qGkWtU4catpndhBT4mxa5Gry7jqa3k/u3JHF1TwFVv9H0eTvfHOgHPu/9oFsn
ARKYAOuyfKcxzVoux1PmfkNk9lKVAzxrKrjbtVl1vfLvxprJdLLT9WyVTKgj+0cg
Msr1CGRdMOk5f0f/JD99tNPSbO77DEScj+GNO8RVoUe+/WtEuR8yz3U5Z4kqI2a7
p55Aw3kHf/fcILPbigU9DuQWtaYTe+4DS73QUyE8Bh2p9beU8dKQ1Qj6n2Qs0ZNk
lstk2okv+QUa1yMF3VIhXzZpbuOZtEV0/ChPB80bB2Jkp1ofgdYWHiVd6RvomGka
FZrAEc5w8IgS72pDGqJ6dClTraQPfcXXUnSR9zy7UTMbFGRh36eFqnvdwW2KAOPO
iHSYFiKVgv4X0YYhTxEY7DoSLpEJRQnsVxOG90NdeQN4NZQb6BF/5dsCceCZJKf7
UArG7Nh23E6ddWcK9Z5ifVjMtfGg2/VoDpn2TW37InkyOzVMvwrZL3WI8Eczv87E
XZ32vtp8ui74WNegbkLJxmrRzNO6Uy+DZqf8IE9piq8iEr4wYsnaCB5A5w4CqJQC
DdKMTkuJaIPorRXcfdrBylQUwTVWvjCAb77KoqkBhauZbVQXoGQtK/g4fi/ZLYCi
nxGNphSShVVxb7YaLa4oqrPeMxZhZ3dRU6e/YSavmEOJpuqcaW75Hv89acd1LYLn
AcUFYUuPwwRJUHrKRnb0TVhYNxZFgOtha1CiS62gBOat+9qcf+yTc0IUG9XmOFnL
d8+aRHKu5SgM4CvzQu0nBLJD/WHc7JLV4Fl2tf6UejJQ1NJUBxRUkETUyGWurbWB
d+Y6oHamnPrMwyDVwoWxE+zRuFsasnGnYdR8UBR6Tc0tKOzFGRe4h8ZlOFBTdgJk
y7kWUhrp5VkJ5IR/+CQQXGE9kvqOqFX0R7uC6oQTZVS+6l+ztmveuUxaa0gGNZxi
yXU0dTNmIWsXI50Z3rLJFW61SFH4Pv2/Vy20UFv2h3iZWfyroSBOPXWRcGAuRrEa
w6OIoCUSdE3dC+vIHiwl6A3XPT/MSGnhVby6GybiCsKupLMbHKuty0LqemSNEV+5
UuN2PkmjozmWtfzNQ8PKYF73Pr3zwGAQIFrPpq9a5g23PVCesbVkK65YFSxGPfL+
8pmmbX7mU+ncLRBlEeg+TPJT4001tB7mpc2jNSkKhLyVDMa4ZiPPqkIwue5zrE84
zc2q2L+EaszrrAYb/Ye5RExyU3kZN21rwuRI6kUuHU4SSvp9bm2azx5DGcKKhdRa
IhFfbZVdLsZ7DToBuOI+Pnf36VlAixJ9PTIqcmbgI4VmEiX36RSO9np5/3nXT5u6
ucEa2n8L/hnvP1m1w1liYVlawO62UgzvrKJDXlJyunhNc933MBHYNImCQ4dRKT/I
acAzAfGcah0dDuxbaDoJHbWRz4Zbxr26F7vMhbKZvNQLI6V7dH7qhXIwjxJuMU2f
sASdk4ppo5/qkcZB9VdP9gBDLL+8y6XXjNE1a2v3MRQsuD8vsxgByEjWEtr7rwMu
mWL+VNjcO0CnKcI92/5rI/gu2nc3OrfTwBAlofZeRQ+z7qeKjYkhXzxhs1ge5+3V
xif4f+DjAMbInx57dO/ZMEyUxS6/XA+JI8I9tWZVFGjw29sMYyBjd5gd5UJc9ibw
cvZuOx0s7um6FV0lQCbXUO5Pf4pf12TCO8vMlHvKg+3LaMNoW1DeInhhXXi3AeDd
contFO9dSPqW+V8lCBv01XK6ifd3CDlpG0ydoqWxrxO2Nockuoyg+GGI7G6XLEHF
Jf23F1ibyb/sECdE5RenPpxPZp+DLR3mbgFNO3djYcF5ZbS2pJ6VO4NX7IKO84z4
00FKEBwxjd08PkTdeSDgop3/4pTLyoNwtuuqIOQQtn5UEckvTRSKfSjIxRxCxqfF
kCSi8MrKDsfhk2iMr6z+MmjRnLq5W/EuJJfvxeGQL8mFwwfm42dajmKHE1OBdMvw
vqLoapWxMEA2heNdAK8pbX8zbVnffql2K/AnLSn4ZdZhEzjN8nhBQdU7MqB9f3G8
cJHqaXMuioksa7r381ndKrQATMTdRb41ZJxTGDV7ZEc3cAjdsbrepvkGRrs8TbPE
A5SCjl7nO5jfkonzJ6dejA6csRU2IdKs8cSI8wuSnb8vkwyRAS+Mqtnot47N37S/
oskxgHgnm3LEgtpEvBhLxAdaAQrJ/X1H7e669DMeCreUjrMsA3F8f+Rj/+hJEA5d
YwGsin4Eese/gof3mVwQ+91bezrsbcf3OOwfqgrP7/63e2l19YCs4LUxRg2AbUMP
S8/9sR6u3cWVixOiebJ0AL2sssug0MizIWnb6m4ofN5se3XbYMWWdJHO/JvHEy/T
7Q47+6vHk/8BZBJ6PnTWSM7xCBJ7upW8Jc8zRHDNI4uf/Ky+UR+zL7M+ALM3b7K7
EnDYNCTJbaiv3S+wf1OlX11aO8uMkljUXQR4/9WwmzhxvyfpT8Ho9KiXELpVNNnH
S5OI3zFZY6mGGuJ3e67leJ9OBO3PbQTGOYhD3KuTAViP4VKKpou+jTPWr366z2uv
QBmpPDqEMFqF8ZF96S/kSDNwF/hhofoWXlbUSZ69jrC+VXLRbVlGGZ3+mbRb+rOw
Ki85pUj/5HeSKatE11R+cwTMeYpTnocBEI0FOXp2LMXZXFiY0TmCD0yieHXli+UG
e8eZgJj2ugIxHwwXcHmhR/QrND6myqydwXNPIQ2fQhPGKklx8UnUWQ2m4rpMfkqJ
GcnBrkYf25CLqWFpZeMNktHGPA9eQjL/wyvF6uea4DCnVIqxoCqOBD1Hugi3VvcS
w/cKVPkxZFi5536YuVkAKABnbO5e0oih6+ECA35VPSPh+ch/fvOiTSVzc6MFpiW8
V1cxTN7MQ8PiAcIgESQY3zuPOgeMLfvhkYqu2bX6Jcl775s3CTqdMCdaOCWXvCHv
tIldzH+Ca7+Vp4R++SeT1RfklyBnkI57LiZ2/j9DxMyIVFEYUIXOS3FZ4/1opt61
NikHCqMmNFoNhvOCcv8pQPSc4NICZDYKhxDZTODlvotOyOSzLPZEBhRLPwLV4Of9
bChcRLsiiFmc9dMjkXqpWeMCOYLd7aUnP1EnllpW2BGdJRv1qDU/wUoMdoliIWbS
nnHfKA+b0wKOoqBHoiMyq6lLSrBU9o099Y6lzEMewfjTdiDv6zt4/OQ7gpBO07RG
ucoLqQb12C+z942NRFVbxTYytq3Bei7V78vL2jZYfUT8bo1ieSwpWbBJlh8JmO4n
SzC4S8F1w8Ha4OyC7pf5eYgve+oKa3GHEu5s+Y1XLxvsqFnQpRPT1e7mNG74janQ
zos2zniDF954CzIHM16zMbgCZawNy16L+TQYRoTAhGLVoieXi0Jv/DyYg8Loqf7/
EeNWod4xq2XdRLJNFvyf9lQeLU86bEttvSKW71vLfTNC7FX56558nj7CSrkaOLTY
GEYV3kuK6zWM4aKGp7JEt1up18CutfDC1rDGp1bmCj0aOz4/J1PoSyE2BHIWwNfW
ZidgNPleYvN0stwqplIEQ4zXYlNM6a6wXl1vjhBr2F8hC6Jy102YDhObfRKd78yL
VqXCbnuvSINSno6g23D6M28WvTpQ8tZpBWJepuVxT33x8z2gTTdvzcnpWl/51SXW
oygWfQPrKVah+W76JLf/Ysm7WVeWqzXK8nDkRQot9iqW0cZN6hKP8xU+GzbkuEhI
oJ2IAKlASDqkDhCUpQIZFnvm0gOHIySF0XJGfyCnRVc7bAZABuPK1l4O+XMjl+1y
2SMAilU4XUxKvwEYmi8/6Yw5m4E9wAv5PDiRV5OXR1lzZjZINyqMedYGi0pGL1ZT
iAWh5A3v0tke3NcA+g5QRX0xTgP5X/IYmv+iKhSFxegSqlL9r4PcG6ppQcX9vA2V
8uvbxbX9zhebS/l1re8+0/ZMVZ94cQ1S540WPdDs8zuPGSRLXonIaITvtoQoLG+x
E4U3GfxE3P9Zd1VMXBgdHT9Vovqejc/UkDc2XWa9+cQqOn9FxHgu7Rivk6qLb2wh
4ig+QAPY7M72i6xInfXp1eaxx+ELwe6mnGp36EqXH/jZkaSzYNzpd5mpg5fFJdlv
FoIi0KKVenqAZCxPjDzNrOCO7ZSLhzef9fektMKehhbbgaPLivK+3iz7/+L0P2kE
0hljQi03K4sFA8nsdCjqGey4CAkh/7RdkNwXaXmkkgf6WSOTidvTgxhObU5FUFpp
HhLQfcw9Fo0FhqmklKbhORjYlI/bUpnzaVVQkWrhoPrzzjcUfgKiwEech8tivvl3
C09TPFU3kvBDfs5o9U/U1jeLg7XyS1JFULi0ngRpwEag+1K8QLijfh/GCNpZQ/kB
PwO1MaWW/06Bi2Rg9o2Lpra12ROMJ4F9mCh2SobrozXjI24H6gGhips806T4Ojgn
JvNOk55FuvEmwr5TyDUlADejOb3RnJD9ccHzwK6V5K7BbILa3rwwe/klILQkDmZf
cIaC2RZrdJrRtzd/q1DsD81dF9gEjvNSZBr5edCnXIzCRFbeBVicsbSuPTvbe/0Z
tJcQkHcxy6Rhv8vOCL1pwh7dXvjawB+99FZKpYyzKxh7WdAoHxFBCnawL2ud0BYa
JMwtdT79iiUOERvIVJD/9FLgcdCRcHaNYuU2OHVXHbFTUyhx8oip9/vLzKgUww0y
HaCz7JCnykREpe7bt6P8xepLyIzYa1LeX7inH7i9TfcsFVvtZoACZrx1qoOeES05
LEG46WrxkTWTf6Rpc63oQdkCQh3dp1mOge5mMxb3KFRrzmlYXysoiik4VF6YRO15
hIhfRsa8k8jc13cO/qDt9gc3u0SFj5SgAchK1G0syJ5C9e8qK9HmhZC4mUYipS+M
YsIzBEegIHW1wEXZcZijY5S6R0NcknCVRXsD+/bkxFW8i7PQxj/nTN5fw2Mp8Ja5
S5q7SWxv69ud1fKYXdmMAHzIELy5Avzz/3l3MA5jsAoqQGE7YgzbSjN3Fo5JosKi
qJpVJHVOgJ9g+y2E8Hy07bqX14gSj8eCZEZ0AmMmjYrG8uqIxbKrXCCvb8PzOKRj
hZAeeFWPPi+9a4mQTjogW4qfhQETUphObGFBy0/PKRFRON6YiSbl3WGnUjCJ46GY
EF1CTefgIRMGgBHX5X/f1MLtkeCiE9Bg9Fzeo6/5UraWmPntQ4pAf7WGHqCZHWeo
cxy7TRnWamE8TsqxfTQ3dPRnEEppeKk9f39GduX7bn3DgoAoeCIt3ARA3ne8rGU7
+SDp1r7KszmU3aIBHu6zQHhYID76RMTRlErXZZvTHOdYYWNWZ9x+vuC7hw1EJSz0
vf1onOk8pIW2fh0l1xmedwwVwqjhS+vcLd+ZToxap65rzni+18Is6nehTFczxEUZ
5ZDG7NodgzJhuXng/q8//Ky7HJreRDz851Gz5XRYAdZ4ySA/yjr2y+knrjC9UA5A
4s6B6hLPQD7SWNrRYdPd2fvWWcjKrm/LFlAxc3V49JoPd09lfM6GC/9uo9GxG6WR
RmLuWoxW/ch/dyzPwBiS4shP4u2VLJVp3qRIXkY4aZSYljkS3O3WpJEAWWBU1OeM
cHYywZX4T2DhC34QAQgIXpIsEydfrY3vLbuZJQadirDXnw6Wg360luiXN3HVSFQu
m+qsNSlPE/zpi75QryfNEd80Vest6fp9ODYaIRKdZtFov4yL4X8xv73+2SLPygHA
a6YA89mSHXJjFbgvNcZMmKG1wRKSH6ahpv57car25vl/x+WwL75LXgzShglHEpmG
ZsJuPkMdy+lSzH0ojUfHIl7uO7eFgRfTajr+Owa0yER6IJXjFrxNpR0eAUbdL16m
AU6D3ifQ1tMBZNre2dijxWS0fCv5yJ9Wn0qLYi/7q9VpzxeUjXtY4+pSt8SFeO66
cZ17ta8qaYU5p9E1bxLWrxOKQUigSck1W/BbhPFld/FLRNDTLjtyaWcsi8mGNDbH
7HxunpE2Vi2Hf7I3eunAAPdov1L8LzHeoUcwgLRrkIirMswZrxP6Fx2owodcYzMQ
mfOkmXDWar6Dg2I39dlHd5yOmcmxDxzz5l1HEnEAZVrJRJErwA891IvrKdrYJfju
4j/5ctFTiHSKBn7vwv6q++hLazySs7upG5kwpT+ht/ggT8FTB9yMcJn+4speEfQg
NAb6YBbmFNAHUDZcdrqU4bGidiwXKeS8eajc+GnOA7LH5DVXYxY6XZkqqBICEhGj
9+I5ZlligRrIg4KByZ2OcZe292JjQ+Db7hwpPBGU/GQY+Jj4RYLq2QwoyecS12NN
RxltSKCFeJ03MQ+O5jgQL7ExmqeOiVG/KxgpkkHsnVPi9vy/4nselwDG81DVjRJr
Ui/kodjf8WDRdsG8Nwx9UE4GJinpnAdhvRZxWr3xSxNz0dqB9yBF0JvOx+vFek0B
TX+XTvYs4cGbfYsjybufzY3fyoBGg1Sz0n1B89KlvbkEZL6L7VdzcM6lAbRNkbxj
i9JZxzRaUIftBtMqsyRGn2FWbslOtI/umj4CFMIUTMwdERuhOGORJXOeZg1ylY30
AR7vUeyuyA0V/Poh+aRBoPj0dnwOSBUjCvUocmBYH2liOVAZJJKNxbJYoh9+OWoj
/fO4NLexCq2pGBI7iZLHd9rCNcmBlDCr6P4jkZe4EbBATF4vvRKfY4i7jjeMr6DO
XhFMh7LaL6qclEIaWcNY1uMMExvKAYL6pY2vmugWN9E4d+WuZhQlUXN3XSvfuQ7v
v8aXwMRnXy782WhU944J3Ty4OUipB07vLmwGzZ9S7U2gadu6KYoW7SWKR5L5F4O/
5xkNfDaF+g+ZJjQsSXsrcCnkqQ5S5bfsZj/50JgctkQ8OcF4Rnsvh1kxFf9I7qI2
7QsTSKz/nAqAoZJ4VSLMqQOFj3bV7fJFyDr+PPcLaYY1wBLCUFptaO2aDFs1bbsM
u1A5c8bwk5zuGKoPrUZU0pkqaLJfdqMmb/Q20Qt1DYdTrCX7jy1jRD/He2zhI3rs
hMJW42K3JnFMVUSVzV+V/zskAqrqu+tn9WDAGBTWr05neqNgyRn5gYCK/ZEhCbAK
iImbH8EnO2QMWo7tDKEff8RPAqxDrr5dha0RVLJ5IRqR0GDq+0BowqPkV+JfwOpg
qO5ISs7WEcyRpkCmu8tksaO+3RjayvAM586PN6BkWNorCwDJxebFTdjMakO4GXG7
X82F8Xrbhs4Mbzt/iwKbkuydTJ/zYr99jz9SdiQi6qOPju2nkYIw73SMKDSKKW15
3qxNUpa6Bi7/txgPkiiG9WXgKq1LJTkeJewFZG0SchCMW2RJDHj+rm3Hrng7D/ob
l7XvCkD8dBnuVoCMBo56vhGs6MXYyLFIjYcvP7tqNTFOjCuQnrItoRO0h4XaPsYc
KCcUteq33Rz1x9ZkxlDu3DkpRaAE4GzrFZWtEQiOADKYyjh5YFbOXptEGjXipVBR
PPRB15gzVuVe163w1BKfiflDpmS2gG0zdeJ7A/oyfeFNTDetzeT8IgAZaPWLk6RO
0WDLKaiV2K7zXesUmRjTBfNeZ/6MIs+XKOr6CjfACa88s8AE62yeSWfTWvhtG0tt
Hl6lJEfJYuUxg6jljt6LQ/1qkmx1OHBh1BIc5NMzYJZWQT5r6YVzjBGscWgnRWSn
uj9J/4Mt9DuYRwmTEsFwR+5rFnZTWWXw6VytJ9T+Cm0S6cr78J1wbgZ5iZCQSiyz
xt3iDd1fDDGpYuHBdVfteMhIbM/+B3RbwMtfucSW4rdKIdi/rkce0cCKJuhoNAnQ
WcayVcybktl3m2K8sjSWbukxtgkq5X1SUQRJzpMz64CL0VkXzsW4VuWxV3m7uke1
5nJa3n5lr2SEO5HosfZt3w6N5FKCD8cA8qEKCIRemKu3g0flaleLm3hReGYxQtxl
XblwU3LkJkfd1YJvwqGNryZhzmbqtgzSMS5LiR4p6MyMlbt8MSuCxAjWwtUKC5IZ
5TQr/QaAZ9S+TnkBU+Uct7E5GabMMVfJihd2JQugEMIqMw3PHa6Glsy1RlHhrS0W
rfHcTDvfn8LMaAEUmQ2HP4JqvG2dtVXNGrjJ4g/vtLEAWFqnQAzA1CbaWO7MPx+X
JLilWXlCCe7AiqftfyDTAuP7363Au2IiADKHjNxbjc1TzuX0FFMoW+B4YR3LKKp/
M6yF21pH/HnfZfmauNxji0tlc6RdimG8MICPO70qWorV/SDV2xNpMAmQcRXzy9Vn
tzJGInEuL265pWcJQoY50j9fTRxltNBL0JuMzmjKD+uHTaEtLDGy4Kpf9Oz2bY4c
AAgEOpzxEFsKzniA4g2t6Vy/B9mUQWwEHGNKPlP54GRya9vNS9O0hcz/9PoIdMVq
ubeS75bgxLFuLAgNc7qedN81alqvwzdXyCKugWYVi+elixgSJhrwpjmA7/Fxcrg2
rpK+m4JRPge+W4nknduO0RCssaotcbZriC3Ea7Ja4IY2NvbjKLZ1EvIOQnoB9c7K
CBLX9J9zPKuwz0DWLvgs/bF9vKzIOUv3cpx0aLhUUKdmEFgZ091hK6nhu5x4UJjL
mkvoGA3KSQVQwKRR39vzKacnNmv4IXsP7J/y/wheH8LZlJ7S7LMI96VRNqTV8zeu
2rEY/vXaasbSfmYIxNRrFYrkBHryODgZCdC+4fFi3iBPEo45/s2lCBd+lFzL4X1E
Se3RBWUfcxk/BvJWOaVn43ca8ZkqOjDJ5ZBh9qCB/SLfxGjqGv9PJjjaaIJfbeEQ
uFrHOFgDhKMazzBX44jTZndCv5T1D/dDt3EiI24LlKb68ZdgTJA+JJlm75sheU1v
4UFgcWw0xkMawVByC3HD3BDKRuAwODETKCRTa2wr9BkwwJyieVvzNKpwy9FjQyTN
18i6v3YCPCcxRMlL/itlhfVymYbphuifAOR0NUkgb1OQ/CX7FwrIorvN+a3JA85b
AHG/YQczyaaOnC5iZbrkqtFQd9VhMEy45EIIvhCZdcuNKTLBQxjf8X+mESODCYH8
CVeAjTHNcjUAnkgEpjo60zhmyICXLITznhzYHTyWjVJSoH94tidddMOC+WfLBY/j
fsei3onZQQ2H7MlhXcIPZzT7ktEbIaWiRvM2Pa3Vn92G1gqHw62OmJkKgsCoh6bN
gxzYnBJTIHDow7DT2N5LQWIBBLEXIVOM71uxS2n7MWLnHwXUeVNtiSILtaKELSHM
uqRaYJ/VXrpX2dAe5dOyp/1LCVxSsvL5CY3182q9vnxTPpuTe2nKah0fUhbY62OB
9Vs458amXNhRRFKWPQf166CvDiE0gXJN2un5FQkN4SPn/wOL1qAKTPfok7V35a0F
Gb9Nf9sv+cKd9HslVCWwZuoAl597XCvghDX0OvvFFCEWsfOIMoEfaQHpQqrzLZl1
6Xg20HCzdKZNbteUZ3X6lMPOu49/116q/b68ZBQTcUYsNOao71697GEIiHcyK8nM
gXSYtoAqAVzH8wyRpkK/Ui6UT8iUnsJ/OrtL6I0n4wO+Irgz+Z9R2m8SnhJSvTXS
uiST/slA2OMDfYTQlJxJpnrrOYhcTEln6QMBelzP0wRz0Bxnt1DfHZkRhxvAZAjg
txopD1T4PI3evr+seo/yZgrwLPwDmaiweZ8eXkZui6CUZ5Nu9BBZeJf9pfpmtDks
YtAxYSXIgRDQeIkQPP+h1elyqZ8ZzHjAQpdV5NI1GXFDEh65S4gTWp2CEWchEEJW
GFs6aNQrXWE54+uYYMQk+i30eXGGzCNMsVAe/e9GNtJPIl2+4o9L/HYje3lr9/Rz
cyZPLWtyN1bRSa9n3Fjrf4YmoU3HPrKaZDLyu7d7xDH7tBI6A/Gky8DS+NY4WKd0
9TkYOW46mku/hmSqb9tLZaJu1bMTCpAR86LY/mBWAO5E+Q8FkyjsFFo+dy9/ySGP
AdMawQpMhD3E8ymUcfuhTha91rHQYD+MYuq+WCLELqn65qkT812xUWQdoU32Pvcp
7eGWTdGhslAwAtphFc99tnUTmi953jZA43A3mfFzea73KvOMLkgaeQlhRCLStyso
yxYOOzfeatl8BOFsyDrQZZRtGki2sknXfIHQKRr+WYijTgJGo2qxAHPVQccMHFQn
eLjEYYHiIdaOVxy9pf3X4N1mO7sZx3Gfh42zBK6Uep+0IRJOGLfk6SfBTFOLaIl4
Sd8CRUVeXgx72Yb6Zb2twwKgWduxNvILrfWTAtYBBAcFS/0pQQZSxmmB59ukgzAT
2g1QR1wWYukyQzJfNJgR6E2R+65NmMuM5ctCqaMk+dUhx9ix2o+LlK0VGC42JD1j
ukxgHpgyXZIKCYgkElkOB3Qyhr+uFmBHfFUyqJVWc76jxBax0/kbOUfo94wGU537
sECxWfPOeGXQZpXf/E506bhvxRY8JDjcZ/m1JSXO5kwU/1OwFo/mTa0RWKOvnIMi
1cReHnyL42Yt0PooMf2eoZsUTm4csTooW3j5gRecwNuOQGLQgB/cMJEepH8iB++2
JdgxoczrlHx9iUffXToqSIOJlSZLQWfJnmv4WirQ9icpM0OYiRqR0vkBtUM4vJS1
FDTQmkKXetjMMD1MUOUCh6Q0gGwxp5dY9Ey2XMsU9jFYMm+c1qzRZTlGjiJcnDCx
9wdBeeIKYs63BZfUmwjbm9HHdQax8VxZqH00hf9ON+SAicgxgdjO+BmizxHj/w/C
XJHgKXWGxGfaDcUlhl0Qyd3SYSCYiHB2E1UXfrMTyoDR4yoD8TC+EOyWABpkqJkl
MUqseZEeyNw1XzXsWmpr6/rQuGjlCV4mNphLvwhtbIvbiAYrD8nHDZkK0OlPBSHE
tvh1t+A+R7n5qaQFd1FabUWXhDrzBsZx4QHWqPpDCX0XOjcJUM+YaXrI7kDA6UsA
uQMfSdL8++YcJaD+PcGldLjuAJVlEfvDvAU8ZUjnXxcPRGAsRfmOaBoBuSAsxmI/
zwFG1gOu3mj2aDmvGjTD0396FDLg6x89wK9Wft5fhubk+se8ipUG+DH9t+WwSzBB
64lgcght8SpozdpivW+OcTOuaptvLTVcPPk4Z1cCmrzAV1g4Z9HToV6plI5SELVV
Lw0R7IsG22VQ4RcLQni79udEIiND/fYG2IjBl0opSYqBGTP95tTj5scfSEwB/P7v
YvEBx/01L09Bb+hm6WdIPe0vOhtck224KsFIEy/QaHbDH7OJRe5EPVqmAR9pUw3E
yfg8qCpXDOthqZR2HxT5p/za7No9ONeecvWS8C0Clhk3jDfBrFLCvcDJ0es0VdgT
mesYKBtsLkeVnIaDGyD37m7kn3+dwm8mH0DK80m85nHepNGqN3oShDaxEcB81H2d
+5WwF7QDl58Kf6ArhbuUlfXbDORNKAyEs5W8DYITYozcbuKg3toOr8J5CzMLXUWt
QcLXTWjhPCtfT3WAo1QXewb+leR7mKygrgIkEUldTnSGAKMVwtDset9bmVB557Gz
TKaC8zywyKKos+R6gtqczGL5j1j1Az2zYSJXP3OIxC6SzFz0n+IDyverf4FEcGtI
h6QVn/yRyQr5rFPdnKpYPlExW2vyv7cWgyhlyN+w2Y2xaq7ICwrlKz9Rz49WitTu
WPr7GPuLoPDHzVdVk4yBFsPzkzNGpAW4Ph/wWlbF7JcGHi7w83LvXMysSONzRz4I
M3wNMpI4dXeten385nMdvPVO1PiIS5CrwQgwz17cxJNbUcD8llkydRqizZaYFH3u
3DClB//mbRSSl4gMVeivxPh7D9PKqwZH72dGCOn9ZwKw1aNoxLdGhzY6YiSvulD/
yrHmcb8GNDW6HFLRQqf4tyE6pU5Jbl9dxnFwVliqOytWg8lkKx5ytvJpTbvrDZVW
VnaL5E8ZroyxSlYmq3QMQCnbU70kihPyry2XdJ9i5wAqQ8csFxE2r0oaFKppuE4O
dLXbAX6GUQ3ArLYJ3P4d/nToBMHmfssCVecL+E/kPUiqs66IkMIk/DRXDpnnmORj
92F2Cg4TXCIXpX02NFu0gmM/8esAwrzg2+nvaVSHUj09Yx32y6mm1bKtLlG0rzED
JYtsGYx2lEJ75qgWP/1KhmlbCIfNnyddB0b6wiAC27Udge/mNhCRAECABtM5OKoa
4A7sIK5gjDhOXpH1uWJ3U7+s7t2v5o44A4FBvOuM3tsC31ByDrEZ4TZbgJTqheVT
xb4wilNtev6xyOtPqNS7nZUNxrCBkH1Wz0gnEojp1gkqb/SpcJ+A0jk4kjyh38Xc
sA+z3S8zQsCoS9r9GVrB4HoZDaKzXETYGvW6siPH+vkXLlTttvcN5dssRP3brNVg
wnFusUqH+2eCZOIQPvYRRaC7btXJWra98H45yU+sNo7Q827HpZdMsPhcVgMWs2mw
2bHzkEWXYAzzXKGdpWLUeuSe1KQok4EEWGqW2dPXEmaVHx9zAxRpKIpj9UqX7AjV
1BlczY2hxSGuRR8hA+BCxCTT7mvu1jSDgPpJkr98AE33bxZbg3CbW3nizthDAiD+
CPHMuINTQOjRiYvx8e7y/X30YkEp7aAzqinlz5kc++oFy42MkSliBiUxBEnn7XWN
gaxKWhkq+FZbwqp/g5JV0R9z++0sva8DLBhRUmfik5G2BkwshprspdjbcAh14prS
wD18cnKrTg9HbndES9x9zvZlibnkwnSkYju0b//5XLvW0WzMfEizNVCxG5OtivRA
4w6KOMe5JuBWV2NgrEHMuJ2LMgmwRCZWenRSM9fzZ7GTblxm/4qzUvAWmDvk2izW
7QdRYve0AVkQH/Oj4Gpfv+GiCRL3o+sHjeXmS5V1BnjBLmTRUihYERZ+YsVxwJFG
NfpaSUm0tYm6bqFH6P1rcdQgisMlZWyPlRC4N9x1eQlla66/fi+q/ihAMAMOlp0v
DXfMVE57BZZwUlVKDh/FqedCaZel3mX0BTRTMPC2T0+PC7GCs1CGFm3n4K5QALJ3
al/CcNy7kSRoHxqrLTdhEltN4zl6YNNyteBGlEUP7N1cM1vlXgnLaIdyVWCeYh/J
krPtjaKOuFaXz+E/XIBktOa6xOe6pWFN4CMsPKKaPYK7mhxNQRsZ5+ppooqKSC2k
qk5XZnnlugPJFOgXK5FPvD+uYTLJWuwqixXMk5pYjTnrtlADqIpDtZl/Uggz1fvG
5SnR3lk5NOfH/FTIon8fcmLhHWpcyvTslud1EnWD2qGWyrsKg/JGrhihQEo3WyUr
bVnyIvLg025FZ1BJNsLAvChPfSH/CFkG7ZyQhK2HzsrhoMnxUFw5pUJpj+04OGFV
cRLSlFcvQc6J5QqR7H7Y0UK1pvo+bLeJyTTP3scfVyE55WDFYy18vMEtDJSK3fPw
7AaHWvtCjUY+9t/Dk0JzYebVSFT3jrswJIxEddyNef7FiT1fssI9WpYuDMhl2XDk
ZNjZfUFBALYTvGFOGUl9a5gcg53X1X22EAqzKkk+3Tqjl3e9H0OlXRjSnFiTZZrs
QPtHhYEQ6OUSKuQ6lwewGvSzgUDCUphrpkYozfmla6X9LbbK0Tmaa5eZRsQCRvlS
FeRTKEvpu+rfPE+d/7XXlifgzAh0YHKWsytoAHmuDKWcLM3I9QKab/NnCT3A+GKP
HIv3rWRjA+tbRbx7z7F/K/EIHzjKezke/b7h4UeyV2GdB9XbfUcan/nlKfu4596M
d+6KRCn3EbV6l51Nz78g1muCdPG6dfIF0q0vPnw50IU1umLsu2LNy/E6vTNwbrAV
+8JW0iRPibQbCdQSsNVBkil2j5tmTBMd+8Ii4YLV4uqwBbHNi9RGa+FyxI/hof+M
djZX88B6RPQ/FmGLx+MJ8fVoauqeNghRaook7959k+as6Ao/hknb99ZuQwwI0bbe
hLnJk7G/zOBBIL7A3wh5M+vFf4rIIaa9hOYv5brKNJueoHcS+h/68G9V6feEiV1h
eTFw6DsQYH7JdCbYow/n92KZCgFzjpFuCPeO+yYZlbVA+OrXZzNPZkcZ/n1onfPL
RM9VtHcPp3ZyGMJy5GJL671KB8NS1VeZTx2HLkDfrkPfzSWWcz9PlZ8kTQaiIWj+
xLAdNjJWiUzOFBSPszQg+XcnxcYGaa5/Ob/0XChEdea+Br8f1fM1CNeKLOgmr5M4
1ZuU+KaefwsdK1hCu6WFtbmWPfpu6MtrYXURY0KCuREmsvxB+dqTlk8Vd3plcMN/
8Miy4dWf71GYDezHEVSGmHhYrssrTsSCeYDUmrWakNs09EGikK+zeLcJ1fyOI0hY
ScsoBweWnK7sC4HcZAqkRvPAMIEpP0Rc2xlcliARTJrAFKZLWOHMPhlYkTyZN+MU
vGg4LNd1BN5JJVAHf1Mur+SAhZK7enECB3XJi3QWAiswejYKUuPrWbF8HRib5apV
5c2QFBdfvfzWmQuAXMUIpsVESmBJ/Ir6+ggV1zcHcygJ96XpoCq9Z31KcjTcay7y
GLlYCrwcMFIfdZ+2ywqkpyjKqIgfr8qAf60uMWl2cUqB5q6nBa07f4YdUi2JXWSb
iXXFftmS4O545JTyGu78ybM48EEJ0cTRV84SgSSOPIxgML58md6Hg1u+E6zmY2xq
8w8IFcLZ8t9DerEbf9FoGCZk+q5Q5x9WfaftRXsnagOo2svUnixVnL3VK2fURkak
6vpfU9Gqu/0r7R01R6L7AJKcLvpQO6JZTDwgMbyhIV7ixYd4QWneiHoaEI5OhHn0
6zgNqE861vGooQbBoA7SwibfWmijMvg1zzotNj/lTK4OVo5iXdYKSR8LLoxOZP9N
pqSrxeenYQH/4jXA/JebV1oVpJiTt5Q72a9VqDDxbKVBo4lFjt2H7BghgJNd83JZ
fshDS7epIK0g1hDQUWn5/k2rtsJL7AjJ04/n60sx8aOpSnxX1uxEmv4aTSBIV5E8
xwEz267jLRFE6dt4pWmR0scUBbovkRHC3/s5oPSHiX9/HB4dyV4J8TdeAP44eHBP
t8M0P0oGn6s28pn21hHwGQs7g4r4NjujoH7RnTgccrkVJw+yTDkaQJRj8EccU9fa
/rHyVT7EpXxK57TCVEYkKzrk9QJ1etOj6jWEXo1gFwa3JKFzN9t1dvY1ZvxRByEt
qYX3+w5sB7Pa0ZFLmBWVJ3HkOKZa3QxGU5gwiFrrpK4fLXujsEl8Uz0IhnVpLKwT
jcEtKfZDtLWxFykZ72M/2DYqycYBWWiUG3m4L8ZGvU9fNylSp98SMYER6v+ZsRbG
s4fAx1xXeD95gxNKuNyyeuD+16MJaH6LtfnKwfmXlV42QFyMTl+DYPiCyuvifPhs
xzSGtfcb42faalsepybLXn4XQ8KXx7DftM7T4XY25xmP8F6CsPHY3gtZpFvzI7t/
n5dPZbcqopPU6Hv7G71LW6Siqi2uxHbaE40SYukeb44dScm+ocIKswwA2WrugIoU
6ecI5KWlE2+UFjCsxTEkkUV4OhKt8mm+nT7VJ6dGsLkVJ+MdJ3VT3sMhIGFdhh9p
P5B+rBp55udbwcaDZq1uLYyUEma7eDecnKUlgK2KPhGM3bl7N3Mb4u+birYjLvkl
XNRiN39eDR/b/LRYon7zoSWvWu3G5qZfONRIlYvTmAJigePIpx7Nt/LpshbAF8SW
+X/1eYvnojP/clglrZXer6bAHivhhA09gLudtNSmOLKex+Xch5i0qvUJWSLNxAEa
a2ZhJvYhIJLspfQX04UyL3EgetDVtZAWKI8aMnu1EmILI7aRsyIOecxTsN++YtAU
GyZ7KDnaDw4kdQxUwQGag0NzkS0GzE/xPB5gSB15omh3vT4pQcWlmBMnsWflQ2W6
1ijTkBB85ybta9Lgo6YiLFoqan0jbo44bgIswDSjqPMslAyKqH34Ina5TAuFoPDc
UFZjy65UD3HC5e71nkJf8HFHxD263sLdPDfU7yBqG1PEmYgtTZbKQeth5WG3AKfp
UuVEEGxBic9n3ynbAWLAMWu9DQgZEh0BU1wxWFZbWm2/HmUpYyWtzBt/0ymbXrFT
2fD4sq3oJBZYhsjBielfpk1pgTNwAAYcLpCPPbBbmNUCPcvIe6p5GJjQiZFXVhgE
Gt8+RK1oyXyUeC3oSlzhtL1DXJjo9P+e5YCtA4ni6Hih4j7Z1XHgns2yWTIzlkED
g+bXkmtXZXmP1NPDQoPn5owJMJD2NxSgkmhZcMlNCQXE4FKXKWgYLGhqOUoUX43A
2+1Y9pQJVgB/TS5XvnP6Hppd/8wkfaH4hW/VMV7NQg+KFEdhANQi96a6dHkJ3JBu
2gj7JlK+k8GSEEFQVArbqYG1fAiTA/WU9yFPkHTOqpIaXRsIVccfrOSd1AYwvWBY
iFOw5RqjHDhwwKbbO6SaaEdbwVs/0e11rqhqbpSEq0l3Bf+wTof854pVFP5Pabbc
O+VJSHbrinmaIKetlyim9n911RACbZCB6JvbGbYQT5GdQh5ofhSmdvruP5Iz5XDm
CX4jaiArpmZdGQi4koWptcgIdjhRgp9aRXu78V+6I7IxJR1847bORiBIoJSzdGgS
TAzAjKvHYw3oG9o3Fs/WhQ==
`pragma protect end_protected
