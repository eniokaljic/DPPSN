// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JRWVuh2gCpOiDkhuNv3hzxle3LigG6cPKHFOtzTnDoLM03YLvtzFDk5EZ8ba/Fh/
VtEuzqMe0TtcLFTDPfEmf1SX/+YadmISFO5UdBoesVSjsbJ9SR180aq3pK7gr8PT
ndw4wcn79FuQyeQ62s/8aiE9WV6Lf+AcV+mClDaVhOo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5920)
ZwrXb8+lWQF/R0fl/Ofatgyg7b0229mHc0prGYZcD9OBHVpa2R2HmNBKD77SUHC4
EXV0uNRs3jQcGe003KwSpJ2Jw+fMw0b7rHXSSO2uFL4XWjQYMF0rnjTF+gpHQphe
FsHUcweNzLL3kJysKyZy8gC3jkHNjmPxMH2irXa4xX/HyFIR7i+XxdlVxzMl5b2J
5EWWUWqTaDlqJRoDAfCUgOKbom6BxexctFoEEUunZpgS24uT81tKdwu7EBMobU66
4HFdLgn4+hqo7RnIlpsOcCRo+M/TvO4W4uWpNFgfjU1i7c26vvSWRjQqh1EwIQ56
G9PmSFHtgc9gPysARlATMBI42K7b3fuW+PPn4UHnc9bjQkZ4zuwTUzs31R9orxXf
Q0O4T36hnE2tQKW2bbtvvE8O7TW/hfmIkRbYcMCcpU+ilKBY3l44LYlaALTQWrP5
uJnh5XGb4MD16zgdSwsr5OkzyyFs7ubAiwFRGK3MoVqkZrDrrZMAumRJSyLw7m1s
jd3+3Bd7VtQFXnJ9VH6DG/XmKELC3E0qeRj32PjS8lOlieS7dtVS/GGr9sFoPr1e
GqhoDZPcGMzXgPcjEAy4QlDJhpjAzr2RXrRrtBDZ2Tt/AFG/CqR77X85fRYslcOV
H7ekT6exAJLdqyPal1uKgBUXsqGiwFas7LT8w3UPKy1FcDJ7p+iw7PH9OK4YCg/C
9OJr7oyoBrvgEcHMld3eF7aIk+NGimmgCjHBh+545tZEFD95y5OH/m6z/QigGDUt
MmFVg6RaEyvUsnKrhg59ZKIIrEis5+ik2vQWTC2kdLsggBCFIfPaivVrR1PFvfp9
s1mQAN+A5pm3KjrjMPrQkIpD7+8XaORB1FWylz/515Pf845itVnOSrn9y4wahOz+
WfmhBEDxfrsMS0LNgo7/dP8wyWHkYm3TwVwfVEpYlmOyNgG/wO6k5yUSUBlUOsAr
6XtNb926AUk1BXKZCYUknE0wCDBcPjUMKkWpOo0WY4tzzPgaV/6K83wpIgs9621k
9ea9eoIJPzmLkprm8Vld2rfmrb1sCAVze1ECyD5p0rDZLO081nTbU02JjdtY2vPp
Lw95XBz9RcDKzeZtHWKdceOkU6fI5znsrE/TQGLgSva/yIHaJY/k4tsIhcoz1WLH
yevE7Hvfw2r8VtVioQjAHulNjzblv+Yy+h6/C1kgT263Y7rBTqO21ItxOicrDIRM
ywbtJVeKFf0eo/KiRk+K3w02tHIsgs9HhzeSalQKd6InMJf4VgjioR8QEcZaPrgW
4ympBieabXx1oXPNya/N2XOIvyhMyW2IM5coPZ5QykOynVpWVWmtBxhWoiVqYHSs
xOdKZu/DExMYBoFxzsRh2/fz9+cxiaImCqSMwHVDS3FhlXBTrjptNenPC4lssfZp
V+MCZvj/jrtzKlCD3GxwqtAL1XPoS8mdnZIC5jyOhHrMbE2gZaqCVb7j78yMno/W
HSWFB4erZp6hIfJU7UUMZ78WIiINjWoSnUVNNWXlzSOyil1KC8OlSeOAIWdqdxC8
arxjTGY9bLI5c6+RhDrd4bmVFPrR2vdouldATWMfsul4a3FTQ/FKD/LSGTSyP8vm
i/r2/Re+T//D5l9YHaAPIyiYFfOGkJRcl4ydNX4PW4g7GXb1ZuGe3W+SVD5A/pNx
Ht3j+KAQFsELBDd8p6fBzwaQ8wMNbGLCCn18va5am7Ah7QCrB2podHT9ss8AWYjO
mlYl5X+4sY63DKnlVWnsnG0InZvANoB4sOTfOdB+VfIaZ21bzoQQCGKZDsSPSTRy
a3nANYoLoFvqdnhJRsKL/uDKkhDvxlug69t/4H8RTI8v35Pu/lyo9DUFjmzw4mFd
IplRWsMhXAwD207LTiIc/FU784GtfzXWu5Vi9dC0hnOLVjOA4kn6r+f7WeWa2z5V
QqYmi+ShN20wvPymIZodTWw2gMKx7EOBP2dMLBT4eI+p+39OHaVdMHwvbdd1zRS9
HqkxhUqTpQB7RIA/nCEjXpWCjAEKn6BMax5fiTHD8E8+csKnjBEzeXkyHP0RpMXX
u67MAYFDA+05jjAHiUWvCBtcbSUbVUzmAuiWrFiTlhcPRQqYI2THS5AE0q8Ysbao
xsBqD2YbJTJo9SIJZ//qxb5HCLU51EZaCQb5v3KWT5JBX1T8iHmBDgUA/6msxE+Y
KVEoXb+U2/BPXqgRC6x1CksG8VVJUzLWu3gN3vmoK7KpuFatJME16T5tHi0VxZJw
oqQJ/JSZ2v8Qk1yBBpGRjBX6DFhlyHnAov0CgHfMhEpAtEoyef08bYpCWdaFHMqa
s2dK646YAoqPASd2uaALRnYR2Lo5fChG6xm544RYx21yApnSAYgpXCmR1zYia7xY
uBl4DI5RfGpwMBADezULs658RRLnn9RFsbeirO9e3ky+4fm+kI97LLpuApN+0LrB
kLQESerHCL55SpfdnJnXCGB8KBfILqAX9uswW3aQbvipFoxpISOrnlVW5O+iYDYG
Fn52lS47qc7okBaZzIj3iA+PFToWEmAslBWx3z8WrcG9wPEAoMHNkeMvsIDcQc5B
84RFx3cUkYJfwWa+LjnPZn7RqFLW3B8+PSFKu0zqTU3cxkT16nK8mJZx3uuxK6eO
s1cbQCJ7SIknO7UVqVmwkB6+qyX6R3s4t/6k7qv4SPfcT6VhL8nXosXH6GId0BQa
yvpeokpKsd0x1AFbSjese/B5DAoXzE8QP6HpZnojWJWuMCDCcBei0WE2VyILurgd
C0fBh3pQyhroShzrg0SaUXlZi/XG7Z8s8QNDLrrJzMo43WAmdlkpUSSj801SiE6U
dWT0Ivtf6FK/NeqAoGARp5uTcgHoln5yEWWtDRM6ePa4JeS42B1AVCbUQkwjRIam
YnFhesJ6GCJwEjx7lqvk4xAXXsE46fHWzHvjz373rnSofTEfOTbdBbetfz65n4u9
ynJ07wJlRBRirEOCSN37vjiRrnxHSmiGPaEbqsgPp8oaTF2GPaRQz4nOQTOcBnCT
JQvqsh3o5pN5HUGjL5atQfGVml9qZe1SXoYjqDuYmO+uZm+SCbbti39Kd+jjGstE
2AyyZvcRrTnhdWRDrigzk61ZfnFgHMzOxjFLEPk0tx2IKsEsWGI72D8oC+WHcTA2
BeY4pOC0JIr1LwM05K9lw6OZeHM80MgGtVAk6JoDhGjZnzmTl5X6xgjrHH1Kxpvl
4zr7V1LZaYSaJBKHx6eMjC1g4IcaeAO/i/RhYGNadmaCqJvvGhNW2uxsb7q2u35/
BBoOp86ixAbCqu+S/sLWhK4dpq9iNCh69Wqxjj2MgL0/BAetYz44BzJn9D70PvLU
1FdJxuxx+uTr86YQ54FX6mzu4tIJX/zumxRqxKD3SwWGYEzw3bBe4OKDN5FJpiki
yR0RRafoxpzL52ZeX8ob8g7xy2mSpG6bTx5sBrdH16udfF7H5OdJU4SQH6k06UPZ
Aq5YGUzZf0KZEWocz97F4Afw3N5nJl/J3z+CFVchFIqFfiK0COnQnQTAzXnwMtax
67ogn+NFvbxUhYNTXC8uSNXeXCvXJmhqS0ND/JA8RO1xUDzDY0trrXbnn1Kkhyc0
zWx75TOlBQqpWwhJPYBHq9m2GP8++OfE9B5aOSw+obo89gNNhwqkaVSe3Z1GP3N3
72Ep2kvWoJOza95vHxU9Ggmg3jL0ePdpKGTj0uK+Q2hAH5E371PosEerNbgHSfYh
4IfcoZfOo0tIgAurHQuH3IK7S8WMYdedfX2pFOLjGCPmT9YJjvw4YR4b03Z5i/Fp
w9QYkGd38HvNJasAC4UrGpPoWVJbJW4whX7A0bG9Xd6QfRqBsMqqiVIEpHsD4lge
9BS06FP0XIQ5Il5YEfGAFl2ir4IH1nQKn/9um2oOGEOB1QN/7sSvtQ0C4P6HHuja
mnfUDZl14BBVLlCfPx5+jNE8/QQN8310VAR/u19/mS0x6QIEoknQQ0+FWR3O8Yzf
z4RdtZwWobfW5esKNnftT7VB9JvbDJ4lPzjreA7NUorfzaKgdcexxFPhcuxxNx1l
1A2We+iklzv9yo4OsBRK/bX8D6R+tk7yB67tpLpLv9J1YRuu+u5OwYgB1xmptyr+
ufKf5fOqhD5p5aoZLjox1tRney2MLjgcGHW1HAmen4rhmdBNa/jylzqZs2r4QHFB
A8kB/JPA636HPLwH1hJQlYycOg29fuj4SUZNfL/LiFgRw8c+LzcXd6Jdk/g74oCP
zFsUEkd1Vl3tPgWWoM3aJGERGXe29kX9uZrKaj0Z2oGSWj1rze7D2KboG3AvWhJn
qsyeoICKZrdr4eH3jhz5PeRE+DSlyHoj6JjnfOk10kt7Tn0Slv6h1D+UXQzn5fep
KDJyE5xxpKhPNNBKH63K6AOdURt7cmEDAursD9XFVqrzdPFJGCT40/rqJENGpxwy
oPCS/rpnYKXfB5BVrIfNIgdZCv+5H7hmrjHvrxUpL+Ef2pPiZSDLTz+CZwZAz5K2
c/UDmKyLIAmTFmWxGhGhm4vqw0QJec0oK60jIP11qp9DSBzthZvUoXWkECDVc0Ae
03TeNqboUN82+Z+CZFroN2tlX4elOcyKzS2nL+UVUtNYAGWTMI/uBm12unOAC1+2
X5mptuh9zU+JoMvaSEtvBggzCt9JgJLRobb04ZuOn4nIR0MUok8r3v14yOMOjTAU
vYAM4Ju0RIYvpqLuBAmBntFV6BK/bGvmgo/XNIjn/6xRupLgMTGfqEjjDpzx7Ed9
ZM7dEsUuKPuMX7b6gqxJ5qunF+bgVyQG9eNQgR5LecDkMDCevZ15HMGE+pos4R0V
ut536NSRvp2rhx0GH0oEwxbJjmhgwLYJdUcb+uq4wtu16txxBc4HcWGk6Vwhul/J
csX8F4EsiUo7oLSkLTozkbxVEZhYjxbxtv8SbOmNJtk/J4/oFFvtJGncbQ0ewQUw
uXK8PKYCHuGpA3i/hNDc3tKuAn4ZMbjOzgZZ1yTVgpd8pQ85U28VoKULBKvy67sp
yOpkRK0d/9fMlDhPHB5bCNqj2YR8N2HZYug+YFAK/xtnSRttvpuAHjcbbs6xv1mO
bBY4ig9XFBi7SgX8v1lc4dnDDLOHhlhEx3B/xUC8ShjncKhwT+4JD5Hi5+m46siQ
3wR/J9w3jR240Q1Xtz/xr+u422labdderQKhoqjefOoGBrvhBJ5znU3lPOXla41b
oj5eApmlXDDY6C3gzz5kmBeTW3MpIJNBfkFKafUp+JxIg8Jr9wLjHwRWCIAOF/mx
wHRdmYqut5YfD6/PV4eEUfyYp66Zi+zIBVP42qw4C13uELyGC/u5U/MGBlCFZnnR
JfpmxHMXJsC2don+xdDSZDhxM3F5C/sh8ZERmKR3N7WHRf9mAYzi3IadAuXVQn6p
39XmkSacf/IZuZFiVbxJwGFv7YqL+ACCrT/pr0AN1go0g7ey5DKMYijo1c4MCuo+
M8cIE+8D0bNqsm0wn7ZlFGnoV2mfZiJl5whVltvOjkNkKNNPL85qlF3wArN5ZwY1
u5Yi7+NUpCirTZQKknp5X+oUeMF+7PhtgWEEnGNLjdOSL10nJgUHHWyz8Oq20SB6
gtCXfr+lEeMHWjE6KvZjeMc0FuZ9BqDP1jIgBSCzhlOorAUsjKtyU1rwsFTkFvxG
78RUcg+oJ282Y+TolgskyPNv9qJdbDjkxOMmWUP0y+O10DLj+G//ZoqrKVNUA2gY
WCZm3CW72ZXns4+7TrLsM/U0dZlKK8lEIv0vac2VZw/WygzhcJdVDrggvGh9Ewlq
RAmotaIAqCXlqCbQ2VvOCXpGLlFKXrKt6WHMywj1nOpnWAzn7QAdzZiAJULEE9qw
efyaP9R4wh2raXWLd1clEI906ll82djbSRWpXay9aFYHWFRzMzK607fBpsFe8lUJ
4sgov3xPK8c1vUdcXKiv34HKBSRtp2Kt/T1iZkOe6ePJChzJALua+5AywYMjDVdP
woFvpgtZ0R4L+GYB+kDf9uHDN9vrtITLMzOOBRX3WVRjpulCRJpc2zb/VS6y0RUC
gRScyz4GxG2a7e88yMPCM5LBX2peZ9+YqMOuDLWr+qhLQ6pDxQFIp/wwuflNcWJh
FT4T+k2N7RENY6PoeXAs6bFghRi0+VZqU6x2qvdTDTcdfqZYL3o+3Ob9Wwq3smfK
pA4XVeHNRQR0zvJB9b8q9Lq1Y1+FnoVosXJxOiAe3nIQrVQHNDy2ArYKpsZGIteQ
t+WEUrLhz7mnTtfX+3ULD94tGfxJ+C6JGj3Lk4XyakCVUTH3O4ke4ih3/6preinZ
mFaSOFIHTTsAPuJua/QW4mfnjTQ8P6pa8FVkH+89MRvWnRLPBHNdwSghZwmC/m4M
zw5ycyL1rE0OaLRy864ohnTyq86itAdoKqga7pt8YEAUDW8m8QzPE9yjzayD9yUE
yqaVsaiTpCMKiLM/2m+wOMWEPfWuzVO+tiesM903tmq4vFQ2fV3lNUQVoAM1gD+J
uMaPGJ0w71zMGoncEv7r56BJsvUAvhPsKnk1t+WoUcfZwQ9EI10JG0E5eln2gxTA
mgiF8pittC6xq2Kl+4Kp7cOlGAjA8Z/F6h2/X6Xt/38sjS1/XQKoeBMjj1vKKYbI
VVcA5X52TBW+W/xvG7R3ixIEtogG190YNDlmawxG8hW32wKDo/DjFDSM4hrND4Lk
K/2V84aRfrv/fNb1mCVcL6eec7Tup5Ge51GuXjyr1btkaLjalgPTF+IGAUYx3qqT
B03edoa/T/hPaxB9Mxth/fgpyFDCyFFKU7lhmqUDO4MjU2/ues7DU3A2PnhMOxWj
zwXNzxae7mtT/osjIgrVxiGS26z3ulmhK6dznqyYy3FR13CzDsBCSn0yzuG0ADUF
u6cVzp1bcHTCpRLR4gLuaReflRBMvJ6ow0TiiQHzRDxDg9gb7bKM/X5ElijRvuVJ
4zHXEtnK4gYuZyGswzA/tKteOKtFBJeN/G070cvOOmfxgdLBe6Nc4y2dZNxEPtwB
845OqvpD7yUkhgdhA62jMzzm27zN97TX03cfWWO66sMylUQcWwGnQZaB1mOtL3Kt
zB6wF7GxClqeOMIjyqwn9zcKWoPJLTHFzeruBq1VgrD8n/BWFK1UTOauWJMq8bzo
yqzRFtzYhqSQP9JODjom89kEDSnk+vi+JQhp4DHqu4dZYlmwyuNAm47urAT/InOE
SLD0lv7Yyrr8TKL/VnoXSurQUG+oVB70zluGLpjbMrO4kc5Z5tDE0pCo02ULmqmB
dlPYxwYSPy208lHzjtSqYqL1R8DmJyYR9ycyCdOYsyamXTOdVl+WvXuXpSRO2F1L
rNA/22CFbJEKoyG6caEPBG8DPBh3uDn0EACbWMkL9aZ2uEfhCjVVK4L3cbO5y7RC
ilG8zKJ74J805MGCVIt+5/+le5AYxbeAdby1zlRwGRZkpVHoOTrUaHUoc+qF8zfR
/BTv5D7vAMixInGWXZaKIw4j730DWNgE98NHCZjvnb310GUmox5QVo4kMm9Spay8
ywVI4HPkDXLAprTWGNknBw2+hc0/16rg++VSHTcc7qoJyMwfI18BMHIOD2d/d9dy
FKYbrJq3jMHjp3NNPcHKLZVXJ9bkmpxhwGgZ9BkO2NuJ4YjHI5GEuG6APJ87kT95
vvew8eSqwQsHhE5KcA2/voiF+kZLYaXyJKosQuDFzNOjoctQkQrL/zX3en7ukWJC
TU+4Pjd1DjpfSef2iasni06pRTLIFZUPSVinPq6/s0jCSpT3rZLHAEnlteft04Cw
NH1F5r5p3y4Cz8pkEvLPYESHDzRwsv+FdScqmzsj+ICpdSTgWrDBLkE1ClnSWbnj
Sj2VMaRrWIZ7+hNy62xVXp9CQI/PvJDBGgAqqx5ZuIBafRx9J7AAf9PD+lsiY3yc
iTG5wtxx+ugpuSrNIDpbuw==
`pragma protect end_protected
