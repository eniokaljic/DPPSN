// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hc5ylgEJe4IMXPbvWzashxOGFgALKqlBnsbxcLKEPMZ04qX72GIQHkDd+u3bvbAV
hcUrgZ2AdorbwB+stdhou+RhZ9B8S4YIneiJtXb+0ke7I3lStZMVRhwDHH5xCqRB
UlXjgOVGf2QRiXs4ft+lPYlL/1ka4Jq17DsFOXp8fxI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3296)
B/Do/IGbxGOo7U2pSkqHTxJwJT2sJk5D8C96cG3Ksqal5gdMjO36jMTSwbUv2E5I
5m6pfM2SdMc38clHnOn0Lxy1HWK0NoeDYsZq//Hme3j4Z2HhiIEw8yO8OS6vxh1b
2pZb/2xblAw/H/e2Ix0EETkhimNTbWCZZ7PsFYAwjFnJqfLBBNp4inzWqRJ/72sM
QoS701XEMn+stDffADl56aTDPHV79D2w/sy017SEzO6H4uJ98eznJYMN33ztftxB
8DgF3/ww05LlYUR16idpY36apTiPNCKx8GRdU/7N8H+ZtVa1+3YyqR6hHhLX7dt8
FRMJCjGiKlkEL419NROH26tHE3GteWQ7NOZmNoX/AQuK1J0SW2HJzLAvIQB2Qxo9
J/t72teGxiHE1gvYxyA9cnlYMtcyHWGACQcsFx0/Jy5jlMC3+F/nhrt11KH+d2G3
ueJ8b7hXdRn5/lrizXwc/IsvnfuyRp9BtUB40awG0hI7dDJUnwys4fVQ4FWzr5SI
3fy96MHkCtKmc9bc1wMH5AsI5vrS41e4dCTULo2Z8b7cnu516S81wwKuEppv+eL/
1pfhO3rX3Khzp9bmD5Fg3R5KmbRJWs1EgBCWxNsOHWUnXqegmDAVnzU8sMlhxonw
tKvv7Ix+aKcrW+4q0cHBIOHMwVJf5tJdT6VBcJ2+7/IiZUTtrC7GB1gs2p2w9lfy
Yhz6qztGR5mzAgYeDUK2/73UVbHtUzEpTgJCdsSZ7XKiYTqamq9wAgPtiL2D6Yrz
ricf5YzEn41MER5NABvO+u67TBx6d+tDYkn6AV0Rcl1E6kdLeRYKH4MbRl8NkNqg
wgcaxlk/3IF1nubH3h42/mpln1kf1pP39wDQklmd3AMjWsJBoTTTG2x2Yl98Apaq
itQokJMxcEWOTCstoIveu7gVQ1ETjnSiW9+ep5YnLgvT+bHGAc/WG6SmRRBNjE/t
wjoHST3H9+X7L4We39S8xi7W2EYkTfwjGR5VD/4Ds4xOrgOJj4KWgNdWNwn8tbEJ
FWTqIpcDnUzpehIwnGOob2dzzdEQjeJDLMWJsKcfEjMRLFB/ITwal86dZRZCii+8
DvvoN+ZAr7oKWtWC5Th/iyipZiKBx0tl+IP+QSebDQ7lEdfr6KyNa+9YyBk/eEhM
tEQOOdN/dj2ZaXFZr3JYCpuJCt/WZKM+ob9412Zx/jo8XnMb+EORedNvpt94TrOr
8S4/oSjUnfqYU3qj8kq0kf4VQ34iVU28jOBmAMODQw6yz4kA6HmicExXiMp3ONnA
bznzGQIkw6OS/NomsqcUq/InhyJU+2jZBbM7ebaxJ5CBcR1MsJRMCCKzjdwwuZII
9GIvrrYXEFiGMzHk9+KPQ/rz0SZivMMtNMpG6fv/XfH05xvT9fYeM5A028R7LsH5
BWC5fSsHhAMVqz/oSH+w2Dd2JB4WxH6kIeDLs/8GX7sD+O9gHqLymOIWByyxCX2d
Qs6QGrsQZ7z8t8SdDXxDs/ZX9dYI0ElkB8CVctVAzRbiwCdlVhP1TCii3om8LtaL
R2h/YjTZ52+1CvTNZeeXq3IeC7xMi+V4e46MA16VftarR1qAfayNWjurE4mT9os0
R8Gbjy7hQzOo7Hge5jNewokxSf/HTYsTNwVqhVzN2DPaQjhzzdHGdFXN6v+YAqVK
xeWi+zFrUVSRcZX2wV5GcntceMbPEye2pKG0KaR9ScXO07sWSy3DfkVTsUiplCFi
kQXDqk5VU7+8AbAsiOE/YT82xufSJeugckidZ4YrlDQhaz5z5Nj6lEBcELjzBKpD
x+TWmFyRQYgu290haMil2EbTzl4aCI/UkIPDpBq2yiHpWJUy6NAOnbqYBINAM9lv
GEx3D/TqVC99v56MRPAwuCbMjEMGkIB4msVWzRbiTlA9fH4NS0ZmhXajWjX4quoU
7tUJXfqqvzO4mD50CJLnmI35UX32EysG44AhjEFEwHdQuYDzXtgyMFg/Mfh/wIAm
/IT3jV2AW54p9ASaNyA4cmXCzJ59XjZyuqgsJ5uyvQ+nmMbxzuD6ISdVbbylmBf1
dBaVLPHwOuTnx2Bh+eIe/76N1LC8eq2THyq6a2BO3yfjUI6HlWylQIYdv92RAILG
czLGTGTHXMVaQM8gI3A4QcYlO/4GZ9A3NRIFCO2BWqbb39JpRiCOhg7w2CGZ3wiv
SOmGXQxYJU9qGfPtWwimGI1Wx4AG5LqJh2R1nHAjtbnfhM7xeRKWkfQEJ77/jD14
+Y+D8I8jQntuCj63aRULiO8Nma49vGzkAzuGD4bz9RBXFwHRWw3Y2invYxq/OrIy
F+//kI6gw6qSZKN59965nbE9EnZ3RRPOA/awswRLOlVTJGuNB3NcIcDSc2b2ucGA
NNcFXKWlEAd46pNG2i8jH/aIpeN2gRNT96Nl2P0lKIgS6K6Z6bJKcnhVgyO5/6Qx
UD9fKurz7qdMowNboiuxWuyVy/jdGaFatVTGq6Fjsg+wbrT646lADnvraHbxsAB8
P4qf+XxA4EuQiwYjgIvIHVN8zXyfkgz7sfrz1BhUU2OYhrD9DGD7teTDXOMOZS80
7KMtqgBgNAP970zf5HLlyLqGmdC7jJpiseRTQuuhPXZgzWjAL4fBqI+SxDQ8yCYI
W0d7zH6XGGVQ+0cCIy4+TUy0SjkPbFukGDFyqnzVR/TzibE9BkSbg/d3AuKx+xxX
1JUtrVtzbLxI7hkJ9P2VRhHx4eKixyCuA/6emDTV+JjX+s7VmcFERrCAnl/OYOtH
bNPQEMV65wcSp/cY2vpNtiOqAEDc3We+WAizCrtIKvhM/sGMgr0TKGYB2vfdySSC
5rloZ0oJ5KqnXEgEi36LFPTgW164LR3QhfzuVn9Jt0+h1EcNy8sgYcN7BZ955RgU
o3ayTThbkPqkRo9uEQqtN5B0k7cHgx2GWh3Euf6mcYKQE/YsfqNuYdZdjow7lE+X
8acFELcTVIWAl77wsenUo4ksgYVz4eRYSD1w91mVge1QuGOejkV4L4YRz1fT4bR4
9laAPWaUuSjSuhXb0XAdUyG5ivp7cDvE9VyOwpqnslS/KQvMZYgTacb/TIne5xcu
VqKgPf5pBI242IGUAVq6Uev6YuD+e3/k4X29FLjQf1EEb9MuOh7rkqlvJyoGc4TQ
m5akyHLUTU25XcS8NYgDiPXyjmx/Z3d/2xvyhVt1qsf4Q0utNilsp1ab1s3xAfNi
W0GBt5L+omAWS1LU1M3KVVGdm/8IJpBOQ+Xh1dz19LaWuKBjiZ5dzgF+Ja3bC7ZK
6AStdHtsODqI8YgoQopMpH75RjYUw4cE/59H+UnOhjHQNRtZVi7/maT6ka3PuqKk
zuy09xL6qvoTVizoLNXC1nnEicHU+/iXp2C8kEUmu7+WzuXqIf/wIo2tXTvaGiqz
cGHAs518G2micyP6xG3rEDgVzBhGBal/gUkm+zl6FLEJinPWw08mXolBJkQz5b1A
/72i0AkGC/zCZZKUoT7obV+YDPGSRQExFXDe+/qy3S7s2WeX6dkQ7BcDQFwmhd6/
y9lGNwF+lExU9cKvneEUkkqp9c1RRx8XcBzOjcSEkQPcC2yw7tSELk7NlK1kskJp
Hb9m9GD4NvA+24jT+IABVtgSvdreMo5cIuvq3XFcTURLPi1CE95dHaHqot/6rquK
yfa88NOXExdLHnXu5VvcZKhHGf7LZMgqpJVIdJXm1JLpy45kJcHnZWIgpSrwDb+w
4dDm0SafNbE7bmSLwk7P1bCPD/PYVgd2L18YhpkUC6NN+KHfMm+mxncG0dL/unen
CQnNFrbOWvvG2ir97InQKvdZxu/wl6ovWpXm44tZClAx8xhOGnnLqP813S3QwTX+
iIkmtwyV9gRADO1xvZ37hS3BxIKwRmP8kMVXE6E6OOCZPy93cc0BarTJLak/3cvt
hl94nhpca16juqRLFwpS483O0+XFavPjwLSe7DufTrniP9whYagjbEYuYibBlqJz
IcNRNywLPRAfsvGV0WkyMA65ydE9t7QZz3/UAzTFmFcNSAt+jOBEfEM5qHzDnT8B
5lr/UABpd2+hqQ8gFYSoLF90LrsECh08mYFuvLqQ/mUG5XhZUUvRHzNgda8pqM2T
MStMqgo9yJ+Lsws/pu7R2r189ozCkYOiN8Fz6eYqdTjJyJyzUTWJxhugKPjrxouH
4oGDJ0FI/wbZRNaGm8ckcf4kshO9d/CYw1JWd6Wl82CRpamQA2uf9ajkTSBkyYyX
h6ulVVne9305QlyjmHAeOpJM08YP9DD6/VIq1gJpc31fvbYbJWvluHzn93U1OPlP
Jc547Gsv9J9RF5ZfpRBJy4jmc8scPaG4EGwU1BNrUazUJe7Z4io9xoS+Xvn0paDR
YozrTfa5R9jSrBG+i3bM00e4E5ZUMye4QZj8zj5W69E=
`pragma protect end_protected
