// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XYIvOl+vdwlQbwD2pVRPI7WS5BsZH8UCdLRdrZlgzsA9N7txqelwIRE43QkYlz8n
AVCF8SJOlJ3Z5vOxRHr6dL/nFezXrmv8qhpVQfR7Ip44wROKZa/CHpUZGfTh1lz6
igN9ou1C/i0tnkFjQL3NvpJpAjVAkVNfu+g3H5T8308=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 128304)
c8bIY36+bV6YuREOJJ0jglx4J/jMJYKI2LzzcwCO0q+HKhTNPWR26ZyXUzIVr9q2
xjX9PJKZDwz8aCPYUxAf4hQ2mI5gYhyhmrm4PtuWWYmAgXUfCg+Yp2WeU2y8pjmx
PdC4q1V8aV8SbusUVXPjfIfgUTWk8O1AMJrwuJLa66O2EpH2M2wo/36UDCdOfD/x
gpYMGjZx3DTBc9fjNESIUHP6zMB7XxUB3g/uBYn8lB8XEy2FDQklsnngQl/emaAA
8oGzeMIh0oGL3h28xEmzF5SZt9sU7YQ4ME0+WrULccvdbcqW97P4IAo6m7WVXX7D
DRwmZHtZFGsoncGRnCi/qfq7VLfAd2CMbgB2G3p5p1xfkb0OLjtZlO0R930jAgJ/
PtTMbgSX132gYKdl5UF6hkDmWY5cpEiuaYXCchs+6ixc9RSJ3K05VIUDfQUl6ZBc
ZgJRjtv6aNLm833M9zzMVZ4DmdbTN7rjPCF+tyWzV+O661d59QviW9WQH3RB3ivX
/CDT3BilKHQ+rJu90PuHjwTF+o3iPXycJ9Mdd5SGebVy8bEQIPMIKIl8yQUJPjWs
0BESdZP0tNbSVxxYwwfpntSCnXyJrcfqmd5xMsX0pvSmaH8220CYtw7dopfdxF+D
Udl5ofDBr+NH0CSqhYo5VJzOTsniIuCGlp6Pv4Klhu+v5xSFYEbB2KqlyCpyg9vd
SOINiimVZ1LCdcX9ZpLozW3jFF5iW5BE0gQuDHxiMMiIo/SMdNaUTVdBhLGR+Lqr
Nk+Hnq+YluVqRNacJMTJa2WmjByErM5uTUAW7DiJefC72sSpsiCkXex/HDU+Jz/O
kRaThxQiaXZNpCrWSUN8jKJ26Ty+wLvVwFv6HcGkvY2E8kFnrnrHCjXAlMNHfqMW
taUh7xi7aunTAnjENvMCtdF75QT6Shuxbx24WawH4ZdxwaKR7Lj5Bo9sx0NFxxDn
BeF93N42J7ip8lSFQfDekLB9+hFH5b2w+pEQG3qDnaG0o2i2o88D3lqrK9sZHhY/
xa4H8TQbGRdnwXoUHYhjEO+Lvg8RtdbN0k0fCk2e9utBzBo/xZYelT3jd6syq5oD
WhpPeO/Re6hpBv80NKwpHt1fVQMlYYw3Xw60d/r61S7ZFCtaCwKsAgggODGZTlD6
BenMSrd8EfqCmrDEBZRUziWvVkl6ez4nOSkbvhyCqOfzwxMg1uyb8iZ050oORKcP
wkBuscyg464URwQCrqNe9ux7a+2ndEvdH/pOdslcx5BcBiwKsZ9NrrA9t3cvQRqT
jZvfsW8AaNzRQtipwqElEtClNG/gpoJy629ilB4RD3yGFtTwsnfm7ema5SPRLjP7
3qFTXTc6CAm9/CZ3nEqAIwlK9btSzmBiTcWh3MzP5n8Xo6iEtTbO/oIbgGd9Q3Wt
9Qic6yA6ZmvENcCRf6diIBJ/la8O5CaahFT/28ybv8jRObiluER7KO83ZaPJoilk
bLbQS+HETuepnr6TEyDoFEFDVuuJEXL9sALOaF0vpm8IVTrRE4npLskWnqyy4nYS
voqsaMCb8OBbSkMYns47hnUpUPzKL925XdMR2joA15ocylaN3/+1jV3uRDu5RLEi
GM5It9RqPurS35spuzMiaB1weE82sqthT7PyKnV1BLYJ5g9uF7mNXC5w0bd0KSlk
ZhBA/rmcYC5Yq6p06bS4IhwKDloWAetLhQFflvV2pehghkmTKeolwRKrC950HaMD
vcpEQhHb26/c1ra8gYptngIDR7xJprRg4QcUhctztoC3NtW8i2AuS+yW35bLm1mT
fGmSdirw9QNCXtpcqGBBRTSob4H3XwYC8sluT2LNZvY+PIxRyiUlD1+RRO+DLLMb
IrW9yPez+s1a2d0PgQtRAcmmcSCHK3YEk/AkQy9QrH3XjrUWR4Bq05E7gBi9L9jz
vy7bPHsIxuzdFrAbM4zrzP/Z8+shUAnNRc5rw6/b1mY8Z/FdfTMk36p9W+vem8yC
aQUT9dIDVaCKa9pPZilhE07JneqxtPsXOpdJtoAuMsuCC0WfHTwtdLKn051Xp21h
GJtCBwCeUVvZoPfH8LyDII6ahy3RTrTvJQUz1G8xrRkD7smqBTBM7tlwPCLxRC0P
ffJV6p7avYDb/6WEgVb/0UqFyiSz2vf2ImHb1uZh2h4mt36oSsTgc6iMy+DKb2Gp
dGvwxOKPgnFwxrULbuhsoaSSMuMa2+ZALDRPSD3+Hy+knpmFJqGHoHX34eh9glWg
utzyET6S7KmtwzR2Gg3O5sYjXVDzXFqP40fsXDxGtorT2Te3NCirzzti+eU4upr+
4HGIF41CykA/q7eZWdpEYjih+I+LeKQmEYFzKNJRrvD67o7R4rhB19sQHeSyWpfn
fKZIiebYgFlTUwcAIPJQI0QpTLlV16Q8M1mSaXB8ceCFPpeR1gxl84psLhvUq/o9
OiZXfL1naesptxnhmgXdZDgsY9bFySxxZIOWTPz/W/KmZuFJ8zKdAiQS2n7W1bPK
0xQ7WgycngJj+wMANWhRqth0BSSO45gBJP3pZ9fsidXU2Fl9Op7OsFRyyhd69Nsh
CrCI8qtWS+asSL8EkeC/vOwqOVHHnV6VjzWN9CD4QMJrYq/HSgl5kIcfdqn6ARYf
Y3hWCCu4dwbfdK2e8sDo78KDCRdXX7E8FPmkbpdJZ1EeUq5s0YC20oDQEChUbmLx
YiFv38RnQ1955tsPO7G9ZngAuMlKkG/aNRDLm+/Ng6zmXRwQZM9z5zJUdsZzbdw3
IJPHJ7dFlFCGNCXU+LNGJ+tsi/grokYSY56trNOWIR7rGrx+WsNEn0Gqw7Acrriq
/rVk/qsuhtdNjEgNI1PABHzennsUsp7ycF3CDL28MYZq6wNPkyXe877dwU93GfXH
MwbI3EwO4Myy5AunW5hX07JC1h/PgEfaRYZRernlEwzjW4jnE7ws6E4A3HY4D7AV
eISxtDvSj0e3k5LYhr3/aB/+iinMASvdHwxyQLZ8WrxTZZnU348ZnLfK7pviFUYA
10SRJ66ER7rfpIUFjPm9KMiKXbNYUL2+50vKqAmOCrKWIg5lWWPyKIGU0faQ83Wb
lIsJwHMH2d+RhXQuBTc9E8Wx1tVVipD49esb0RNJGskhJj21sBL5upxXu91y9FL3
41CBc4ELQNBw0RPtFs/a9LbYF/ZBLB+WmzRlil54gumdhdl2yE3Ug9OTycAnp+5M
QQ7GxPy4iGIeQxxCz0pt8vQL1ORn58MlAJxZcOD0K2/yahWRk2T5atH4soAV0qzg
85FGrmczBn/6evkhA+ZEbWVpGJ0HXptwtBUgrnF5FQ4k14yO9hhT3hvS9nGs9rkH
pY+JlThedZSkPjRYqIpcGZNpmDs84PtFvvOFVy11+3/Yv8ZHiuZjQ6a7ucwtyUwv
QSxn8D3uqXzzkuimjsV+5gBFvlVwSWUjH749f72+Mffi/Q8QJzbbm0EhGv5rF7QZ
ySR43sHYtEggw8lbWHGotl5OfmNMUhrem1xoXn9CSpMbVhsUsU+0LfhSmYWmM4VK
JtxluM+YGBbZcjnf3OEx8rl+onq1MUNs2WWQSPgF5FbcbKDLwng2kwf4TJfndG1x
PCDwzbkWwn74flzqVbtUzp3npzDLeuH5B9tZfYZEXVht5nKxGEdNGc85mHOGlNZ+
pwxNwCav8wdl09zlwy6TIevEixhmUXwqH8y5/YZBxPDBeRfaeL9hi9adxjYYuJGY
URmbXY5VOD5ORZYKe8Ua620r4JFM7Kw5Fok1I1IphuGj1TM8AvZ413Rl/P9+TBZs
sdwRMTo2r0UFGxThLwoPlcmow1gDkjnQm+yE7RtKeXImaZjtsEb0JdtRCv7gAlAE
7Hgb7ypk3nQjwlvIJ+iJsDIByt7K+32ZV6QvliC4uyFNNo4nG55BtQ9Duye9jXYw
6z3OUcADm4OisLAQVNjIgr3ZSxuc+f2DLF2Gadk5yQ1Wh5qzcGLfckCD6qzgNfkZ
mc0YJLLafO68yjcucsZOhpdFTeluWyB7+6+oHu/AWvRv4BJFmASmBTIK4ufy6QOI
RE4YojJnewPZXmoZCtoGdI2F3bH1KJBqp7hMuyE3soq/ST7JLDA+beBnYDsUUEZO
yDHKeF0mIcYiobppDZZcdREyFWccq07Ji/1LI6FHgM+YmXFxLx4cWtwg+ARwAcqm
NsyasGbnFZMX3uk9FVR/eCtIP5l4mNnQlUCwj3lsNLooCs4RVh87vFlXTpsIojCZ
/AWwcmsI3VJdEluHPjyDuZn3VtuMrlCFqv89zVvrqMM9CII6U7MTIK38adRZgaUW
TA9Y/pWKwwFHPfcaFA5wUuPSZ1YVe1XhL75BeP2jLnDqcScMB82SekyrnX0D3Pcg
pPpEvMrDU1JzXEXqd5jm4aB7QBnRMajMG23dcwDqbn1mlZ01jAofO/PX1ueKCymF
h+9XuYl3LxAO4J1JonObJwFxswaXxaMF+irFfYlGDY/D+3Y21EdfsdZuKS5NOefB
JVibp5SZ6TkEv4M0eFY53cs++EWLZ/t4yW09f6YKnh/O7UrFUij5n36A3U/aYyJF
RfCVk05sf8X7+ltD/9Gx54UjrcLrrJv8cLor12+x+Ady/kEa4DjnmUkYBvIEwlz1
AK2tRI3Au/RUjgEX8nZzvN9CiUPwW29Diztej0krafl+gb+EVSIlbIw2TbmhYItp
W5wz2ZjdGfHh5ZXyqFgEQ3CVMcTzQt4jlyBTO6axnDp5vOXfeXB+RcyMuAaLaC7k
mvgoyEaqtQL9Weks4r/h2wJVeRE3vTl3fpd3jbJ45V/Hk0tM0fT39QrI3Np8xGzJ
D7z0FlQ//4X09HXcUM5+Jw1f83uX9ObpPrkbBHGhANO3018DCCVe2+4kXzZ1VdSf
b3MJrFWxYkE7Or0z0drAfAV1slj47dqLTPF7fn/YhoYaBt7pBiuFFlBL1z2mJUO3
UGKpZlAOLFYdT51kZcvLgq7EwmqP7IZg4LiMWEVABkzonjORprPqF/dP9RmT3kAs
Q/Lq5EeRJOHk/UFN/NRQEUH5G+zwPeHtkNDvBLgo7jKsqbJZUCwCpzmdoGTFtN/3
IIzvye+WeJLhKzfK1jm/j5SEKXeiA+SDxNtMgiWQ8Rj94KIT/Gk5kvEcgDIXRBnq
Pw4kknIIb45+XHEnf0O1P4B08h83wqVKA4DwoIbuG7Vmm7MOJua2fK1NJKFi1tEq
dRDeg6Q2+WYwMirhMarA2BOxseHOi7ekarp13XMBRWcI8kf6+OkEveLPfZh143Lm
Qv3MrjbYJ+m4RgOwvQ/OQC+h/iqobqePzn9sbEocLyQLvNdNS8fbyvwunw0v9VCM
7aAavxfA6qN/rp3qegaCr9YS/2cV8De4rZF+qPTYci27pMdbczFGZQw8ayhUAoNu
vOQ1WZV3fy3L5MumtxBYTTxHMp28IStfDo3mmo0TEYIGzZkhsVM0lD5oeXV9kGIb
ilDF5FjQTl0hvdhccKvAUNu0jgO6toZwXP2IWdCpx+G+Fbmyaz/j5fyRoIPbOjvQ
Y620Wz7E8Du0+Gq+CBRJWIKKJofkNNDafYfEeCQyvJ3NihW1MjSXbrnW+lCK7eEf
ndkl/cXzgTR+LwVV2FSFzpkU0PR4a69U+yc0slpc6x2sNex+pnOGvTO3wpv2RUWK
lkhM+vVVnTWWiax8mZv1+kAcmO/hDuQkZyp7cgwAq/YyW5CNjryHf+opr/N42KMK
/OSJLL+yqbQZKcJUobU4ht0BqwMGzEDiezDNOfmofeA/zEznVxF7PdWZFPzzCS+i
iRo7f9svzx+MLfKRyclr3hXuOsOpoqCEjjs+Nwng0q0USdEvKM9OZk1Z/Y6dGnO/
d/r9MFSMJJzudTtfvI8648lrM/UlN6o2bdFaYONf5BtQtto5uaKTxKc5J62iwCyP
qH1bSxjryjERZsVcsjiVFqgTnENyV/AdXHsxCDuiPrDs3XqyZYGIhxFeacZNZXCY
QvksHMIUs28LMq1p4oEDMMFaYQ3Joosej2I1ga0HWIWDa80Z9oh8ILT/fw6S7ZnC
N5Kq2pTxreWrr3yC1R3KUnpDJzjjmgpfOMQIhrtCYdbwGnz86beaKX74pTzxDxe/
4V4vm4YdBYE2HL0OWBh4BOl4cjYjn9PhMT+FJj6SyJnBNcCQ+7vJ8LiBTxhou2rb
GaJMSkmBiqrUtmzaIN1lj9d6xwMxwSAw1mvmJxMN7Na/VXnlRPQO4AGleu0F3K2T
dLiLx+jxtvflc5r1+/maYa51HZptDgcN6TYqsmk0+aQ8NUGDAnMMJ1/KeK40A6Zt
le+UJvfM4vy3/92lnu8UQcU8Os5IqpsiJcRKBvdcFNdPMT/0LQ4uQoO3qm9Hpp76
LnRPBRiyZGsG7+aH4TQHiTEld2lR0ntQopIqgv6Wx/1iw2Ib3BqTV9eiJ6XM2yph
VJ9zAXnA9Ric6RCzGUbdYt5Z+lpzPxnZBibq+Vcjgs/Ma5conDKLhVPEIYcnkmcC
5Fy9r/BzgO4vKV7n53mz2wBScin9MWnmGjF88MR319T+EIE2Q+SWDw/MoU9IMNw4
pTC30khmLIfFNYFyUqAxfkxwZgynmotnhjgMXHSpphuGCsMa9yq7tART2MOaOH1m
ebnLRtKbhda9IYLQlbS1l9S/DAkGpnaCQyd0lVr1rUqWYwcX7OGgOIedpVVVQ2Zh
qV/yei/AoaJ0YjNAFdjKiZNuJ27J3ZE7ze5fbWni08GTW+Jye3eywORM1VsvCT7/
vZnyH46hajFYvlqV769e1c81ilOW90KV15TJLSGYg41kY++SHhzVnZA2cw7nABaO
6oyKTp8Xb4ZBGPsVN1/R2piWcAzuaBU8asoDvmemn4ErzKZbjqn7SQrz/o4E6jk4
BS59Ryr0c2M74K9kqF9q8sKSIryn6pEKdoR4EDVY06lPzdWFXt0K5Al/ccXgpjom
xyBVdQHQFMQ3vL+Tk3QYjQv+7OCoYfMmVh32DdsTam7DzL4EN8W3B6smZRxP8Agl
uFpKFDGrJ/JKtVtd1Ciab2LcoRjsP64d9yV4osQ58QoNJZH1l/lpmYC13RyBusCD
LgOhzO7zacSULjo4/zcEcBFM/pdtCCnfd+8J2xFmpNYztW44U3pn8ZkHdfKrSMUh
+Y40DRtTYorMrLOpQPrhL9rJQw9x3CDYL1m0IZ9pQfnVkZhqgMJB6+ur36Eu7ynP
MoOQR7p6AA1/0ip9A8lgp4ayCuJ9V7yhF4ZpTHn9aPRaJtY6LWJUH9PzyaSDAc4x
GNr4lDLThMQUNqNml9EkPyuWI26EIOlCr3iDgeP6bIh/SzC9mTohby9BxePw9f/t
ani9yukYUzd8OBIwQJYFAcw+Q3hXwDZM/98iHV/daQZrYjtCKV+jbIVrsijQxjiD
HNx+LxC/zbcokAHY64CExn4s3pNKeOeqsjze3UsxWCgFWeMoEmDumk66cGliSNEg
4N/Z+Udo47apukXqKx+d1NGFDDjZSxCrwvxfzt7Aq83nWAa0TFd6w+bIAbJANfIS
Xg+XSxaviKYXYnq83HF2qIVr01pCXlPWysFej4dTaSYJncUN9VT3KFD1Tz2cE2YA
wdUUVyo5W4tatAzM4MOYlNXg9z+/LzvnGwwtNXB0yk42YWOUmHtW/p2+EpfqpA4x
bcoTAZBZ3rK2/VwSOQwJt85Tf9lNRIukhQ0KIWK+1yh5sfjtczSFpgesBXoAeRwS
Iy5pRH1PUQ+dZfqTCsmDdYlYyrjfqDjdG2+KN8FqyDNa0gkZK42AZ6NNSN9283LQ
KOmtAzdje8YxINIAotrcpjzlVTgaWrD01/LBjxqTRGb5BpB/ueGrmGr8bP7JSO2V
iCEiNsexsd0Rn9x7fnQFgQBIPCgS61LQ4cucFcWFxNsBCdwn0yWRaFVnWuVG++jn
BCo9U+fVSGYIIbk221s2FlKYDitTIrhQth68tEaMd3RfKAjBGUGPMBO/bgp05Th0
0mqcNs+F47ihUWXxctLqOIlJGy2MYYzm6R4KoBxFj0xezg0Cnk7I4IeQ2Ch8xuvm
INiNWLUbBzdcvGaDIOvrCWe+GfA0YnKbbrNeERCzRGbh2VQ8lWrL/bguGe4xVRc1
3kNerqckJlTR4red8S7b37QScup32Xz3t+ZdjpglRG4IxDFvMl0gQ6xwlM8JC6iC
QvVVKczVOtm8HdHg0cTCHqUi/9XMEbqJu0gK6aIImsAmOBm944v7CQcQxQ8MgUC1
/PnFlWHzyAQTKktAx9iROoDcFKZ9kQzWBhSaKSxWiQhzxiZK7B5mScwhxFPpmg2A
UnfwZo+FNuyNeIBgTNToctiCZlTgbOzMUR6DjaB5NB0bQK7pBDvRcLyVr44mrODj
ugniio8idten5R10p2TEHCfqWgqfx1kZCU55b0cB/acFEshc7CgzQQMBnEXH+0j8
yEBAZlCyDkpM/7u6284dsmg5TgfOy6mLrzF7KT8DOHzLqs2z9LNKgHAuvLopeahU
IhKCOREeHWFSj/cbIfzyZR3bika3aoB0jB3fi9kfqftJg2WzJ7NqKBoKMlBtBimq
6k+4LLAJZFykqYf5STrLDmphkdUrH7YBTpqKo597CdeMrEHw7MaptWIwI2IN2Dyh
qIyC6AQ2MkENXvGdU4kIOSpqN587bTnLhX8gIpD5tLKZWQ18jZHczXoX55+ehiUz
OzyMizWpzjxEVt89qvuzMqRo++zWqZENzDnxaZ+08rYKkHDQ96xR+DsA4h7hLKck
DfjbwIKMHCsKpDlgGTr39zxcACwX7I9HSTU/AVEvD4Y6y3iNn7/BhjLLl19ncfi9
G8my6FkEtU1jmGGAaPlzsk/cjrNK8sKyvgTClaVvUf8vMwdgGT4Awch2CjXu/K6K
HKPJ7SEjjOhx7agCGq8CQ72DF1ybDq1eA5VIlkWeLQOPAxJwIA4yIE2aJZ9a5nMj
lXzPYKiLIGobsApCN94KQWlDtDPInKRtNTh1pUFWeN9Yp+PDIbIgYI/K/Q5x8dJL
2z4XJeCDXD3PFwNC7s5zJBkol7fQO6aXJJZBkBDef89O+N4AnfYjMPLxNBQJVjkS
/pxHm2oW23yOfCv9qVchYL9OP8O79KhtxKQyR+p3cu7G8r+CvI6++Khaa39ewKY0
z1XVZdrl//QH0E+VCm2RrFIOgg+wwPiAVflGEXdz156EJcgOj8BDlsmp2H7d5lGJ
6smMN87iy0QrX1S8Oywjl2+D2N6PqX3VeUWsIfT7NhYx0/AJBhXjC0A5IO6znI9S
dq7U7q1obY8yupVYfS6iQ7+lsHaXnoEriSuu8ZjwSQnBAKC9VnM53SwwllitwRKG
g3jcaC/IHhrspKAosnPkT4hiKXPH08Saec0YPR8vDtEbnGfs9Altq+YoZUVxbdfe
ru+SJ6O2Qa2N7QvkNctTfMd+K95cJ7oky0pCypyTllq9afv6mF9caB9DNSxQv4t5
sGDEvFj0eX1ntyajFH+J532lWDpjPMM6GbT6jzn6qhmKIWcT4u6yxBANoXGmsqF6
UZcL7KjQv3Q0o6EVfaXt6uSxH51mHRTu1+uVyEDs0m1UMynDUHY8M73Vs5xip1zY
tuePaKHvUjjO6ovGih/JnMVCzwzKrsyf2TYhEhf5Fv/WzK8EQ8TGVxFdgh+6+tPi
1IMwwCSWcKeaj41neuGviF5r/fCLThUg2yV/wHQ+rjbkcpsLJYshIG3Fh4rKpKmm
VgIZE/Y/vN35RcK7NOT0QJUr1Far4zCXVJV8GPlfL8ouIAiSy75M5bVARjyfp2HD
+3BShvpQZ8nMEWlMO65RFVsIN89SOSGh6g9Qx8ood0mh7XkUhdzpwg7kTWOityEG
zBO0vbZu/PH/VCImw8NSMwUJPsXIwsHwqX++9rWkkSz8SVbs6zwcXW6QnOMFJn9a
Vk3UWtVQGSB6/5ZukNuzcbQ+RbIWk73nY4J2UNT+XR2TGitlLkSs+IgEqUsr/6XN
PrzEO+tTcrh0FhtrfudnAbjtxQmy8OEktEvQ9zo3OS27xz/FFI75oUD0rHvNNK7Y
wgYUzkC3I4WFYRmvqYFmhLujwY/DYAKEJBh53QglDfvAiFfztOWohv2U0vo64qkQ
Eb3GlgZHhISC1zDSdIAGesubfFNVb7sXGrx4hSOVoAUmTJwbe9W36UKktZSS4nGD
hvdMpE5Vj+CCkkq+/CAtTkKN3m7Hx4+L7R4PBlR/NUDUzzqk8AFQvyTa4Ob/DHNX
kJmZ7ACA+3RS5WPCHIkGI90L2Jrf+D49OIxfkAeOsoB2vfw61rmCS/A+jcWfWeQ/
l2mhu190q5DDYqVI9sMt2CW6WuXXKLMSmYNlqhrYdLg9lZ35hXGdKlh1zYeTX5yu
89C93Vr4G6e6BifWl026XA7vuJhxteyXuqCuIwY66TZqKkPsrJiwmm6KMn0hvGJR
7nuqON6BsMoNHOrEztnztcqL3Lzu5yS0emy/Xl0hCff+ScZZ92tjNwuoOy5qrF9U
tLNJn6RGeUZLVv6XvYH2M+8FcWO0PN4Xgg/osTxTHICuTArKDb7J929tx7A0N/+l
8/DIz/sbUZpGLE/23xOtqiF8xtzjPsehGTqCj8chAA1NBHcuauibDqNwHA4Un4AG
0TbcaDjansH35b3Q76LRhZYN21gGDVvy0u89v1CyGLJMQGyqVPL7SkXWhE2g8plF
PqW8Ym6wdrCuOJLAJsrWELedYNhgoTwEYZ7K2R9F8K69Ca+U+IIDBJp7jv3WgH0O
culWfMJiqYCG3Hmohy8amwBQRAdg+SE3uzVySev0iYn1B4K63R/ICL8ydF7v/sTV
0s26XM61HgCLC11ziQM5IcCSd7Qld4t5qAvRNwhJ26eEfmHgTCftXEYqTqUtibKq
xh4gm6HTeoZaVXVb/j91Iy5xobPECukzCogTzkhJMriHj8kw9mJ4QdkzLNBcHDnO
nTvLILdqhTauCZQVGmd14LJFRpAQtWTQ2ByZw+gKrycHOgnYUrHcvE3U/Ek+a2A7
fXZGKyHy5I56B8Mh3if2jQQbrEVnScGkUvJ6gwTmkC0UygS+yXeUnVwmB0nXyqpR
YGt3sLuyx0MjpcdAUWE01iuFqCiN7F7F3AHD4ynMdjR+o8LnEAg1vrMH5Ex+8hp3
dnCXtkEpjrWfB1lTdd/rsRAOp2CI8oTLiqFPMtSP3841+nE7Od/RFkUfLDlSOzKM
+QeOF7o06PyQqKYcJ+jqW2O1gdOCwgrVfmioT1AlAtdEEb03yAPf0c27Mu/KiVAQ
yHZk5lZjtPakxex57uMJpTzBMBZA2gL0RdB8I+lJipGUzBUDNLB24s9kQGUyl8y7
dCb5v0HXX0TQm5iqSoEujJbciNZWyiOvH8DxBNJLY7ejxiYIq88wSrXxJ/gtK5TN
VJF6ejYLlM6Xti1f8dKxzQkGqIOWluay8flsd/H1Tq0X8xFX2No8xyD8x6ZIZ2vU
kZAM36DU7qBd+RMATuKze3IgH4CgHqV1Y3ZvxN8aPbJqOnIJOYd35DsfjlW5Wf+t
wz1PmMUmSYNYtOUS2Ez5psNXzoAaOLhEF6wgt36mR30CHt8JIQgD0DoTzc6LOrY4
KghtdExojK8n/EG/MQRdLbrjD7m1vVrC7MsA2U0By8D5KFyNwFStjZuzhU6knbhV
9jfx8eWXn48opy4odVlnvChvMATiJGK+vF8+nQCXqBANawa7LEwEzkV9cX6qcNnL
hY8KiXJ6sY8y6SL7S1sJDBHHq1vVjUG2xzYmIVwR/R2J8MFQx5wf678TMHzZQxXc
xP3axa5b5LZUyV6lzkz5v6os1Xiw84xFTS5sD49kKGboIOg0LMQvvOJa/ijxzO5g
O60yp9r1ve/NDmBYSbg7PCTxicov8ZsVBp3kCEZha053y+w54skKOOpiXThPk+0r
HIF0LwnTJPTgAM6s9AmC/b10gqMLpni/0+u9p3i6My8my0M82DVp1yBnGsYtCPCU
wEvRaHyY+PAhJ0r1WGWlm7cybd010UyFElTtuyt+3Ymp6/2/RTM559zYBFvAYu8t
cDPThaGqz09tlgaZhOUOaE/H807ldQ+vjZNHAzWsHPDPKrHRx335P03PG9I5BgYV
uFm0qoT8X5TgA2/zMswU/K/2bg8Ekzguao67OhSSA/tkiHrhh7xZ9+yTcnWq1631
FVTS7vRQQYT7fQeNE4ArAnrLnsMCPKRy7ndoD7QsyjSqgrq1F+uUlB6rsKqiADle
3sD3D5SHBJv2qfsXRuajjXqcVitAno+z+LwytlhfT8Q1gslIdhJyV/gcAItHuUtP
UmopYkpO8tMmushnKq8sYhkr/+zLp+ocsD/9TH4iG7lfzauECSVF61mTh4V7FOs9
Xx4hGvvY+X9YQGQ0Lnnr3w6sfEEV+g9Z8ptZ83tjPTzlU6/rhZJcCYnVvVxLfGaw
RcSXolZezS42hYQwd6lUijX/9LJLuCOUpkpl+RqEXRIPhkjDfAe25WQgKF1HxEhv
R6rMXPsVOne61NNv1YrSg6fKkVRH0P+NbkyBh9St2Z/PmAuBL6zDvHvn9KyQobuR
zx8OIkqdZkzaD7/GwBkviTV6BCqVtSYgdini2ZAW/2nbIZ7QMQYsWshGSsr1uz6m
q4Q0XdHB15Mpb7cWd+/wIAuX7VL2wHDpde6/ikeZqOhOCeke6sMsYA5fMfDW5aPE
BfbKJ9G6HNKiWNe4luNi5oZEMjJPE2pRN3UhSSDJbKxCaPsTZ0L98I/lPVns/62A
Ad7EzuH46mY+atfwl6mm5AULSGMu4c4+35bSIyUu7LFXnOBXx5+0LJV8kjfIp/Mb
BZIlKwWEkMtI0F2BzxEh3JzFkfs89xaGetUw7fNSmFcPBlL5zYXvLbH0ckRex78j
QlQalUK6U33xDU9YxVviQtd/zX/z/v6PbF7kqpceohqGrul7vdF/uiy46uR0gPnv
A4DzljsOaie+AwhzjUbe4RYxsBl1bw6ERWfGbvhmksgE7zp/rycRtrlUe54vaiZ+
LvHLssgjISx302sbzvUGQFGS6odfTTx2p86aDEUJjcBUd0ARojGSWml/ckSNxFWN
U+gHuYVSLFaJqCBf2tMsU2WTJtrgcAWscaTbkPVEdspFYO0TFX2TB9FdvRbrbrt9
qoJafl0c8PEnqTwPbEibAI+RNQ8RL3XBbWdGfm0fmt+og+805H7UBh6683MZIMm7
ZClB5WLk4RUPFnBIicJcGlNDLV4oCitPO0lvLopMyCzGkLEWQTxI+GVRZ/Io0CA9
/QoXwbgEnGAdNhd/xxi0usdrpYNEuBAR1aGsqQsX5Rp1jNhLekBSbFhRd7RdGeII
IVe+2IYiomhrXDTklD+gTyLIBEVjwWAQtypiT/J/cwuNDM8eadqMRG1bLhTkOn9T
+WQznXILvI56R0uWtjt2cr6PHncx4FRsB0gi65kzL7VRyrbwysDetT8h00Zg09C3
MRwaydf1JzN7xtcSOgsE3yUefsh9CL0dikuDP6HLY7cxWg2QpSdM2kp23M7L9/C7
dbTyPc0WRadl9uUvXqa1lWrNQKcgzHdhQu6deQRiJXyqHElAy77EhRBPC1RX35Oa
pyUYrcDuKxCwUBMSch1b4dp7OAZtJAau1ZeIyjkcmqpamVFgDY5Y76KGpaqaV/8I
9NZfFegI9Zrz26MbbedXE8cErodn98pa23bqclaRcjHSMF/C1dIah1x8x/6Ot+WL
+mvnoGCyk6d65eyTx2bjleQU717hSIqP3RG7T/ucsHU+QUPYiBABUbtZaqEG+0YY
GG/Yh9KjklEirtULZLK8HM27ItJvJXkYuR8ItUR1/2B8vIjAogsGwWk4znlecCya
MG9U4Go8BbutbKwlbMbuAi8W0EnTbWNiIJZmpYaa+NXdTu7w3bb+R7tXJtUc6tup
XXECz/xeUTqFONA+kIQWnj/CSkVhOH8RD7QctYXEDcWFv8y/ylCfVcge0Xbz/zj7
tt3MHDJMg7P1BlbOJ8QfUoFde2jFivusoGs3owB/ZzEGPugMwkX8GxxRtPS+oD5x
T3k672GWwdoBoLOkJM29Jqix4BlwsJbPPMCGHIGH54IDBoNM5FyMX1Wci8v2hSBx
tbFmrVYKuszTHyL/cCHY9nDBAJLoz2kFWXdvqRzN52FzqIVBq6PKY2VaEwWiixvV
XCGHsgykOiCm7T+d09VAwZMxEubtPIJsf4uFrfbDbK9UR1nNLZ1sTt/FS3htRkz8
NxmVk0mT22lQEkzfe23DQbhq9GHTAzGi5XXd+jxF7gVrWnBgm2JWBvKUF5t1/J57
XNZzy//Sd4d5bk9yMl+LdyXeR6SvFWJ0B5vhOIZtoHYA1+b6P5tnPxUT+rtQoO3k
sseaXqwTK8RIrprSAvn2mKhRJEUekf2mB76+bf4v74eqDvjcjDn5mmWSQiH0jgnw
fxxuyCIh5rNQsRmHuIdZTbVR6sIb173k8DO6Bf4h7n8jIl0iWzfC9RVCnzpKENoD
gMHH6pI+6sSS7gfQ/2FW52nMSpXuFGREak6WZzF9asxyZklH1maYAi/Tmz5oHvJG
fNHE+tFVNxGJzm6dw4JtnpjJmX/7yaBTaVGcALfidMCMNWbrpHd3tIBrBAFcRgla
VijmoX9wJDRPFMRIsbC3EdUM4jjeOOrQCSl7l9PFntH5Dsy1XRKSPGHo+kZc8m+/
xVRYNWGIYocta/1rXKLf4BM08nn4MVuJcgZLEwCY+MUXzQacfdFkOohmTlULFVex
EwunEOhP7JenxSmFps6x+W6dsEI+oANmNHxHEAVStIDNnzZ4WShxffiaB2KayeLT
pm8hoyZnHqUl9RIFYp2w68qqLkiVB3GpDUQ2YiQfwxi3DemgfuaELqVsZY2DyUMT
0c4O5xvAXoqECnDaGO2qoddDSlP6SpyUbVTaUM4mEEVmwniGj3MmuSR1f/QCs3A8
bSV8wlw+DzmoFc3edgZ/+KeII7WJqpyE9OrzaiuAUWnLrqOZ5cAIONPUCstuBiW9
lRbs2MnzKa7fizID2z1wG9KMNS1Sw3mHHL19DeL/zkJdwTPla1U50oIECjSDFSQg
oT7PxXnkYHaEuq8PmoaRtADheSAOwC7LqDAoIVoiJkyojcLP86UyNtGdX0xeZk8K
HjH4y/Hf5KvJPkaUtnjB8a83G8FWSJM2nKKtrvO5UHctHi2K8yv9HuPRn3zmEw3o
iwfxU6gfCr1L8La+NnnBYOfFCi3uzYFF0nh0m2RZpnIvo6rItVk9oaffja/vg9Rf
VT5rdHJ5k1rTu3WvDirPOXksztQhvXLrpLpHrhJbK7v3NTH50YF8EA0ioIheP6rb
6eQGJBTvFR/BaZg3ixPgZ6ncMz3hMHwwfrcKdAEsNKyvAoMUe1oeawh+HglCTmCr
722FVl20VJ+TVGn8/Cjm0ftvE5AEiBRNR0DVtKnuZ1gt8vEO/z5A4uKwvR6iiXe8
9yUdcZY6mIZzpWHMbdAJjdnTgvrAuNbZmJaGsm/+PA1mmmrS0zOgFbROIa7sXG3j
twVIvQMjHITtSwK6wlaJWgmkwSLxS8tx3+rhX5hrGGCCRfeqDxMzVVnsHZYOAKYV
2ocHo5igU92aMRSXJ7uQeaACyd5+Ea2DUr0VmQ7mItG35XJw0CqwoXv+URPufvH0
Ae4l55flhx75k3fAXCT8q6Ck52f3f7eP9yXbHxYFyDwNdxydN6qeZBNaQ022NAtM
ajgLn1iHBQD+LsA8sJDDnvUDrWGXV+j3AcBpLB2ZeZ9FC4b3GvTs7FhYPLiI4VL2
7HG99c4NlGUwnrnzQKO/D/2bxNpnXozsMdWi/kIYxyWSg+T7aWe1V+u3wvRkH2NR
WhoiTPTcOYteCKwZ22xBzO5xnJTUKCxpCIRp9KiHcYH0z1IlzpnpU0ykgYWHJk0I
eSy3QtXwDuDf3TkIbL2yOSob4xBaCTrfa8qT36BFBDwPTIF0nvNClYcHtq1FUgwR
5dI2THAF/A5istL1mv5YdrrQF5YVCQ8Ci8zl1xDiHHIswJlSU0swa0ARFw+l3aVe
4cy7mNeefwn+6gQzVMfycwctGeHwWlh+18Bcpj4pZ7LBbliJ/C9WvSXerb/7GGqi
AQeBgA3Qn31qTEoY4M0CPf/E6azHLJh7FLlByjAultq7MG5v8xEB3n7MQAiS1gOl
m5q8jo8TwbgiePpauXghgpvqElOWSubpEK7D47KasHV+/pG59qKkS6//zCLq3kT1
rvNsSvKtvB8AsQYCDU0bxPY1kOijPttPZ3xQSM+nP4TE6qMa1kJlXPI/Jbos6NlC
pyJLGNGsPs7bh698TxvJCk3FiOr4Gj2UChtYHczU5yPuKBY2oDqBiYA2yPesyTpm
tnCvbPDb9pOFDhes7x5LVJzT6kIYKmHQLnhjFchBD0ivf7M/UoEEqeaN0SomMcoK
YL9QpPpM0IdjMupN8qsVYP79rJGfxT6LDtgJbFwKwUiC5z8noLK5W8qL1KHTHDGy
i2sUewRZj0nFa2GL3ho90ixeNiLnH+VM4J7xuKjaZ8BQ64+zwKfo6GbBgoSeA71g
6+OvRxkEnOfR0baEdFdwmAsW3f0CPFTBwolrQjDNcu1t8gcafNo3VHpzfHHmrTOj
3HkdZYB/0x3E1bzXPtHpJk9a5I4Ig7CHlOREj33wiwcLyMfD9JmbyKD6DA+yRTKv
yn5vMcGg28/reRfQISxvtOs2iLfwbEIjV97FKC22Nv4Qwou91uMVPp8X4Df3CcSl
YEk7QJ+t5EuEx5aNkDogB1AHrfcVkjOou6kbHxEkAxR+KeHrAjE12w6x5Ga1p9WD
poTgmMflMlQcsCFq3DY2kLWlrO29jeo0VlN/r99S7eodcYi1sxpw0NDm/nLm+rmC
Ht1q5+nmEIigwehhDeB51VUHYsBfjuYhRy4n8Mq2gHPamp874YXsHm0Fi1zbGc8K
LMRYJQeffI6Si8mvLVrWp7i8ggkYl661szZ3Ei/5e4x/kYljGBhLLt9/iInxMqBq
y0wykXCHgojuh8H735hhBvcv2tLMGwPVqtClCis1z0+DBX4W/f+TO0vsAgOoN/0X
E1f2R1Kvcjqfs03hccTGGfrF2DvmH3llPnMdYteFF0e4WTYz+KNT3wGX0mAW0k9l
DXJ65lCqla69qU+fj/OyotMqfEtXMlt1WPRgQKPD0zjZTGh9JROQCTiiEP+UTgbl
10bV82itz/40I8veZq0SqSG6uCNpuLS1HhGywBSPrsXl+3CjsPrSPquBIcz6rSSd
yWmNsf0vHa3+KHzdvWwVichODo5mLANbp5N3VyAKCqbsq4fRabsGmwfq70OJD1zM
Ejz8UyjH7Nu9AMt4Gi3zbXhhfa4Bb5fQwij7bVkYqoMnm84yVBl7FDf6jELhU7Te
rud9UppbdHRkuCIbxNWYM5zWNdoSTTy3CG/n96CFuw3KqOwbQmmAZciOMvTJ49Hz
Y6rBwpQc26KsQuquWyDyuaYt5ZQQEXzLQeMQ0zcAUvyQJ60KE75Y4xq5OoydG4/d
uP9w4TBLhGe1GUSw1VIt8iF1VMFdAd69DbsNY17Mmdt+Rax4Mg2CLpwaZeH4dvjy
40/OpwwL84CQhtWJA2ZOmL5kXLOKXdI3mnoLcs7yd5xsjYwOPxg6Ld3rF9hCNOZX
ljTs9gdUfAJWdhENArazgJ45FKTaYYSiREJ2cBU6c8KksbkAlO31aN7f8FjAPL+I
bc8FOK9QSp3JH/E6aCIvWWokboJiIPPb3zfbPi+YsFjnANlTjo6yDAzmd5Ytqb51
5/FHv9ovWuA8S8SslGGGsJIOVlzGj06a33JTIeO1dCzzG74w8w2u+huIlZQt5cvZ
A3hERclr5THz9Qi3wxO1NChqYBG9tImSARg4+3Wu0gOvVxHJqdWtNzM5h3PRXxTS
pEgULKI+uYxXmmdJyfVpViYVqWxZgZ+4YKSkRmUzka5i3qX8sKbhwBNmIIGGkdto
0GyedlN3ZrvUKMKNpCNyURMHOKnVmWGOXOQ2+mkhE99gaOpXHsX3oCYFivEwuiQ9
FNtkH+7Fh7Qg+5C14k7tjEhd9QpOWz8J31Qhq5ybqkXGZf5iXgaOUsHNkp7q06A5
HycAtqKFKLKdMTPMs/iNvmUpZCYIhvd5tRo9ghUx/X0lupSWfSVLIUZ2z/EbGdgp
w0fGPsXMudwM3r9fcnLWNQtEksF9jWQAXD8pb/BmIV9XWWqFg3Kw3jItA1qnAgIx
Pp8RPQJ/socffEy0igxJzluQUwGsEjC3+yymnri9zN3WHkeeJZR3rc/Pt/2IUH1M
5ES8HfjfII2HPxP8kquVHyY5vY0hmFhuL2kaATqPOfEcY9eEnwKSp/esCMu5j0iL
mT2fdHYyWA858vYAbdB+d6j/OEr1ayu714VAhiJyD4ZFF0llH4A1+6XXStnOmVVe
s8hMEEH1zFtrNUBibGr2RZ06Et191Gmzn6Xe1tp0/BPgrQim6jsMf4mvp+1uukxk
NldqEx7EpsjCkdx+d3CRkqX6Vv3tTY+O9EduE40Qy4iKNzYuA3BixjrXdTrX/5Jg
sOdP/7cobVsiII+2sscGYmEJLaUj2SUsVHO++DW9tPJ7P/cEApSNWw7FFK63OBhB
fwql/IdJBOWy+jqR54BytpFUh3OhqpQ15W9Z3ETvbDXJ1Wg4obHARnB+AqWn7Uis
tx17K6K4mdtFSOr3c92aewal7tGKV0n5zSdW8kprQ/egjpzFYBpWp13kyIapyqpj
PeGKea1qFF89gPM4naVvVEq4zeRarnE9JrA8YjjLx15vjtvg4MKu6h729RyCDsiH
39z+s/FdDXp9pNJ37NXpmELMFQy2tJSn9pf0q2SN52DRNneaUBfxRaCvladdHbc+
LY2OuOjmOthtdF2g7LJDSxVkEig+wSoo7SBBi3aKrP8sibaWs+SK5zoaS4JKmcTc
PrWWluGJGpGh93MX6K6S0VvS/b6s83aLil0Lp2/bTarGy2l8PJ+i4CJrJFSRIRKH
uKXoIPg0rHgGphkLdDX05CkMLg7Xz047cXfbR53DAOasct7YEubChUHJprbvnvk3
9a1PmNaYGheiQLXhdM0QAD2XlaG9BHxRukalfjXtJRpsj4FECQABeTPrM+fBon7d
Pmvz8tah8COwVFL5Qh39ynxDNbc1tsP7GmVmM8VmRulXs9sauDD6Datm6pHElPo0
eEm9qyYt7QSt/Xq4kMS4K99Rv9XoWfuapHgmfZKe67FNbViJftpjQozEkqvbUSch
Aa4LbzTrhQWUmV3HDY6Wz5QMrvZXbQHKgWnhqpQmx3qCi06gWnTJ5Zh6oHWBwiUY
nbYjDKK0wjiEtdbQdP9fkth4DFi2ajeoCqgUEP8Fw3yWLN8nEbs6pF19FffTF+jM
Cr1sDaqMQqa7C1afGPy+Ti6IH1pCQvbuwLZzwO+iTWf19uWSObEZyDbqwDlR5EAS
x12M7YNd9vcZZX3KY/P8NA7wmOzf8Yc8owz6A1cITS3pzgvR5usMwL+DCw3yufjT
bthqusXEh5h4eAaYiJWM5qRvHtp0fX6nitd+UvSm/qrKTEHu85oeMNns4bwDs+6o
mm9Ply8xGWpcUUea2v3Ioe02aKwguIDhI4ofU+tF3IDPdmugcX4zQR/bv5vZLOtc
erVSGp/urmex8o3VPN4IMQ8mrmQHNVVbm/YwGVf+Me1C+Nr1ThNAII0Ep5GN18Mz
FvYP30nJ4ixOkQwM7qxfoU9FBd4E0IBtDcO0OPtV6jib7FT1SdK23lGYjKYnGCmW
BhXWXrfzlObr4IOcHr2od58lmBxH/8MgcbpFu+XLQfsDIFJxGXNkDDKdo22SzX3x
N5lKWa3UQRGJo9vQ30Fr6vbZuOROxRMHh9qkRWvS39Z5h2cAusyjQ2UY2Twx3jiM
Lg9Q61yspcBp8tGQX9rXshMLTFMTGVvp4H8egDnoknS7Yot9TYhr4nJYVBhwzeH6
AqlA37TFk2/mspEZJe7oYAuQEHfrIm/0D/WuXmFToeyzSL/gqxU6w0J9cb8W060j
pKJdWGFI0UWUcICtDnAXLdk5xaWApJJZhpL8TCfV9iVUg7g6RpC6nVM9x5M1Fwu9
AAKrJLgsh71byMH9s8UE0mvcJuIDxlMreNPohMCAkYQWMEp0CwrOKJDII5xZhEPf
AJU3igTk6mDSxyFilDxyqAIrFvbqwx/gMyeR3Pn3ey7slyPrFos+zW4UzI6utdn2
7LlYV6RViDR8yRlvf+vM1TWwa0Br2avYvU9VG46pEElXgTbvn/+c1M9sckC/5W/f
rAZ2R241Zr5ZrILX+uTOXSpLBnQIwJ9xtRBOxNpfaTPsLdXXC7OcCTO2CECLHnso
a0m7qZ1Kv/wiMmtm2mcIK1cURtKMnx6nN1cfivtevFn3yhXq9y4mrO2s9p2odo+r
EQMm4b5fNbJgjHKZpSnCweXcz1XZZtaurxmkqZSOgmLx0hrUNPQLeWUz6ljW0KeT
fbSvh0RLGCCzgjGEKntbzdDOHgF9nwpS7hdQmvDie0CNVOk1/5VBRVXdXBoiWkzH
Be5mhKmw7sIOqeqvD0cspPeoVZRgngh2tYErvK/AODpq/pYi1JmnNcWwHnnYXiOP
8frjCQSa3Vj0AQ/roT8PcE5HoDeQJQ/em/9fqfurygfmqMNL5eQ3AOrIa9nQeNEj
6iXB3YfyACdW0+5DUwAg/DV9sCmBilukjpnI7EbD1mstDX7O/m3Ok6Q4RXAt2/fL
SMIpKUjsT2aTmVARIhIQNPCuPZsktM5RZ0Dxb07ltur2gSEHmQCGBJOdqh6PVrvY
GqyQ5lUPa75J1JsI3NxZPT3l6EczR161udqUybpfFF7hTGgNkBgaBNovIjs0BG1q
HmxNhw+Ox3HQ30x2tY11KIf4u+FvwG7hQNYL4HiR14yJ7N4EU8BioXxk/qrw9DU3
7a+T0NKn+XcsbgQLxm8mo+8nA/tuyd5kvniC5ysFHAnCKkVQClGEN+jYnxdIvPo+
i7Wa/EzRoF5YOtiyh2s+pRTpzYgN1x8vsJlAjnKl6mO/JARxTYwhNh5Tm8EOgdpF
1p8HHuoxkAiWLVz4xZlEj6IzWW0lkRDO2QyfET7t8Kn1m5cEdxarlIYcV1j1AcEr
FmQQSCCn7CjaGhMspeCTXSZhJIjskdTyWUsLCOQToNzpLAh04iCtWW6OSO9rd460
CToV3f5W+CKiCLcgZ6cafWqiicmVyys53Iq31F7+VeOSy1YUe0gbt3tx3V4DRQXn
gK5L7oqOobivderzJmdYQR5Gi7pm/QtiSj64+WgHEN1nD4QI2YhEHcOIsYVUtQQY
9Z6lSH5Tv4N4JgRQZc6jPST5wfAHjGW6B5uuzGfm1J3Ev9gV1HioQ205Yifnp64w
kygnYdxjEVERoOtuH0ETZFlxlU2zPpdHmplbvVPeLTdNVAGXzgom+HiHhC5kwiDZ
jxnBz0LqAqQs2u5/ITogV8Dgfd7oHBVRDbqxUc/UESUP2yv54gebe/9cVI9N7mec
qyyuSILUrnHSDy6LQwGMqgcnScWGGcbhvRrw04S1kMJ/wtz8mlvK9h3o7mnt8qQi
TXGdoyWKbntLAL/1m0DE+zGb+buafc44XkstL9o7cpbD/hMpguNo+AYwwpLFgs53
nO/wemIzjvYdNGTkgjx9w5R/Jtbg1LoQfjiAStP+1u2q5dUmYs8aJD3/aWDtX1zr
4h/KISx7vmazMcepx9AuQ0jZOoSuQ7w7pSk59OawSMiH5IWvIzbTRhKwlxrHoLPm
PYMWf4g08bf0Bb5B58ib2oFCy2+8v5Wj+YJV1rQ2xLAhNGQsf+/c9PTFJtBpVFJN
KAmRaw5XedOuqAlt/M3ZIUOPY9bSN/edy1yFXaJyqL2Hvm8kTT+i4XVG/0AhzqcW
lPOkf0CrIcaGPxdshQLqJJvYBfqu9/p4VM9u5MT8jX5p4dGTuv/zlBTsTolb5Luz
pJFM6RDDnaraR1VkFFQU1vvmawryMrNTQ+nu3kUkwl2OqxqFC1QZzThdFjROsn92
E+TdKNz0S0eUbr0DEGmNvRL4PuI4piz5wR5j0Z76R8BiSsXAE8LR8bTOlO9sZE4b
TKOQbGzaFHFChLWpz0eMxPE99VX0FAbv/b+u1PVgedNoqurapHK+51FInHkf644D
k8oG77lpDJBSNhFiHkkf2EeCqj5DH+hXiT73Csce5tCe6fLt7d1xsrk6GiQHtlZN
KyjcwcXbcxjuS/gd3ZYoypvpY7E3+ppemNkgH3Sgif+YuejNFOQLdy+pHwdK+oXf
dvrV4oQZaTvXCNBQHYNWFlmZfWG+gIhdSrmiw24Cdqlh43KsVvWefhr8K6YXCaMu
Fal2uGvCRtNAgkYKCGRtzXPMZPxc5GF6ODB4pLZa8qQ2modKTHpRzE2i6to9prdY
T82Ut83d0cOzF3pl2Qr4qEaHiD+gQQ2f/UlNdIKDrRLpJcD5gdWjKCy1x0ThdF/j
7PiEBs7py8d7/QfaQLISA8gnXoM+ujx8ZdGYZfoSCfbPUOk3d4YZL0cc2xici8ap
L1UTCTYc0CXKOcBPDWZYrMj0GOIANWdultH1cjPrtJCe3bZTGwdtuUWdNAiJwa3z
iEnkU/h0lvDShHv52d92h+TACmQC3bHRZnc4/czRA2C8c3DERY7BqOFT4VBGrTUt
BWz5U39VcnIPSrIQ6pYb4CupnFaRLrgj4J/uw+r+1Isl9rgOubTm9+K/V2NKYfoo
g58+582lVETGo63mED3bwmiL+Eb6+lpDOzHidImrbjb7jmi1d/4sheUsM1Y6v3Qh
wJHQhO6i6ZWLwoyox3dC1z/tFIF80i/8OgRbslEsLRnZSpnlfkZ4ZnXX3aUNxTfh
BFTkAc74DYNaKlnZFTYCZS8zfZFlJDc0604thp1Stda+r/91QXCzkJggTd7vmIZi
aJZgpFmBiQ9nD4uDYq/5qTgDYfs6qP6busETXJNbYbTOz4wSuF2llEn7eoY6H/at
9z6tYi1Gpc+NsdqE6r7Jsn+34MSGfNi/FKDXZcDkCwvsHzYfLjmeSE5+7TQfkC/8
SArhzzFBrMgZr10EEjXelpWZiT+7dqoQWHXtn6qbocZbpXoaD0ZDh/A9hPh8qHe/
EjAyp4lZZ3L4LB4t4zDQT0TCphvjaGOyUEaMqTDvltFFTReU7AnveZkHmiAZqzH8
t9QsDYe/MgRfOHOQbw0P0KgwwzyTPX1iScZoWOY/1jtNlt/nHsXil/YEWryCiA2O
2WNXD6wdX0azGWRHP3qY6mwCnKiWAT4rUzQWQwlr0hnMqp0YfS1kxaeTT8uH6Y9x
3FMnBqpXNBChnSg6AqUADI/kHma/EqpJa10MVdTl7pXezCub13n5EJVzYBrEaz8c
ucdEu/in60U8+LV0VQU1esykzHz7ojeRH6xIm8ZIBcrFvoWnaph92X5GZ3sIgl02
OkotMOcAfzqiQax0beEeml70BG0DS3Sjc2NKnrDg3aS0qabhge9FEtXNS1xjvAKj
YZI+gtQikHAPQ2SJds46nM/fU5z752LeiXIJjLSmrIsMoCn35WlMRavYmoZz1l4x
o1JBA+SqjER0WRNi8/Onu0XgskjtLFzremDLtMrReqy7XtlRYLabhOp0Waxh4iRN
V2FhSS1ipNEfmCZkVax0nUhQO490vfsnG5Fg4JcKR/TcOnNPUNlWqlyI2rqKPC0t
1+6cz5CaTuw3hysUC7jB+b3ictI6KbfDhs13dPLTXWXst19n1vQO94ZTOy8ttB2f
uIaUu1AxCgyMMuCkmG44GUdw+i6HX83ig3T9qIRSTQMgvXnhWvmW9MGDrzES8Etn
35gXje2J2PMy/CSpEezOTVLV5anhWcKdSPuv3upvNdein5bNvAwz5fp4wtabN9o7
hRT2Q9UGUap/5UGiyuujJkYjhIe9q/ZLgdKDsNdj+9QAZcXnW4HAvFY7JbkjLjEA
xZYPX/u5G9f6PfRhlG5D2yaRXLOl4dtnw0Wdx1kF0vHhW1+gZOKLGQmCclRCT2BK
kkDrCcwTnpHa5YAGCyr4idKgyOhIeFMSqS+p2liGoG+PSu0UiNT7Dv2e9m8/+4EV
tDI49cSlHvLLEbdThc5S16baDvEHr7ftLbYcRRvvbrkNNa3otP0C5XNFM7w1/PL/
Ae2/5xnnRTCdhMAZlgTOJvqhsmdjDdvfESYaqQqxEzexgbR2LsQNp2cEHUGLR4nR
efeyUpc73E8ROjYcyZw0FraWd3+spei9g3m7GQ+vNM1xT2dCod7uphEgght4ahiU
4IkxySsmlsu007RhqOOAHZ2i8DWLrEkY0o9Gycees9zsINwl3nu/QnyRRoa+/KzI
Av+KoCd6yndNt3BAqnw1+uV3WNj9PUM+BedZye42NbK6ovVE1Hp2W2859+YZu6+l
E5hpJ9GxDyCozbUUoaWHexAbTaOKioonHjgyUxKqXjC3S5IheFzlKWT49ABILU83
6Qn+01sZmvDYYrGApcejEPp4B77ZXm+sJWmFqY4y8FFeNQQQjrLHH8fpneCt9xFb
Eu3QNfNxnQVizVM4fODCi3he4R9lNcd8tr1lCrVRvcOymq/6RXe8a4xdWV1fz3Jz
Er0eY8kEcf1c8sLfTEJO7YhN/NmKpjRw9/RMoKA2tx+geXmLvcSEoamGhvxH8Du7
wuip/QQa5JYzUw3p7KSTaOC5Ga4seGYnIemnOwgFX2WdI7iSfbsTERgk1zEb75X1
KPy98WdF0JWSWxMDhqrIKiJR6UppwagXBjDSZ37WkWgNyJyXo9oeMLaYXyBd+o4t
ex8+XGJ33d1t8GNwlMKk1zVkDwv9gaE7WLUtHLW9h/A8tDYnHWAxV3DaZJyIV6wS
IOcr8IjtgfNyUVsi+gw1A0MfeovMcWSstGdsFVL8FWg+rsq/dFbJXwzp9vx29wdv
uZuuNGB+55sZTej9sbSnF+c+kdlwECIlFEbPXG1+JO3pIT17zVE5xhzLvzwPCS0A
z2iTkxXNVm1pr8NAeVAZVkP1wE+bOmk9J6n8w9iVkbF0GhNH9h4JFa7z6K5cnhUs
0wv2tGPLr/Fe9hy8Fui2e5kzJ8pTZtdJviWs1rOrKy66t7qOldl0btdu5+4UABWQ
1msb3y0pVvtm3wSAeOgfUAHVDrw5dEmFj+KIkXd7Ryve+JgaRMqRD2pWomBUc2oc
0fc9du+Dm42UrmEuKfV8PLn5++1I2X23usoe0HKiuRLJXUFn2HmQQhEsqwUI+wMp
f4wFwg63v8CJIKfKqV/31OTxzl3geVbwrbpYeX6fDcdrREwlkt2IFvllaKiWUt8s
LqEOc26txqm6iRPL3jFWBiqBtPSjzItkdfMFIW9u9Cy2/mgjKKmSAHF8jXrFYoty
p2uLQfX9h6ABYrXD7Zw92P0WSVYyYv/I+kh9hF+0+Xmt3Ji89TlxqhphoqDcehZD
sKyz69S+F5y7kDSKJoRD5HzTfMGKaj/99LDPi4XanwpaMJ2DtrLhTV1ZWdTzYuI1
h0uo4FWfgx7o4EzN8QWgVMfvgx4LEPvnxOrUppsQdh1/liJL/VVV4GM8sUStl9wE
3X6w+KV6pyM80C1SMlywWRtGvA1vhCxyMG10Bi//zQb1ZDQNdWMEMEb4zV01AcU4
nvoSTH6w4hoVENA8sC4dygtplZP7Jfl9vVDP73lXxe9TjfAHJA6VLbL3x4jZyRho
D6OFHTLJALS2l1DPbtPAbvicmUjo0NbHSeGupzDWNf2n5kfVBWjiKCQSqy0kYDiR
3FnM+HROH/6tzbyGtRVgOzQzyylrl/3f4jcgiNjSPGBtQaa8zo8Z0R2AD+hXQPub
k3/V6NoiiXtbAwDAhRpK+gm8+Z116SZ2pYhxPzn73HMs4W3imVsm3D6iiuFgAYBV
9u4wwdZllHYcI6n0adbjF6MkLDf8QK5mzbAVlIDp5pHUJWwXvPPWUqbW2xCfrsE4
mB960mb0DtzE01o1KDQGRahPA1fTHtx1AU1humvK9hTTGgWUyiYzIh9x8O1z+Gc9
gUYx3xK2t74mjGyftImFj79CAwNLeceklMkj2J8UlUPK7e+zYalZueUU3PGSbOZy
R7c7dhoT9PiZMoiFqo8Nh5wTMrMJurSDTDhGQvoUb1XKcQdCUcv4J3I4Ar/nID8J
MVSLnE5emBGiaCCyMQ9cSAl39tORV+aBg5B0Qj8VjcvNhDzW6TPlhCMX9Jruufo1
1/8uMUsYyLXfrUBCRAf+e/alR6+p83GUdVlkFGs0BLoP7djmiqIHBFYUAL4PNtNM
ngDeHK9GF9pP880M8mYCjj2Q8FesdZGNjV+sbjBZsXZOwZcdzWAvyhIABFvDwr4b
fTaRBZ36LuaScT1VDoHjfAY2Dv7bqZvadIWVuGznNnNDOH5pru120WOsoo9E9Eec
TPjTQy7PTIB2+OZAA5WUoPkEWOgzMDXISM06QihV7hNnkhzqvl/M6GG/dqZ14LHQ
tDrAFtqS0PMVHI9MunOdfjsuYoq5K6sSvDWjiAbj9rf6UH1Wg2YFOdmmJ5DqkwJE
2Cf2SFyV7AwrWQbQzt4/sI611u3SGXJqURP//T7MnSpHbBiQ1FG/LJ/9Ah/s7gJc
dJrSqRNUP+q3cYtZGXdaZRu1avfkUj2chPkHIj/NcMFn2moR+AMIcwIi/v0DB7ML
zfm/3md6Xh1PZAg+QgPneJe0Mt9y1xCU36rsMEkMMzGUKJSg2441wxjGkY6yMJfq
XYNURwZyM63QHBq0bmS25WZSZe+hlhT5DLiArBz/jjMx1b22bXx/Hnucdvta0ZKN
EXHoiJMOstRbTboIXNPfT+AoWdD6nuiU7LQdDSInNq6G2LkhPRfvrDFF+UchDdRQ
U4xbdFDzB8k7bGTTWHdPv/95imR5SZ9W2dLJHcF+GYkTQlfmp5G7o3xx6LHo0son
9je8C4JTY3b/SccLDIdjoLwRicFX7FnbSocpU5ylNfC/+CMiNKaT5cEyjdc8YQgx
B1aU8DPunkYLV6f9s9g0bYNIIUkaODF4betOL98ch+HwiEXlxfHN/vAO/Mze6Ftm
4uJX9RPZKzXNH7o4hv7FMrP/Fv/+dpPVRvo+OC++lCrS2azAgrnhXoj2fISTGXrb
YtPlwkmtjcMjKEp7cHMS1EBBwrmMGBe9ux/SIGpXPffJumEZpCJYeXxIKHF0GIkH
QOnb9iAqTVoE1DDe5j0EUFfIczm7e9t7UvwptTjOdnVANYp08luhLWGlHGv3T5wp
4jAPnKkprWBRxIKCBQcJJISuaUN/hjvf1b/t012JYM657NwlmTNGjVlNOPpLEIwn
dCpnWnXyyi3y+eFJOxTmNs6hUN7tnhHpkzdTJzqPFH2xwGalSdXDcW905nqBxuOn
Uvb4TCiQtphcT/JKzjjH0GMdU6WIpNvdT8hn+vV3DV3+1MnhPfNQZoHiNMr+peQd
/E/XECjsv74FCpL1O+1VuK7kirg+3zD3enDNTd8o+sF0OWSYs1cbmdep2shkjxAG
2NpFcdYFk3chqroey9R859MN+dCWd2cXVZSEAZZ/c1JDeIzEDOhUTRphd0seKU2u
Cqg05a5lK3yDskdINMZ4kcdKGu0JkMD/3056Ljx0W8wB4XRCYvP3hejG24tXzKxF
NGsqPPnbxkP+PeCTSjAHdHWYnVO5YnO04YzRB86av4IUE5JLROhPdkZ6aAdSXoAs
Cz09re1fH6fesdxv0/+oiovKA0DwMlHcwQtrMC4Kbkl/5FPzmq1GxA8XFg+FCOeX
eTAZHXwbyB/9oIfwaaWtRzFYY7Jmb44L5gva+Cma1hObF3VEWZFKkQfoQAKh6TvK
0YK9KEepMTWMAkfms7AyvJcHO4m9kjeco+7cQJTh0LIIK+5xdJde+bcKy3RdxoR+
lBKX0XLiiLAt1/8BwRU6pNJfH0D+lOp4r4G9VqlvcfWDta2EEAWPiH/gvX5d/sCb
xS/7exg40C+NzzRW9ysTIM0gVBVUOf8n7FN9e8slaeYs5Md3BWtl+aPWkPE5fgvm
EdKzBU4pdB74FN1mapYGtTeNSMsey/LucvRI1+0DXIrYuz57doQRD0BBJjIzANPS
uAnqrZbkNzjO9DiGlxCUEPhb02wtH1N4uqk69zWCvbKNGpemjlzB2G4EQNj2uIEw
TVvnPP75ElB0f1JRfpMr0wBj6P4FpxMgRwr3JALeHJpd+b93iU4wmmbDT/BEadtF
nyf1yWTmApCLEv6lgZEQ1Nvo0NBw7ckEhdnYH8VwLgYEhB7XPSUpi1qsJ3ey8TYA
sxyClan4G+Y9+d+yF7LilHKCCMZL0eWOyNnFECinqnAq7Cw7A4auQaoHqMT0IBl2
Owf3kZ4knRKTuqq2MA5aN8+2sQSM9L0E//L3XtqGDah38CFPrwhua3oeRKh1fDf1
MSc0+PL9rN8yfGi3E962oWRbSMUHBQyF6LmG6bimNyhTNcFDxd5B4iVsgdXJVs1a
hdm5Ar3VWDFHptoXUqFwo3z9jDUyYNzQkXH8wIdRJu0mqo7zS0A98ecZmBNUZCE0
JSJc0pZV28ByIrnoYyI11NFY7LH3x32ATAPwoBrnalneKv43OadlCTNKydA7Pdjv
PaVeHR/ygZGouxPZbB7wpNdVAaFxswvaQoyBcAeH4WjqiVLqSMqpQpMuU5R/zx2y
8H2xfzBVNAGrbkhjMFUtubt6RPlTlILWbWHxrY+NZQu/1csQcKR5n+zqoQ+uyewF
1TVAocSXH6ZW2RzruM0N/9S72S0wdnMUm9QjJXgO+//xZJNHjABFK6iMZbOrT9zc
6bEUIyCz86LLqtqU/QmGHAptYqpBNtD82fHnBnKnRlfhAgmYbG3NBMEISoxjPeWM
T+I39cZ+gDrOTG1wxvrwJ5mh0VF/5WTfY9QkS5B0H62bWs5mrt9bE/1tsb99LX3E
HlRL2Om3KK0HxqN/LhckmeyOYTEpRQYmhIqIXflaSuUOesegfo3lvLR+HBBBk51L
fr/M5+XzPOKK49jmV/9Ga1jcx/F/IJHJElGXuZAttISr/2uauXptrzu6ePTmf7p2
tnjcFg8oqit3EthHWT4+lA7tN54Q/oYP8v7r4DV0r+l2lR4jY/kRmp4clCQQ37Zo
KE/5gcxQXz6iAumbAxBoYWs58RPEYyPJuyIzcXME0td7uAiZm2xy08uCLj83saod
vtdGie7H+4fWyBNIiarRvKDJRoUXzsQvQvlYuEnekuM12ayNT+eodGoT+okiS344
iFg6ZEOZJy6G3ul3xoIypl74etuFbC7ampjYJm/EVtLGcDdPtVznybeUAx5YtVS9
Td7Hapg0thDqH+vNk3cKcUKB24tV+98MC7HDzeV2pPvAGQtFlZLhnocrbaJaXed5
snHaJhmgfWA07NPVbWN6KJ9buZcVppJpjU4phzAEMaVkDr4CbdSikxwkzjWHFzrQ
TfVRJVDlBfXpgqaC7pyQVCNmDSWPQcrKM6UN10IciUUl5qVcBak+8DeqsXL9Jd4d
MsAr2kwlL6dXWVKArxmgE9CVoDFtS/GECOVv8FhiOvC1cSo6um4nZQc6sEDvBQ60
8YS/Vy0ATlkZHmZLEXTvEJB1LksZHQXJtvwxhN4RwjUXxBvX91lCM1HsceuPRjGy
Q4x2smNIxJF0+1qdr4yXyf72Ty4euEh0ymhxwLXXYg3hMaroAxOK49hdnLWEU+af
r6Tn6lbE51b3zjZ30qFI62Exhm5IG7aH6Nb3QbNRAUGgTk4aC+9tNQ5XZLP5CJJ2
KDG01ObqfRkPrymG0ZN4qL6Q9FJwUWHyVx5BKAerV+VI4XQAZoF6BS64WnJ2ytlo
MowK9vn8D/78Mwul9sa0I+G5V1gSuL9e8NVxBPdZ/hHJUunUR4jZoO3e8zKNnk/+
Ymkgtz0scmOjcnudqGz9uYJpX1VKx6+XU/K+mKtno5r0Im/A6xK4XLBwkkLclIzy
oUMT6uBcdIRaDp4tzgfRJDJab+vjyHsAyPQU29bj3KQ0l6xH6zG7OU9do/fTQHcl
IwKYom4V6cQrIbhsUMi8rnu7Pt7kc6xKKmEiuv1dHznAYEv2G3CTjcs4K8bKEu6x
Uxin2A+glT5a6E37NZV9g2mEpGPVT9sN5Jc7M+nsOE342gYQjOoE3EKGR7EDsNTc
Vv2MlBCjWY7e7k9HsaUSIVP4koxAIBRlVtMqygaRGqjmYZndi11j2PLGYFr3N/t9
WHxUqDpLdqT797q4BQpLjYVrchQE8Br2iNEU1ysKtkyaxYjJs40ORRA2a46ueUSX
THGS7I1gPOn4NaGfkN5gBiFNzMVBZInQbe19af74L3ioTJenHMwOPl97MyXmG530
iiT+eqT/sC2ZuXDToJC+Oorok/QsEzJvD7a35lseIKiAJaQKQ9ntMrh7WynMntxg
woDfgQNFLG3pQ+MmGlG6gKDz3GD61LtqZLn7uwaGvhFm5UeqgUTqQdXbHVUVYlot
VyUJ0pCUaiiaoxKtHL+v7aWJAcy486nocoqDOcv/Q+O536/EjfL0O2wAzKYOFPnQ
dUtnaiPV9c7wZOWn6EP8Aglx24z77pUn301ZCvCOJm8tdlLHVSei9nHTK1ybu9kz
deCyjTYL+W0EiyPoKNffZheCw66LcXw9jBw2wogdLji1nWQj7mpuAc5kb6dfrx8e
uSjUMhBUiGDjYlBMCHm/4av6+7C3C76uU/H9MBj1Hf++eRvxKqPNY/K5h5i4MEsc
2VbBVS1uDSuvhpYotYahM7yAIDnQ1BU2D/R94A53Pd8sEtMSEr86bheFxQSKQ6ns
1gSAHMbJxj+uXVLplfYRFgQgCEZZ+7hopRfaMezFImU8mrHIGp68L30SfmMcCqRH
9mbv7zfRZn02IEj4hFt+5KEBy90WqnENGFkB51FeMcMtFIVQU59ZpDKcsJDvvjt9
oKxluhfkkpP3BP8akokAewlEzcSDtq2qun9gvxCLBHvcX9vs0pfTDmd5LqFJ7u33
xsQmmV1NHsZN8ewnGQbsoT9YHoiPgprYnZTA22M9wVm0Y8zbCotON8DUES12yvI9
cOiUDnGtxGX/ipuHxQw1Iigx9fQwnThaeSLkiC3jkgo+M+MMHmGsW/NlEaU4h8O+
CPL9CWNaeblL6iNsy7x269YL2URV1NiKD8EEwImvbnGE8ggMdftFEf4eQqOs5qMm
FsKMo6VK2fH1xLvu4f7Db7fK2Ai2TdUBkffyLyQHmfqrRbpf91lZewQ5u5+5kbrk
15Y0ubMzbo3VNRAzbDEZdu6XH0J8Afx0j5QzW3XHkz1zjHzgP+bvIoNADPY/wMpL
qgSexCv9wOEkgl+Fb3zUpMiz0qduPlT/scainj0lIQfsmizVXhH4v88PzK2T4Phe
o1hbbnG6bJj/WZrCaX5oPrOqOyv11SQv4kPq4CAE5uxolubjDaoH+br/YPyGDpwU
NSWwNA/Cozpz1YpccrL0ohI5rJgkWZn6Ioi3yNazRX8pbr9as8f+EocviSpXXToD
CaM9wt9GDYNFx8davgu4D99aaSriIweR3HOvxWhhHRUbG+QyC9TPIg4vxd2kZYi4
jGSctjwqGgI04SoVX8rbZaJPCnQ3SsgAwcvKPyahykEPFrD1jEWTqByovRCHH8XX
nczsWKE3lTYQtxE6/6stjZ6KBSFwFAfKgZ8fWKS3upF+nWS9zbEoMcdbOGgTOc1+
4XvM01lMycYGJjUGNOjkqtzTxbutIiHiZTXX8py+jZDrfwR7Fnr0EnSKJXFsTRvD
ZJmLV4bFPOWCdzJsfNBpROcucXaeRRl+fZPf1M3sbvyXVjbJQzRbD0KYO3b1legC
OoLZ3K2bkF/2jGAQMxRjnwTQWUTcvcl+cg0WsUKtt93IDQ1asBe9xxz9GExTj1mt
Wgo8JkQeve5iHOvzXqVR8QeWKr7aV6Tz3rUIHliTxfRh3nhWBIhEro3EK3siFOnx
0jD1RPLs3ZN7GTRq3sXV4UnJj9wPC61yIiSew86sQU4b/v+EDZ+v4wTvhAIEQkEr
lrVFceo2hYuUuB2EDB0BPurOICzUnYS2Qxf1LFnssXgMuYqg+BIQhg8UyTbFfSjV
yRS4wxSfT81z+FDHRk/zKsaqJhQ6RMlTzl+vxQVCxUHi/xkZDkcnmrFPgctY3H17
q2wEAr4p9ZWSmpLiXDx1w/lVNOaXuEspPjUvRU1ab3jzr/wq+fcRKnanb1J7WZtY
6rqFRfFblT0muqXmi9rZA4Q7V6QrYLnMKAdqMcvInsepkyBwKW4S6EjnAjIdS4Tl
dNdcb8g1vrOEq1AzYHYdEPolCcTE8crxJpGErAyv2RCsdzT86G6gUbw2DvcVUBmM
XN9Cn6qUXuX4R4pTFk4A4mNajDBTmIZ19gg4hShDiv/eHILLur3u37kR1LRxXLbR
cYfJSMVK03gEVx7xLthdIt0Pr0TJ6Bubf9iWTet86ggPKNZ6zomADdy8puL2ZjsT
rINeg6I3JI3w6RYmq2sKThK1ecydN28FcucnCkRfA6MYy97s0MekeRnxCQ/1GBcO
bNletC1evGNN4WOCO/7rkAQ0KScWhha45cFbgI3qMidcE979+/z8v56NJK9Sz664
OKl8lkvQ4J2RJIQj/UU93g8cGVy08XBP7qF2y1mDF0pZpQRW8euICQf1Ee5L2zG4
LroX9qlgj4vWV0/9vqEvGkrL2PWdyCNezwgTcJn4d/ACfEziQVMxT7H2xRTB6Y3e
BPX139dCdcvLHR3yrvw/33f9PuBfS4cSI79IGLNjlqmeHmOW0J0hUHmoPeVoRG3s
KP7PDRIaVEKH+GI6MG2pyv91CaREytSn5vTtT4fjhQrpqoqzK90eAZGWQ+YiohRW
pUbVX2FUvhvMCcVg41MaJTRghlNhshQCZ62wFByKoNdlYdXnyVoBccf1wUGxvQsz
EYAzNxwSGBJOSNEVa4lU4sOp4CYvEBRGhpt+MzXFqPhCosAGGJr0LRlwerSlb5wm
vUUcypDzrA71Q6wFAR0wI5oES+1jhgNirunLHpNFFIoMZL5av3qEJuX9pr9JRi1E
dJr3WPRc9RMCAL1oJK5bF5pLk9tJypzeEh7F+dyxxkZ3ppEn3AKFelMDjEx+LMfx
0fS7w7uBul6PakLbPHYXMNrhivIki+UBJwv29S23paHkwp1l+uwQOvKmYGMTMV+Z
ZyVsqU4uY2dUMe1R79prJjT9Z9U3JseMxKhR6cl+t9iUilnsSDbVCPmo/3RTnAFP
mER0/XL7EQA2bNp9tvkkOWxhcf5WXoSYKoVyb1+Tn05HMkeWfqBWsmAljSvstvnw
kw5pk6RNS7TRA4ZI4zFDWpoTeZGsnu4mbFXMX46i0MSrf5cuH4F+Y9iBsbcek701
3X9CFhgmGpnE3xRUEJshlCHK9HZBRDCxw7OzYWsFPVIF86LKIBmSb1U3KLie9Rv4
bIhRJX/PPV9RH/6Y4yOfdlnLyVLXJisMwXqP3Jtu8urd5jtOPkR8kBOyGebV65ae
z+xMT0u6b6Klly3qvfpiewopYHb2/XxN3fekCIlr7NdvNwhdWDT5P6C7rmvRwcYI
GU+OOi8NXNGrbi5ciDwxGDKe5e6M9ZuCe36mzFtn7euwnkyD9ETyDi6rLje6Crca
xPFqxS3VCq/W4cVTeHTO4HwHSCVeWmQpJRuRVkQre6bzMnggVPXcUAMx3wBa+JZI
rsN/01lWr/H91HOUb/NgwDVhQkH9owjBMbYfn7JziKLJao2XkHurrosTFJ8O2DwW
VGgAC9x+wORAaVIsJSqcTGXtV5bV30WzxzECNBX1usMSFVY89jZh7MIX4ZkIMM+o
lpUSDHiBWX87N6uEJVxudqlvUTXsTQvcgomVkE25GzznCIeJ89kj0xmtv/hCovsb
vDbIDwhVb30xfqZnVW3D/vK6zkfhHdq0hCFevCIjulG1u7KyMsDESdCioU11hOP9
buzgANxVjuXbM8YXyYgJYDFD37pO2GFsruYfvWQrx6056d4IaMLYujv4TutGJPRp
i4IbF3ZZ9eM0noQeaGJe8LIU1WvFNIzZ1DVDmOsvZhL2zdsuWt0iuuC4ShoaDX+W
UCno7rdK7nLCYie9Tx3qjpbkq5Nnk46gyJbjc0MS92EKzdaQmNmoQhfyZ2G8E6ws
KdtT52kFRkszAcHehKInDl7hH7zzE4kTQzx/q+jjxqpTRHf/Jbv9OC0EMzePuN/S
rithNWJxKaQ2Gjy2L6sh6u9uy5jCEGx7DsZSkUoZE2qHwygl2j7tQYapeyH8BZUF
ksNcPrgjtL/Fec3gubsGH/6qnuKlaYiG3juDeH4oZWWWyJQbASzSYEUQlkRSTxj6
HDWR70a1Cn9S9uXJCOMNRb7qEh2AnblLVEJFuwtfDFLQq3GFf+vfhbn/SliS29sZ
yulAjXni/qLq+/NwhFW1A/GdwdzKTLLBArlO87gg+w8AdedlBH1L5dLUxMO1rPdu
xDHpuKiBcx739GwIBjDt/kcKWmDvxwXAIsFA9fFlhLW5h65PIuNjYgmO2AkPvtVp
hqDlnhQII/Pd0sSUHB1Pe3EDbWMW7M3HN6gh/Zk1f16hE8E9E4qJEy1yLF2sxJD9
gXIjP1rA5Ky/suOEazZlBjgGq6n6Nhg+HgeGdLYZZCu/yq+ePQ2M4Xr2f5Llm/r9
JyoxuDzIIQJ1M1roWrqEmsMjYeXoL/hpC4q4xDRyjtjimBe8NVLkKS4k5n78nTuU
iZjON8YbX2G7JoGoAnfo3XfeDdhjcgqTnOsvaUVWogXYn6ehOuTaC7vSObk1HDZS
Dj992kDO4wXpoeEC4UdEYwxnnhTdAMlcAdFY3xwchi3BRetEy41DpZLFzNvzyY6t
TFlLTOOGnkg8BQJ4dvJkZGt/lsNuO6BOT+EEqZZQNbz/NWGWEWOk7Nq47p+ducP0
q40RhIb6ZUVgfSvO8wX9g6XpWBk6y6266zmpJr7p+2lzmWc1QtjB2Nr4G4cz4FQS
H/wtJSFC9NyQ77brJU2OzQgAG5il7DMG32KF8goVqEWmnweGwUCrbDpR/rhFSF2K
DPgq6jXJdZc7P3fOg44NMIFqCLE2477KnbR/934PLYvJ6k3DwlGEKPTXn/X1zbzi
93Y3szx+DP5AGEPf5AjspG7AuITEyPxTGjpZdbflpFNbUP1sxLlxUekq95aria5E
IW4S+c3tvq1TPGjkyRwbSTu8hAR0+9+HqQ35/6Fmd33xpg2peW9xFwPq3CLEdStK
PfHyxvaFCKBbk1bgKAjOf+fpocqaTR5tdyNRPR60HmkkKHiQfDvVJJEnkPQmf+GF
RH6KCI4qqnWSumbxkDxcTGV4SCR54dhvTdTCPlq12lvMwh8Xa24o1QHqCuYBDTsy
SEkd6z0zO1ag01RDUrWKBF5wcJUCvwW9XG7vPgkKqrFHFL93Z6e654w6mLZsr8OG
o9tTinDuo+4CIXbHp2S8YwP6G9nwkTZMYeh16m5GF0MWIj69fU1wET5CYOtgJoqc
pLhZqDLMQ/VD3/OV0rQcrYvGjK4Q7tu2QgftLZNsM1miVUaLZscCOo4FCCKW41GW
KmoPTtWK4fxg8hv2knMTlgynkaxBTjZ8brAxjhORCqG+wpMDzfZb3OFo9z9L7yWx
zXijvngLz8noLLHpEbIBLCwDeW6C6eHiYrGmG7wXCdnT6icnrhsey817TCaCwQWu
WxukC1UXhdTRRCFjx6xYPX22w8Hb4xFwKA+od6Ja1j6FhWD6GKDY3E99JRDGQxR9
3PzTtawanPVKRMrKSK2L1/W9fPov45cbz4LIZ3/8CaqsmIwL+r8cONYdyDguBGEp
wBZqp2DqC2fuNzjQnEjbsv9tfgu0G0TBUzBM773Z8Qfxt07VbK8E+7mGx5T7N8vC
BfVaTDo8UTmIVJNIFsAr470f8VzJj6PnVoEAKqc9R+229171r4RGrcvnHwAFSAaO
ghFpAAuWiI8dRWiTlYEi0G4/AFld5Eqx6ju/dU4Ash3ulrfUQ7/2KZuGJOrFoZQ/
DGRPPBdyCr9ZWqvDZl6nK+bpgKNVFcWPSNitZRFVbIn86EY0OJF5O1JHFivqWT0Y
tKsbSUfNvcj7q3GfidOrOY4ZVjZyYU6llPk3a1tHw6d/95hoNpen1mZFJRDI27pj
Rft+M9/l+MlrE/mt+QN1PL33N36d+qgH5f97XadLWTW3KvqnO7FeUgsgZZvMVdsM
SIgY2LZNH9m4fynpjN0iuvwk38xq/GrBJGt+cndsRzRPXzgJf1+YksqltOPfKFQZ
tENL0P3/RzIGM6+BhgehGgXokwAd6t7Rl3Q1nRfaPhzYc5C/hsp+sq96i3oaPDdF
vfYXTGmFGQZAOgbniKQUIEm3unb8DNcd2mypR7HS08r3b+tV+yOBs+aE21qAyCr4
kFdu19p0hPSrJ0lnD6QEdeVoY9OrJIUA/fHcb/oOgaztn9ud1cpmelHkGAQhuy9S
8Xt1ex8towLYaDLR0EpNcxZ3VfLjpUGhPZRoPWe556wvhanBOmRTSz+wEP+mtmlF
rJxxLHTskPJKkM43PG1JMrDyQlmBPbC6420FdmDnIlwauRlxaSzO+T29lk7vrzT4
N9qlESb0Txc4hbrm0KQ1mTXiXnYET64JF+v0Uw6PBKKdYspg0+Ae2kSj6RYUw0+J
fQwSH82W5294dgYJ6PGlnLCtsOSRSNZG/Ya8v1G6kz51D6Y3Q7g6jMZsjKuyAake
IpFj03iPb0pkIVMUbjYTDDfVsRlowEgic5zuJOAl71ysWrKBgXKOAFhYEBKuV+aP
l1lm2u9sqiTSvITuTBKlSbUJJVzSsKLNchQy+LFRGkEAlNPHtUSqAYtp8E+X3SXZ
HQMtmCbOy+IjQXAD3nbH2UlRsbBC4fF3MK5lbctUvMQ1mHhY8O6074tglT4OUhuw
voAHX0tooio5U/PIHwuhvgNg+t0m7xSP8tTSzTUDgngCYhBHK3T2QdquU7fosI6Y
jehP3jBlfgZOLbf7kUHRU2ODYsOmkXVUMJQK/jHc6CLio3e2db5E0E9ICdrk5oPh
g4AIuUtRZ+6jkoDQWyTHrJESRUjcsJC3YkiEB9dtHThdooo8/Pp+fXVopSR0K5ZN
MQZLQW/+35jwNzyKwIfsFoVU2XCwaR+VFlCG31jv1L+Gp1zcCjo6EgogH1SObswv
e7m1jl/UDUj6UFmjbL8CNLHd7jeVGFbXoME8wwrRFpXWWS8RV+4ylUQOth1Y07uN
JkpOdw0OX5Co/p0EfhFOKWOyFuqCotKiKZ1SsBbL0u19hHUjPmJ3ZfquUui1amsj
+8vUok3uH9rvqKQB69wKVL2OWfiv/XYPyGp//ASNbb8UziCF1Nkr8fwdqEsbnH4e
U3wxICJ0fyEVWy2wl9e3en/xjKX8wyz/fmtMfcwHZ+0zq6FCRq4Y8ee3npt1AT1T
4XT8P0O2OHg7lozZioDEp4ZcQKjCeJtrZc1h5PXHiz7/JaKYbWke6BurMZwKDUkm
WJ+NBoxJwTMQb1kqFU7w0uKZ7o9t4KZp8hV7DpdV/Y0zJNrh3gmw1mW74WQ7Yi/8
HEnSo0ogQohCO6awpyCmG6LD943PFijRDuKqR5HhXlz5D1sgZZSvsZ/ofkcDCKpn
XTcWLfYQ+Ek4sWT+KOX93OGRiptA58OXAajG95VvadhdYwFrfZClt+NTXx584nbj
tz3/D32uyZ3hHbrUGfLEb2mkZwU0Wu9CzMFbSG24/NvVVELLN5YY/UGHfNtvucYG
wrCdhk1o4rQb0sWKLdenNMEdt7ygR/DuUY/O03m8s44Vb+EF6e6uK59iCl2AwzMp
0JK53MXvufMBM/iVHj0S0P/CAkLue1xvNEGpuAG9Whj5FG5ydNej+ErDZUvxi75M
x/RHD7sLsnc608YomU5bP53N04wexbWMekWCoEq0yuklt9Imbwj1Gp+TWjxZ4p0J
8MRPNdhbzjXcRvJPgyOSCWLpK3EafRAg0XHaxBRFsZzAFQbi6iwTUCFDaNH4rSZt
2RZz3OC9ztCKKQMmGxk8pCR2GuvWamjQXdZJqmtifNvsZZaKSgG7m4rUUInu6rT5
5xDp+kDCiglAi9qarpJJO3Jo9gSbIByP4BZpsdI4ZB+4xz8dMr51fEzV+yMaIgzp
4GzFM2iuAxuFnPZc0BzWIwfAsATJ1aaBeWDSm2q+NvsUtmOlcX7sVa4TBZVAdxwt
q1RXlhfX4acrv2IkPLseZE47yiZUTIaXPcDNZIHB7tp46FMld7cN+v9JKQz1YO89
YJ7blMt+PnSM7HkEdCORPHvcGVLK9N/8Okw87B10Sk1+eVpGE5PDQDUcTkP9Td8S
iyB3nBRe4rT9kz2mBb5tqnjyGiQjjy8FXSbhkniFrEzf9dzqb9ZbXpwPERFcU6UT
eljx7E/4EtH++JaTfjpiGC/60/Aw6lD+H85SfAecUDpj9v0b3HNoGCrI1s2FHpFt
PyqnX5JNZH0apK4QacmME5px+pe/pSKsJCFKF3FJdnGt6cwwkCwORo9UarpNJ+Xr
jmWM9vlZ7s27Z2xNc/OVpMNafaZ4sKj2ACcXa1gldF7oTqOJ+ju1Geujrxw8hwRd
f0tJlFrbf95afgB7paFCGhzFPJtmIKQ1rtA2wYdkk0P/rrcgxrNmBt7jUE5AuKgL
R94ZTH/vXsVOgHuCK/HgX1wxWtiRs7W1AgIQ7vwRdBpB6lf9QMnjcaHwTYs+kQgt
Ra4HmH+p/e5EFFYTkjf4qEdAuIMcYiXZuPS7/0C0LI+TA5C7eTevmpRUg8Qu+FGD
PmPZXmJ5sXStA1FTRhSG6RaxKZePxtbp+LdGvv/aj7XD0BCKoaualq4vtklUp09G
6jmna5Wfm4C6gg19hd/EW4oR/P59IUzOLHAg6akNjfQlNBNEWxtKpHgKiEesv1sR
8INbB+PrJWzDQAWDRoQ7QQJDtK0eSqPR10oQKH0EWRMwRaEtA8h5aWegR5sg47Xu
7yFUblCqtHf8OIQMW9/2C+xEGemSW4L0q7zVoqaOcMNFGS5YOnERdAb3X3t+7EC6
Wh/m1OUGEM5Vp/SaEL9G3qNEO9FAYtGn1akJyufzEO0P4jkTJYZFiU97zJ82JEH4
9RxI0fvaOlJIhUiEfBylXi83u/+ab09bhi2Qwt6xvAO8XXvsjI7N2JbVjEC+hyK7
YqvCGSKT1N+nJuyaA7asQHlBpWH2uTNySbqrPg7+2TqziNd1OqEuvLLi2fM0lQEn
yu82CsA8Dsn3Qtr0MPtmScqfrx+iBiAi2WWF3grUm3sKaZgvpTMI4qEAoLnOSs+X
2c/DScJCHoMt/ayDazzdFEcc8Uck8VRNCbYGXVKt6jcrFFMBk6+ypqIuKGQdyTU0
mvvP9lpkDRH8CTNDijOSxTNT/do+2IU0QpdPvpSaU/JoyGy4kCVt2w9xYx2eBRz5
rLpt5eILuZUXzk2BS3n3/6a7nmBOgBGmId5AM2znlrJHFKj0Pu5VIsBHrYPy54ni
Q+veeqSbAP3XlGTu58yb85/Fze9EXwOu3c2YMm6tcBPeN7CcS40bc68SnWgBk4Qx
2uv4GbP+yeaf/lNdMV8w/K0hit/8UTjjZdQDpMpjwInLd9auH9VkQCyHTw5leZQp
Ka6L1NdwkfmGHc6Nuivw2jHgzv7nDtc18tXU/ruRkhqw07k/FV9LuhM5+7nI+IJc
ByBe1Lvo/f5rx8B+/M7XWgax9psOoWC71tIFgzuvSUKAMS5CAQTRr/pWDGCalybj
f6D1Sy0d89R4T7RDVHhOrDt/nySUlCbAKRyCzWhNbqd/EUhKuemuM+t9qeWYqj33
O4jZ5+Kgjsx1aqzdaDbu8JNswszDY4Vao2OA/mo9KLZXcGOEXKh8DXfPjxvrBYCI
/4tlZzVWHS/j7U28tRQRGt7GuuafEnHUD042KGcRYzr8BsypLtV/+vieAS0IW6GD
XSeCVENHR8whHyjG0ysSxN1pg9HY4ksRphd3etl8hpoO1FYCAI78jRZ6XPVNuoL+
Tl37mo1zAFfcEcWM7frjaMSIXcIasdFBW/Baq00W/enCi0TxCSCaPV5/0cfdYlNI
jk3G4jZh+Y986G1dEmXvrreEkQaJax5Ne3xJV23+YPGOMJstzcj67fm0Gv1S9A98
Ant2qbw8vLaxXVmPBQ9hAIA3bP2CXAGvgBHoAS9VGJWPxdBCb4OPGnjuz4BL2I6x
/xzlAhEwOXbnEKjp+gWc41cCvW9De+lGM1nuCz0lUMTrwLEaYcfXhTMijDQk1W3n
CMgWarPlATL+qoraMhQeVyBLHx8Fpo1mZVmrcrF9cvv8viIB7xJ5JXkg2yCnc8X3
UPfNpGSYXQ4COlUlA16f/CAoqjPVcKH/pmdY5RXmCMznIROChh7QDXVJuZYq9KlT
kBwohIe8w/5IomF1JqETh71vf3tHR7jt+9rCk1JyYTmfGeEj3kmuUNORIsdRNphe
cxzEBDdMQAOl+r0s7+X3XjeUZrXdR4H7xLi4107Qqs2Zk4pe/PPFZeY7Cp1IlU1a
VpzQ66zzjubC3YigDCwmj/DX3pRDIbXhI1p3XnNxZPCGotQkIanJPtVyUXB/xL7+
BS8QqWmhpKsEw3IYyey1kiOiPhhkNsxSMMNFPc4X6Oks7fCtdzZtwi+4SVCW2w4u
37/0Ci7RY7U+vXs55TSA4zlK/RZ+9vePZiuOuxeBucqQzONm6Me7aXpze7EvRLgA
1mgQ/hlC65vUkSefZyqB6o8ktkkh3pKnZ2C7H9olTQiUTzhU2oCr6O7UV0Tocpav
X1nwLE++B/Rw71GVQbbiAqp0CXn/IG/hMi9p3WQR/cwLSrdx6MC0yURb0c8WKcWO
1lHPT30YK4lw45OMYriA6vpe1ZZWx6m683KIaYaXPtvU+BzKXw2z4UDqCK7f5VV3
wDjie4zZCAPwGEPEj4RnnaYqa2a4akUzM6PZ+X3QDrIeaGXQk5HojZFlGwvKI0o3
UxVkh5kPQFIni2cdeIgPP0dmMzxuXWEPMDmOG/uSic0h5RGqcRY3/QKg2GN7GDjY
ICnKaiB+MIeyzbSRF0zZzEgAksao1o04s1u8HBwRCWA1BphcS45mGcpOYV0t0tnb
FkvHtAevIHtHuZbjZM8H/cQEdCnD3e4ti8lMrGGw8jlId0bZwWQDHWpapxJYisRp
RO1GV3DmpHUFG4cVHoPAdU43LAE9wFqCpw6oal1hdbhwpO7BB5osVDjump15MIBw
VgfcI5Ja0hgbN0hleHF6OMcXv7gcQ4wdPoSR49B8AMCqaQ3YHSVQisLoRGVYj94W
vrgddco9RZyrLSZ9lSeqizX/c4fa1oPbqqMl3S0TKunbS9IgF8HhJ45g3ptjr04v
6MBLGAFRbhsCS3FpmfjZSCEJjctL3Zn45A9Ly70SzLgsPQI1FiAOHve2T5s9Kl8C
xOCMqdZQv87zPF9yZSA9EWztejIDOTl6+BEItsec8gyCSaWK+bUgdNkIQGXAxGO9
2adYneegwanieL/igmD9a+fsMjKQ/bMBs14v9KpUWyPk3PIC0AXKjWKoXlD8aZgD
tyr2tXzK6VMqiGaHiKt96yjinirYCnWJjrqYZELZDz/el7Jz3L6y5QUfBS5g6YGe
DeUdj/ji0VBQB39SsfWG3jFWsEjROgFJ0fovH6444OwgHhgCNRXZrMmPzVQRgDTG
xAvyef6iVfC9/JZoNpU4xO1xud6oK8zCLYZKazrVmoxrJJvqq612hW4Qwl0xpd2g
fN5Ae01n3Gtb2uxcapqzfCafM7H+1vqrcjW927dzZAjvX/wgLixVkcZmjhg52O8V
sX5Y5ewDyQM8nC9mF/859R/dkKpKEsU4xFNDNxOlnHvRfQADofvBq4Eb2okJl7hY
En2OtMJ6Tn1ORZojkQlAnUxLERLLQoSIEjJUjmcMHIci2KOOw9ab4KO6C/4Ue/w2
KY7J7ipe9SmliNfP9sOy5vdXVFy8D4q4wuG+Yy4tEbP9WteR2SoekbuoITulnB49
/nm2/X2dCs+GaWx/exF25gTiNPduR4xBn9ou4fNvUwpjr35EYDwxPrxWpzyEZ+e2
INxTcy7iQiulNZDbJocQs6ZtHcqwS3T5+P4gMl9r4SeXRdMHiGl2A3NSgsXRBF+S
RDky59EAINLlVj4WSiAr8g98n5fkLfW8W0fdM/eYrG3nzvuqDSQIxTMIKmJfi9Cv
qsH70O00zo7qqTPj/owilwMh4TtNi1sTcs//EOFOq7qk59jZsLeWfV3dovEU1qNr
lF069pLppFgfClicDUUE7wgsdX8EnExOnnL/ZhTAjNKaAzBuvFeHtWOOmlEM1KE2
jAT98hDWVCU2Fd8vYsa7abCVNs13xRPByc8TzxtIDafvDpkVUAqxBwDJWGqi5Di8
RfzvWuIB64uMf2AGGwA6CoutlOYbxCLPRiHcGsGhVjbMlNAoU2MoNtsU76IUylb5
H5wZIeeTJek6Tmby5NKi80ZwZyVyv8ZALl410HZZZyATuq9Dc8nUbOtncQ7w6PR5
2UiH2LEIDHjxum/d5ZQnjGWCQVBtGZ6fDsAlE0gp6wN84PKRm9O0tjiStfBTQCyj
BHfrwQ6wKx82OGgMTE4hrDseKvLJBR/SMaP2JmhlQ7SVwV4lunbgwo2642/bxmSu
qP4eqd0MVmHVnXUadcbgJSl0cwRLj0pzCxIDMLfVCK7qNAR92kAW0TS//ogcEHye
AwWldmb9OZp5b4/kqF+APXx/XMOTmVN75alek90pZRkRiVQmiKOgAcY+gr03lM/P
c3Wld5qqNZsQZMAVEkaZ2sECJlt07vOh/odCwgsuify9d89pjLu7cahGAkTegE49
3JM35jU1mA7YeoAj7WVkC5FfFzFOJsqGARMp3Es9pV9JJOsMUwTqgE2j55USRtUi
QSnNFINYTcTVckZTtCknwK5IImUDJSTZPwmW8b0FQxB0hK3ySkKzoU+tfNxRjply
uyktb20zdpKZ/DJ5K6/Ywnmbu8M0Cogj+vFZAUWsQ6mKnCry24IvqRHFnkTDsGTw
tKHCT4p3crnOaG1CC62wG6K4Pe51I4zc/M7hDaAwYBYmtnD71G3Ghgn6R6thVZys
gS2sgW/xiw80bcAbIXJt9GOZN3TM9fQQg72ki6xF9v7lxUX9b980+eVwRXQDo/QH
3Cr/dKmX2L1DQAhq/WOPnoB1YIRs7odc0smWvEMWiG7ZN7pFIaX41pAZ6mmgb2yW
18IO6gfEFfu2KvldhgaXRt9EDg0yItXoa7v+0uc3DRrFTTVAOCQbtMZSTB/meaec
S6dkC6k9J/ddJM25gXe4HkNfs/W9b4VzmfuGfeR9yVs1BVlSzXEMjkmTzLeqURrd
W+iG9egvPZ34J6T+cBaFq8lVy91G1HlvFCEFveG6wRDfBQqvg3MamhOiuipv4dsu
LEEc5Dh3wYEk+QJLmo3t1/QV1lnVnn2fvkP7v/frfHGk9pIEKNkfq1zCwTq9xxtk
ZL4mQlAsgGs/cMXgMq74esRH+wvF9Myc3d/GtYFcPWmGxkYsQvwYn6zSwnGpj1+M
uKVD7DE4WGCrDTJ1EJ6nS6ZD4YfhVgGWfNsKPbt/Yq6SLVxWLkC7NNkHi1F10geN
Ddcf+s7M5TtcxuucdnLi4bL02h4hMIxT+x0/jeYnPIP4TeMDqgAjc/oTArRbaddg
060FfuPfqTV6hGqtPv0pKCbula4gSWQ86F91674znrmf3AfHIaLj3HCcbYuAoudE
bOyt3eTFoYgJ8Cwc2S326llxGAgJ24Ff0R5KHy54OvUkGrrN6zAnSAvmqvM8jwsm
TA9XW+0yJx2G/4/rBqyjQOII5/DSrhl87zEENmwMG+/4YSesXxkHVhOBTqPdkS4y
ekcFKCyD4inB3NyWmEEcqNts2uXdqhjm2FQj9fl7k7B4txWjXa6J2nQ+40AUM9AF
m/2zmkF0+NAqhW8RF6ZanHXwncni9LvCyKMCX94MUXiwmkdyR5RtRF/HsyjehFhj
X/o5CsiprpnaQuB5W1gLwOVWuy3ahs6cprwv/RtVJo4fM/VerbkT8uSGXqhbRJRS
UmX2wuvSJI9Jeck09LuXMwl0HGFxH91asIgL5Z6OWL7kx3dxRj8R0k6xdj2EMxZ+
GPP54bdIVGMt3zdE5BgI5aUr/xFHmw++rZ70hM6JvrtMQ+LoRNTrsuK4n0h7cY9w
omW5DE3SXMx/BYTU6/BO0qQS//gmChrIkPgBsW8v5AcNUjVsxpaV88li7INbN+Za
uUlH/p4LTWAMn5QWQzTsjwcJdiWxD/4Qi0WnnCc9wAFQFqQpVdkq/rKI3tJiXKrQ
XizyCUnZMrxWYNoY8rPKV+GyOyO3QvZ0Wo9ohJlHYY53zWm1+1XRdb9XsIqTSDoM
1Ow97YajCB+LKd4eFUe0IOxE/oHSnaBSW0sXElFSIhD+3/6P3g5qTcB9rUMPbGTx
+slXzQeFOSruCL6wyVVPyzvj9UMrU/g4HFdIK4PCT+NRIKIZBAVUSGFnWzyOUhEs
S2ttTk0xeJkYZBm+JMsN6zpXs49LWUxCgjrpSCt+8tpW5JsfdhFtaZwS1ucogbVT
Ht/jExOyq8ZmZnmEA5AXDkr3U6MEPxqyvpOeIs36/ghhyv9fksC3D4pS1aZvJtWi
abbY9OH9xKREBJoPZmZ+WScBStqTBYXOCMhRODplxNJnSVxwIQBQ6UGQ2JGbrtPH
r0qdqP6t++ogA2Q8a+64wFiLrHE8EUjAyZiIJz+sawJu4mjNsxvBonS+GBYowo9t
24risxSHqlzbhTO/6w3ACb0ngPOhcSIlXGY1x4KJDLrfRTpKBwPTkLFuMAfVAZvN
XzWddNyx5DlFw0aDrEx7xCGIvTm6+ULGa5NwZGzkiFhH6LBJLuEB3lRNUOBPNhNa
8F2mX/P7b5XieU8DymB6zjXhH1lscwKM7z9MVyogXZBPPZpxWIWBrfAOTIHxGCPO
ELqchsUmzAHcy16T1ijYlNGHI3GSXAelFznmQM63aqvXYTrUV/n3+nW1qZLNw7Pn
hnoV2rmcns1IIPlybbo5zgHw84YbeccTexb/u+tCz61TLSNofiPR8cPiwu0lAVCS
Fe09cUwFGmN98HeeRUE0iPE7Fa20V4hjEiKz1Z1XCkUUABlA+/DyOiSmpk7L57TH
nw2a+TrFTbxNz35ubL820CWjtSH0VKM8ibs5ygqmD5X1yblFJ6TBGMYsP6YpwOtS
vVYAWxvuDUdY/laA7hLsoi/G2ueGtGziqKMr20L9T4ayOC4je66loOodJxWFOx5B
71at+aLd9/mc+i/+xvR45k0iuTkEpouhtmEkZNC/MJAKfMdqgCEyjx4P4Db3sMTe
Cby+RZjb4yGBrIylua+7+Cwz/pVYftGeam1LIFNYocEbl5b/TZwufZ+8hDqKTerL
9p2DCCywZY44tXrJLZEqP6CZFC2PuHsSbzVMuwtPVTzBvXJSTQO2HraG9QO5ly9T
0Npn+lAeROBHNQjJ7XeO9Yu4BMWqB3iIsZs0dEici2EI88IBQZNWTbcGGNtKH00J
nuz/QgICp7CCrY6SQ5YAufa/AV419iTgIUeWIfCp68bk1+Rkh0g7r+m3+z5xIUS3
zeZ0mI0LEl57CDQwA8trsZIQjv30za0dF4pwejwNuMsrnUIMV0oUPsz/b+/dV4H7
XfobDaokKP4I86vp5m2IFHwHH3aE6UNvDZNZQdtQ1C+xNJB5LYx9glfXO7+92Mic
NO4kmJm8EAZYNjHfwY+Q/pC4tslyhcXfSlrvCxY9ymbTPKxOCKoxZdIx2ILoLq45
4RcKHGqW5jIdtqgnasKpDPNtto6nQLmGhff5CSLF7g9vj1me8nvICWwlj7S7S/xY
5lQmjnGDKDJpc18VqodT3HrXpKvVXPRf5r3NER1zVEjmint7ERgH0qm8yin7KLjO
Yqeu+Kj1tmIjHhnKy3JKG/QTD7cwPv5VbPPUs5SkKZnqmROOKeKWnCr8+pfTCzAC
efNPt4xF9PfW7rQiNBtgjbUBpZjYoSpRx2Q5C92DfU/xf9oAYWCJe3XQyjgXKLp1
aUfe/A08XGaoCgjwn/uBu6Vb3Ip1qBJUdQjNMptTj1KBctwM6evMEzqwQCm9VWMI
9TcZbtSew0yEOcWg8bh9yhiSZurh8PHd0jXYvRvWGQfiHO30hLN1FP1p8E4z9m+E
aQCbU4CLjJqPkT7NZnC9eqvAIXXUWQsSrr7eQFJIDSvjXtVuTs2t6r5byLmWYz3D
Oyexx1UZBPWtksX90UVUe6TzJ2yJ+g/mp0Ez8/1CjaZKUkpmr0Rh1vDW88bdLs9X
YKDeFN4DAJJeJAVwTQBZ+Av1morsnLxJxd3HqV3hd1lEiw2/H1WDRm7/XRrjf3kW
a4SHszXi7ovIbh6xPnvLLpXE0B8AUH6OYOGMlWI9rWiF+pnwbry9ih6Qa0RbONM2
hdMt4G42jIFigU+53qA3vPL5kWVakKDb1b+GvGtGo99UdXudV3tnVD5AvbVVN+oD
MDYimCJ4ygabIGm0WaeNVC6cqD55daw7PPtJnJCZVONth8/gPvVWVSGzJIOddtWf
A2CbO006gq/EK4xGR57l6NaIVQ1LSfrZXCbx4C0AT+jEr8uPaZhbAKfumz0WP9nN
sJpxnlW3/dU+5kaHgt/u8MA6xck5goJoqppIpnLY/OPVsEm/n2Elf28oX3zVI9xg
82Jd4DnWVcG2DCPWklwwtWAuB2UuQ/loWC3X1YOFjTweOGVxSGseZ1UN+IWget13
qXdCXsHh6JD4bNYJFAcvV2Wwtwfwlf+MSzOeu1wQQLJggA70wZeKraJwRq1j1WT0
46X8/51osxg0SQtnLRm/n/KYkZn9OQooThU+G9Mnce5w3Ts/0eh4VdMs/tgYlteX
GacSBBj05zV3z+nlYWlvyu2V7+1Ibi1evca/0XM+8lkVzH2q4nJKqVBkMgGC5QCH
2q9EDY58xHSDsmhNws26NkmdfpPgKczuRT6esKdHQCzV3HOUlvyHlGpvYwBGOADT
A+W2oltNYzBDteyprZlg8RyAmQAj2fAmvd9wQqXA/ODxpzBEc6TfOBhj1/oUd6HQ
xIRg2fCs9Uq1gxAf5WoCaUcadpSrsw7O9hs+OO0NwIo0ORFKL4hVj0Nrkq2Z9e2r
vEgecp0xxHzIbImKwy1MOcDUQUbYviUbtmFq9X3OisMpK/GWEC19uBajdYTu/58A
CCfr1UUFs7a54yKY7litT93LuiBtfgGvk6te4/OCrxLit+HrWCsyjtPuPWbzE2Hj
yExW/044hF8ShU6FWnUmtqY49ZJFCe35APGeCE9PMdDzFLQK2kcwyycN9jjGtzN7
R87aj3T2/czZGXK0k6nUOaSmx9FfPXgUMigArFd6uSeAaS7o8r4F7jX/18TIvkoc
fQufmL/6+3tbO4mLzlf7gERyVa0hxKpi3aGilYexOMs5R6nEzYAm49xH6OhfMd3k
cWuf1cNYDYPug6KRkTV7LQ+n+9PIgq3Yhz3EtkRrcsRznkK/EqYnHO/BeaeFexAf
qyn9+Z4hKHyr6vu216vA/EHFVbLuz15S8VxTZJAPkCI16pW1WwsEBnOv6geEnrNN
G/XU+wE6osrgWrRh0e43/UaTjjZJk9mBnhZpjZMwAuhJvoxkUqMKl3/DYbo3atWd
7O43B0Vax60OxRdrqUwdOKofyFcCcUI47OykqNH7A5mvexnMpE4zO1ZX8IgH6kDV
mrui+w+5ker2TxMPb60pVDc3vTyjAEEup2iFptHTzPibax57EOoG4L7p/eDMumXJ
eRiJ1n04D9R0zvYN2hGgRjAoJWksyPNDKZoU3kJ31l+ySTuDSt6Z/QQwOb8dumuf
23n7vSiJuy4iXaSK6pb4JM30kh2UfhHXke6xYR4iJ/M4RqKMdDuu/wNM8iJTNE2B
VPsdj+I0WK8RLecSX1Eo9OULpX+RrfcaPRauWBUyW2cwk46P8JaA46T2d1TC2+Dk
WSDDOWNaOXjt9boAIe6KQy/WN0gv+GhAeUQW8zjTB8W8JlHYizHoeUbUcVBdupPo
rvyeIUADjBcERbP+NhRVpWf+QDNpW752m/kTkfBDWId5pl6tw83CJeo0WCmPN12M
FPzAcBsuGPKTTTuKTUVt9eM8jpbCTUkBwu8qejexiDuckikbq+z4f9JE9lw6OMnS
kuH9nD2NL1DBccBUmTr/sr3tF/FlNvsrHR1bSE70XklwDVFXsDC9u9YhvQiExIKE
Wk7RRRBw+ftNEiJ4hrudigYpcW5ratVXRpWWMbItAqGmtxx4wY5RuNjyr/jTU51G
hmvb9EBZAiJ5ToyLLxVeWvrTPeaff+eZfBUcrbXEYHb+7ZLRIrleqdWTlG5UaJ8R
5ZFbO/vYufZkPz3fP43FDo6w8Hh2lkrnfHXYYZ/jF+Xx36Nl1XDDK7v2R4rBWuE0
sWrH+lk5prVr8RFgx9tbtw5aX2Q6ucQhjtyBfkXIatsK5ruOQZ7rsAElymW5OtRg
QvGRqH+IUg+vh2odo3h8XwrsruYWW1HpzB9PKP3PhySx/TTNAtwOsGNulAxe5gvI
6AAWykO/e/PgrTV2Mf9Hg3fJH4s+w58zeG7bCGdUzgo3AJ+tYmMDgS5dIGUUlC9t
n/pN9MORhz8glikAdiLsw3pLOsChN16fADMBazgokQ2rsb/3/7Rv5jlID7ORSaLb
qKIBnJwUJCZ3xIHv5Nb+Cs+iQlQAF7E0vS/60Lvme+uzM5PaaD7JmwJJimoqGw/9
ZwKjh8dZFPOoZq+QEISTEs1WYSnHpmc1GE3hGE7MvjSuZ1991PmqcUHRf/OSd0mf
AJ53pKXF/jelsIAO+fcdmM5iSzS2xGOlG5T3QDzy3JuQl5ouna9H2DPk+1H33R/E
JmY9KMKeB7oBM+AohrSAwNWl2/qnVRZojusiwvyeBs2+0i7eY4WrO29Py7D7UGcC
fWj5pD5F3MOooghvaKa41ZZll4olTb8PENBv5UHKB0Sy3Y98s8/34Uy8UkoyawKt
GE3tWG+VIThjVhYoh84hNhrwi37DHZKHj2hasicdOxoOywWbaVds7gErylJBKVnX
g4evrhTelgum4fEmFt2Gbrr+xfaQsqfC9GIGwbqvrEEnphDT6HGw9XvYLNF/NFlV
771a39I5seLDmRJHidmTDWTwaY9LR/41bO3gdgUMin3/EWHO0cq9fYy8gZr1D03/
hc9/XeGEChdzsDr1bre/SUyUIIvIbsdPKLd9PZAMSJ85VsBUc5NGJrvdXbbBN1yU
wxzucmukB6Wt5lRplbZeZhd8AI5EQsk7QahJCDugVpGKM4kabGx5lzN8QZlycS+h
e5wcLsPRGP4KKhxtkhWK5vEVl5bocdIFNs51ACbuaqMC5A0iENMbBBpGvI3ujmms
pjNEXX5fSs3rvVH0WZU+VS95nZ9qSuntwsiDERcY4CgPJSSgS4FX4DigrU9F+gdI
FMOGjNVme3I/SsgLMn+sNYTumuC/MDuGnjHZZaUgNTcB+PedmbafGQKszh4rCAue
XcmZh3ReEUW6mUHvvj3Yu/cc1/U6CA8I4LidWdiiaRmUTPLcxmIs6aXRllMR4rxz
hlgiEo08HbdQOukGaNyM1XEFm/dySNjLw7WSBmgCVAQk/kPG9S9FfVqgm/mBvcnH
x4ag/VCe77JrKrHXO1ExFYGP0UlXDMfkrkm/YKI4TFnYhTngR9WvdWgXgy1J5VNj
BLxf7rIGUG+hOjCZny0W4XAS6YtOtuF9STDH0p+K8tlfsvdeXtY9bqtZQp87NSnM
O4ll2cJIZEATD/07BzW2kfoYA30ahNKrQuPGuneALSZoqCiR5+pNre59+Y0EOncx
N4yOLMCuMNk4KVPhqkEbNIJeLwbF83YwXXtcTM0noG7//v2agXxaPeeQ28z7SywD
3CVoxxMvgKOigdsG4FCJVrqU+ifcwpf17MpIYDyzGz/7twsjVvHze0jAFHM0IHn3
4krdHkvwyEk9eX0Xp0UnYH+w5HHIn70OZYs+uIOH3RZUp1YE01wX85hN8xGeASkE
lZIRVKHN8M4vej0m7Ntc1MHR2RY6l7pecrosXdW1qW33Jqm8wD6QHpEdlmyrSFE1
AdumGeduEH8twGgnC2CqGcKFQ7LLMatOCHcQHV6YGSqNIbmQsAlNelCUtqBxwcDv
j9Wx4ZjOYj/GNkcTAooHrxFCg2lHP20E4JTtN2VUt+7hbpKiZ60HTrYEvumYSY40
bpflsl5pQ4kFm6ItSF5rfeRNiKB2ttM0sviedLsLElC+ZHGRtnMIfcmNT2vvEBML
bFQ/k15pVzWLV85TfWvMByNUDpFCqub4fpUFRrrhJo8+0TedSIMFS6My8VtcgQHy
OAeEsXqh0hzjDPRGvRGvJy7pAAIjGfQQ1VR9pRL2K7WzO5Sn27IiWC0GM8IO26og
B3Y+f0RfM8l6wHEkRRWm1Lskjdd4Si/xY/KZAumKzILYatY40ZVCCufxtbssE90w
rEed3eTfiitj1H1yFSFbimg2TvwChkcEUFNURnWm4Eag6Z3V7T51ZkC5y2ghfNbx
BmKrcrEmNaVqxuWDO5MFoJks7VpEZg7kvRJVovfhLNJ0NtF+9s36P49U6rt2SSrq
Ff0tHRr4/bF+2stgDUF3o2fgJKt97ETGPTJnxoGkytBZRxQq21Qtah/yxzYTMJxY
Zhi0zzyn47o7L0x7cD98xt3DRWsI9dYS5TKbAv/Qn7EzCvSFD+bEVvMJt8oxF0Z8
xOYYkwBDX36epu5LfHXz2DVJCaeZadltbSNFhj6j1BtiFIvvbso7+A4393SzyMuk
qNRP+i6YuQz2jUPtyzbhaEj/XHNpByCCfyrwKiDtAnNQG3QMeN1UZexMij46PpIV
aT4g7+EPMYsPUijDGhXR6BXpwEOX/P84L2jAm4naC5HTur7icBkmB3owmFkd4rNL
0ikqi+bTndRvnf48B5nd7VD0MWOhxl5YPAfNHF3OFRmKMgxUCNf/nODHR/xt9jpK
7cXi96frizQUNmBJQZDGeE92KpLu+kfwQEHRPCjBQHwVmZc1nPhuhJrqMomzHqA5
qhFyaGif9yDS5936VyWk/5U7DANZScy66eTtFPAgpwAI4i4rVfqgZrxhb07zYR6w
9yokg35Up9AjLIu3VsE/+XPo3x+qtsH8vxq69YK53jmNF7h3hO5nAgdlWoaUXmt8
2i1r3Pys8KMN7X2QwkbhpLP9DSQOu+3XjtvI6RecDNZsOtwe9/2YfiZZDj1aN6B7
MouUOsWXzFaUB6are86dJDdpp0dB4ed1CX0kSQIKTCFS3jVTM5XEbsjjEKivO5xV
o9chfL3HVA4SqpJz/fl/G8SdOlVPP0zsbcNvI11he4K6jRGnga2SnGmskn2AV85s
668/p06LVNwNvD8bZ/yH1hoEF2nHGcywD+MEam3vhGVTConMxOxee4VdC4+JdjNq
Ez/9UZRG8X3OjIrmOl74VyqOLH05HlK1UyOUxe/biIdYLSzN4A21c1zf76lwb+X8
zCr1xckAfYxXbOtrtvFRBNpn28oVQSb+x4Z8MClS9r0Y9+456mlANhrvUaUnY0aR
2AsXktKLv0GsG9MXFklntIfU+TWITU+A3DxRHaz3HUL6s4Tyh+jycb3FFuDTzreT
yyiO2Pf53uoI8Nn6Sb669HDKtgtjuJrjaM01GIujor0/PFTZW45w2YcnTzmkXBzB
uywVmX7ajAPwBzbhpFLeJ6sRcidp2FcXdxFyB1Iwa7UzM+Y6gtHjsPPPEfenMqrW
dVszo7/tx5RfDXB7rBMFZqVTJ/GOTo0AwGdDeZZJI6WeTbweWQaBp+NkHxaC6bE0
LdjIQUpDdryFXcOtxqD9MsnefYzsae5sByMiiOFwmyM6TBZ8b1dd+ISu720QUEyW
5LSyB+aSlMdfL1JFSxhVG7Y0WSUQpD2F8b9sPXG9x6F0Ku/O+tNaCtwVCYLhrKMW
+XtkKox4LpKN77Xa7X4iFVk7EQy9IzEnrKdzi8LEEoIgIN2r6sxyrBC1w08sfWra
jik19VkFDoZE4YJ+SFizSAGYi23OIA7fHiCXYTmdbFdLd+yTxA07QTO1rbidN5GM
euxpCRd39kcFGttvGKEm6RoAg5w+OPLm4h2WmTamxqAEUpjOEwGejGRWJEwO/sR5
hrv95htlpJiW5aelLpTAEjYb20ha6iTjSn0/sNH2GombpNYO5dnogtfu9NTcjruC
fM6D5D5KmFz+s4K4m8HxIs2aGJiWTHJImd5hHUhWljCnM5rLcmtQ2t2KgX35oM4v
tG7hPSafzP4UYFQLgWKrYiwGt+8X+Xw/9vAcERIO4z8DOxgHJpbLJlsHlZZMg1SO
8whkmgLabiiTWicOc6NHBXU2Gd7d+7XWbEYGjE6/Ad26pq4KI3ynaFj4UwPcALD8
KH7BLPhsR31fCvuj3fiVdN4qmZrBt7n2jxS2+JxWVdAKIQh6gaRnKwTS1JKhKXyS
sAx1oGv5Zg0N8rss/eswmaML9Xg1+lik9PJj4V1oxRqRXVIepOxPD5x6j1Ya/MbI
zEnHgUz4jXrr/y8VoqDH8uCGOddQXq4N1h3Mz7H7nflDSwQHZtCIGI42mhygWY6w
OsyAQlK0b4T0NfTZ/1jS8wgBmkDTCxS6cEaKGP3wMDgS9+uYGoI0JC0eLDJsGQvM
69erYd0BL4+KMKcr2crbzfvtJ+arw9ECSeEcScHr8+PH83fxPtsGUtSQMDeAs+Zg
8pFMcDruAJyPZrXHv1Ay6bmfX4DG+TLR78dsKnf9FlfS2Pi6pJNSUoAubg+D+MAc
mu1WzZUE7/1CLnP72ovvCjixfOrulxbEw0McEtsKZOjo//JwTXBYtxjTT5AzMMG8
KNapXU9oj5jWJL/PTkhagcN94A3bJCRDUKrrpB25aew5g9VtJ2JGk2PYlb7PX5IX
BdZLT4yDBdJdXkjTApt9u6Vmoxm2U8hUFO/OcU6oLh8wMw34CoGXfGZcgEur+oQS
HerIj6yn5uyApnjQ4QUHJ0oseh66dwzugn7Zt7OOYM/lJYyp0P+IdJP+L+7MCLhw
BssNuabwGSb5rzaYkY8rOiLyM3E8tgtQqjy6DGbHbmytTF+Fk0mPHqNOW3a16yQV
caoQirT1Ci7ApQjCaDYFVh0C9waoG1QUj//XyjUJnRWghZ1AYf5wyT9BCSbmlCI2
PnZpYUYhQJDq2pEwcK03445FgeUTKbnb2r0PTPFFkBrnK6QdVNLiqkqIpS/oMQ9f
3ET1w+PbJvCBRFUFnfLO54CRNT8EAwCWS9UP2uGJmSaXwfp+ALFnTJ+iTy2/o/m4
79D6sI4MTewL8B648Me8ZUeY/I1vLbHhqWzxTF6jWww5nyT/TBii0tWHCeP8qfLo
BywBnZ/v8L0WgOWBJYN5caTFDBe4FiUHFWb09kClXe2K6hoX/v7Gm0dx+Pig81TM
184v+2thu5411fztHgUbojYcpq+xhxo9Jxj9qjLFTB2AZQoKupGOGKUhDc4TUkVH
ExDeIpMoL9dXI1Hl/OTGGdKQVjtEHN0dvwKWdHatO/YUGDMauRkdHf7/8ZQjOILs
5a7p384vv/3MdrgaB/MT1GTJyKC6XLF/iCFFdawpr/3auglHd1MRcNknJG4Z4Spg
jJmS+gxwlTLxkKVLU2Nfw4tTuy5q4zchZ6ok/3XVRHJIcz/4ZOq3S8NSfFMpbhBn
v1K9+TJU189ixjJMD+zy9qohTf5HYa/+8gX75FdQxMEOGkf779f5e9gODjryVvYc
rYRz56X9irT2+vUVBaRb2yJ8+rl1y7UK6i+HiweODeMb2BZwI5nOBfe4URGC2PoZ
GSlybcLkAIGarFtYw8/xwlmvz/HblImkDw8gt1CDM9lWG7qv0Ryj7k+gBcFcmpKK
IA6F6AR6VRrjcNiIZ1Dizdc+XA0mwEWlDr9/FmSRJpBEBM5DGHn/uMNr7KJ844k8
qCaGLLSXkPx5kuAhNi1Z9DQWbPvhbUwMnB8aN9HAxzaHDzdMOZco6HiCRM9mF0Mu
wmWdK8VVRXDzJQNMhocMLHWbzxCzKt0yrBFoemGC93JPfKsz8x8PofIMfBAVrMAh
AyVlP/uQuHwPPcxepawW93Uc8XvTOYUm1popYiU7hwZKsFaMSTrlf6xqGn3V7O8u
R7eVBCGpn0Q9GRlZ+AROftkLIYYyhUn29DGItGwoVZIRqkswpgLyKkP4r7M5vZz7
V1vQRT1tKKphKr2aJJxerjUY00OPO2Rmuul6kL6b1h+mFNUerQDSs1aauTO8X56/
z3xJ+lma86SpEvWby6zOw+5TPKUQy7ebfmX2dCRyuPWUJciGK+TN8yLmv2gBPLT5
AJgLD9SxHL0KchsepdZIhFKt5N+WpaIdUW+h/F8TDO5pUZpUBftkMjJ45hy184Ws
z+NubgCSwuQTaMiGPT3BzdqUtQ6C7tDUicIfDieV1vq6ajiCK16yAhBYL8zGmXbK
K9DdVzf4jPS5MZoGIwawVr7ovPXdmvwDyhlU+GCDHidpjdkoY9vvMnw7xLxF81XY
dOXtFTIDtfHwB1AkUWjkpeumFwaHUooWGspBVdBMe+by9YE/rKStBpdXMzt0pZEN
ae91UrJcaH6GLunvkCAcW9dwYZskmc5zdHLPTq0+Zyd4vpP9aBFw7jcJI8pU1mgj
p/I2fUkRdRp50iNei2xJeiFZYNrEP9zuNf5hRvjwcaiHdSiRdemg+0kQAtDrwmqp
ridC/uRK7aljn6uzl+WcBBgu2CV3ZGHy4PvOF5jPZUeCKCSI9RbNszgdJBzCe1vU
rtbZ5vAjoOziwjpukCGMWLy401F7Gosae2+tnyk67SgpgrUy5xMtH06XB6n+UFvl
yeBhgxwsXznnRZzOdRoep+pkdkx4JXzdBChuXxeMwrzu+Q9rAgwDrIXEEGiztnwx
636E5NkgjO2Vsur87DF8GagSDhNxT/vdGOU0cpiQkntBB+PenLd7OtIuwmXmzc7l
BXJTYGLT6USXxaDEgW9geH5bB+DWqArnKMQh/5/EKkDPCoeHE2DE+TqCr1jXcbDW
ZB2JUiIfeBi41iY/D4yT+qWgXvfmUrWr/YX8upgdD6Sm0Y5YRs2vZpySdsVlMsIA
96ZJ4/tx416hmuyr2NqOD842eOVhEUeaEQXkMsyk0vyPm5Nodrb0FWwUcfagpUp2
U5Zk7hNT9Hmob0BcQ3uYgeI5XHiKRto+5S5VxdgvSIjDmkJMFuyl+fi0ETu8S4ek
FU0o3IHPs/hWsMgr54D4fTRU3AwWjJRMd1RL28MXn0LDfNgCTpQO2xeOyqAxCju+
TC+3NR3At/HprJopWpvPH6/ItJka9h4Wit2+pDGQ+R47bjXtqe/n3FwPHclJKiIb
Hi07pEz8PVSw7crX7iFBZQE99Dygnh1MPhiK2TXuFYgdF95+z6CF+O4+hr188Ng8
jxNM/rN0NNr217VtrhBarKjFN9yEw43S1AYceZqOdcrrMdfBZsapnHkjEYGd05Y8
49uWTzHhHQkkEZ4KDPWPgXiCW7sATS5gikjvwq3yCHETXzTFoFctKMD2Wr0xnRhv
t6U0QIXnQutZplbilepKSFVk5bpFOsq12bTCHashry+n1cty7lNF5/+w/2tL1TBu
gYaIPZXGkBHeO71lBjV6rntQCGE/Bvr6F68ooIF0JCOzXdU2OQ3oU4onojbH++Qy
9Nzb8vc6Z819yfXtqvJF3/e+DahpV5D3aybs8i2ir9RKpX/WhhGcFn0i1r2ysqo9
gxvSGy2BGQQPb4OP3srnRtXn+Ru4WwajpeC3VspvLhniHtaKzSgA3aWyQXSMpETt
2dqrJigbFgtlFoN9T6yOvaZWsgrRTZ29xgTC6hUL2IuDCwLLfKNFQBlhEfjfQU2s
AlBzqnGBQx2ezzGRiiGeAUa7zj0/3qslxfH9xVmk6z+FZpy8V+o36aKxerpY7Y73
sXrlzJ/ZDhUXWr9H5mW4U4kJdGgVTuR7O64jCrmV9D1BgytAa2jLeTvEwHxViTiU
sNPgizleYxSy/s99Z1gPiIWSOtPUHLPOV6z3OsWxGEFqXIJGTcsvlp+/t1hX/mSL
LgkK/B3BdhAcWJmDkk5hmgJPF7oZEGJ8cTA6w42QcLzVGPTzEpkV/f8lbLeAnhSA
I3NE6t2tDfxcTgcQbkdhJu9tBO4EBMFw5s84EgE+Zpk0ghQokw7CAa+ry/CaogJo
6f0bMvcon7fRdi3evSX8scyDE2f0IxCEdQLu9p/9siBYKIIfBhq/wyP+5tkAWIso
8Gv5MzLJ9GYdrd4HJ100EvpoLwSMr0bVWXY69Z66J/BM+RiYMPxKwYhUwFcZD4Id
Mo5jUl8Rb46dcQGsKCV/r+eqo4wiZnZu9h0nm4OPF2V4cxjWAUhccDpnGk4WA7CT
cdZ06Yhe41UK7GCICMVzh2Eco6Wfq1gQ/tdVTJKtvi0/xcptKp9gChKJgSXFbYBO
A9emG6QV2edISrVA87xf3l4nquzXJ6SK4mW7XnXYnQJa9uroyWftt5y/x6KzYHDO
N1l+vZqM9dfuB4Sk3BqGOEg5PjiEXN4AIWD7k/Dc3ie7D54OhHB3H8jTiquZu9Cj
+u8cYIB7eBkesLwWHPDCVFzWigJdyNkV6DvJ3ACdnoXFpkVc4ovyAQp3/fkeS2Gh
Sq+OdaGOesofD+dowGcS7ampiY3R30WL7c4vIqvEw41+g4YZ6xH6sQ3hBBHj3vx9
C0bpgmBbeDS53dOoiKTCmdyLajhN8kI4ri2DC5p4y6dywFw6jqd/wyD7DPwUZfG7
91MTWzY/e1YuY4BbxpJoI7P8GpLQMHfRqWUODVKQEkxMJv4wA41dSkZYhnHQHNQC
WTn2MLvpPtJ0LqO0IYgxUIFejjxt61p+/tilkFDq5WBR8edvXhU803c4quWtme7r
jQnNCeFdhNhwZzY7fVGKqMjUgRR+9wyUs58/mZKKc5kVNfAIMPbBze2h1sXq/rv7
S+PzYkaBFV0The5JcxaYkUs7uMN3oPxbxtQRd0uYG6xLwITAfiRN4ZUBB2GuFNzc
8HO6vqNt9nHs63gjhQmYhrfglk/ym34HNu2lPGbsPd2psSVvs4dvJ+Je56fHSZ5i
VyRehHmR0dpZ41C0XefVpc3qnzyGPm3+ngeqB5TAudi1RxSMMnjyPshv6leSxDbL
uz20pZt3yYAbAVCc8qBEP26G6TTPIyfuZXAKPAmO1xk44xHgqib+XRU6/71wqbot
Q3DZsOsOXjiU0eSgxykxfSZvzW+9IeKmHZMVfLGVvyn2lJuR5J/oMEKw9Oc+BWEK
82EAG10ijmbYikXLi8SaQ9dbCPAz6cVu42CyK1pmvYAPxfrZGkztmONql+pluq0o
Jq4qlOCpOvWsquXUHJBmi+3fSkfy1LCjNw4IU1xfRaCo4GMBEeal1oVtgZwfcy8t
mauLuwOpk8Ixf/GUvKAGVc2Ku7ZBBCrymH4r9G6geOdX7Gpk4AWwDlg/aUgagEUF
vR3CaxKShSR7erTglWTWPsxAvxrFLyyk9XsTYlg8UvX363kD6RncI7obFZn34fFL
HxNPYJqu6QdoVZX+halBF/PH8cdYNwEt7ixvddEwt7Txic/HV6jseXtgvuk0m/FZ
cOrc8Cmo2oCpYElpBpASadinh1TMBfolj1UyOj828hqzFpBRIM0OQZkUnHuIQASr
yALM4dTLDlQUYXTEnHwkhhekip7vpEBx1fcOUFTK+Dk//itCURD7fg1Gh6zFICPI
zdXhHSLP2O3+rtdAptqf/TMQnOEgb83XZob9EpbrhySCiuzvWMl+qZRhw5PiMSGj
eqCwTZeDbzWS0AwhIuMkg7iPo+93Bdi6x3Y5dBsfLFo8J1jG8Q5hnf01ezd96EgW
pog1gz842QwRFbHzdmcCPcNQjGs4k62c1qaqhghEHVFRwvhgo+8YK/Bs/X9M0uvy
dD1J4M4Gyy+nmNXhFc86ItDBrLQyfJ56ojqfpFdlrEdxrBrq3psp44VyP0TCrG3g
4CzN67DJTrUMPNw+whizG9zDQ8M+M16ro/l0YhM75EZL101SgngTQu/7hEsooJ6w
PruUUrDeggIYcoQwl3z5nTC4cW5H0E851+WWzALuoSqfnYoZB2p7K4WGxJlcH7Jb
i1ioDYF6MB1D32wGQVLf9yvX1RUZyeaquoK184qi2hGNYs6T+TMMHUJN+UmAT3do
bshYzavTGntFx8J2a9zXiXrDSqx2kZ/jjyN5bPcw8EjRLyk1c+BwoCyVyRv2aiFo
igV1sn8ScxciNUXnNAWnUCL6fmjnabNmVhym30XfVnRkUoqN9Z+EUqpCDhM88cWl
LBjeIcM7wgUEhVAMZyvxgkhZQR2Nv8Zk3tTCWIoQbTq4xaPjjPPwAgudec040DtD
x7uWXJiZ65seR0FanY2/JwPvFL4GVNsKrRCD/VSf4Ji72vKafFzFA7Gx22rkgt7J
tzAgJnlr6iFTLm2DCaU+y4ygnLErbTYm6eC1FPM5zYYh3ASzVA5CWmRfFeeorhWH
LR3HDWKE1AfrEaehcrDGpkdJEKTFkTF+eEVPXBRzwV3rnKquId6+9OeV73ITEK2A
n7S3qJPYfLX/FkIEQKTjq4jCBXYBzGw1ndEDNYj8hiPauOv9i/V0bZNQhmL9BP/V
FdqjQVDffnxRo9z/OyWtGqL3iPSVEjtlQ6WDdK836whUg93VIaWAGd77oinIrsYY
pwRZa55Qyjp/w84Le6Wg7OXeKW+p/BKnkv/TcX+LRn4iSGAVuhx05dCEDznD5mC9
LdojHdxQFLW58gW3wiVGxZG/5vCtsEuwiX5lhc/y9hKpLEm0n9R8VJQZ7JsWTDe+
KBNveZU/OcITb/estdkQgT0RDmNdjtZwAax7kBN+27ig1JOGvu6OW3jKuc5bkOSF
UYwsrvkaEzKib1FHpDzBqwQqGYrxYU+1v1HE6I0+QYBSVm61lzvt+fMDkzzX78L5
fnY3rBqzfwZ9kpkkcWBa9WRxdO7icMrImT9ohnpnQh/dg5mia/hvW5XbC3WXieid
3ZX05+5znHnNLJOQSJIIMDsQF7uwv6c48pNQEDjuFy6MYeECzXz0YomrZcgsRcoO
yZ0uq2jn8G3T/mp8ZISN6X32U7g1Sl7TYaexnWA8zV0DjSLiWE8Ch2ONb9xQ8rf/
huFFQMOzeKOQy8XAQ76ww/+irejmSG22S/b6f8NPjsr4n6sQ6Y/KWR4bK7ajLO0H
3T4E6TjiPS9gr9yh9eLKTV31Xj2B/qNSRq6j/Wkct2GiPFxe3dy3C7jZtiUmcF+w
cpD5pYnNDmmeKP0Ma+W77SMLCLC1rRo6LywMruhPz1txOYI8rlldVebs0Tr5fvB3
T6sp/xoMLW4lSpUqrfUdXU9ucrm6oDQOpwflR2PyIIjDLsPA4OyjgKQimpyZbVP7
7dixXoL2yLTXCKI5CAV1DRiufxcyg568F09s+rbkXU9YsSU3QsznVZlqIFYohgqY
TKiA1uXma/aep9S4WLWQjNknvB4pkWB6C1NJypWUyFS2x2u+jiL1bpkg9gYw+419
eCjhmZWp48LlunhVgaO1h2qM4gPccyU930w5F9ItyXpulskw846whdWdasFejgK6
nqGen0Lwx016xq91zWn9zIricD6RO9N8yjxDdqCBlEViB//SUfuiZinxtiqX+xR1
F9ElmSa/26i4b9a535yRgyjGLGfOamitxjeqLEl2LZ4F1fGNgM/sQ/fhJ96taImm
h0Z8Ewwf7+j/d+3aGRz4B4E2Vc/x5MTTDDhaxqfy+BX3NVu0G14DwuFa2KNsdTPs
kq9Ecw/PSejwpXZAVI4xQxFJ/nTfdcJm9Y5KNvQelVLxV1GUAei9lVEh0h/1XOYA
6Rhx9Jso0Uc3Y3gQy/xYEyV1yL68zs/JX+Me7LxQXVwXsbOxC64ZvyIHlAqUXIr5
WSg4dMsE8VzghsKzkZBjluugZuR6F4YH+U4G8Gnh8h5Eoa7cjUPnH7GywwIlCB81
eGUChgGaJHZrpfaO3dSwho7hv3KzpRTR8bRnp+3B61LYHriGuJsrQN8QPqN2YVyq
z2seDRILNi/qCdH4sSepNblV44scPHpOLYLbbcErA9oZZGTycoxvze1qtWa1q80N
O1jE9RGv+Q9h7BNmcXmicWWaESuqWisnI86Q5SmjhB4LWZFBTHZINgErA2VJbUAb
08F2YVO1yIm10PyLZYSrhxKZtV+hSPfQ0dyR0tqrdpTRz5YCwEoDkeSKLTaytFrj
nHo6tzb0ik+USih5L6ky8P5f/KoeGFQ4Mjab44vqyVpM/GbgJGHYXTmSVB+2STZr
BxaHtSYDQWBqtI4DecLhutBiJDF6+ztFe3ghMVOO7OUoQauo8xfT0WdFJl35Ra8U
Fofhz6DuAH5wAaRCWwpBygaMOPiobWMAjJ9qrJjDCLGrTZrPYRebxi6B7IQ76cM9
lvkU/2aqXD7gddIJHV5cFXCzVoTqUz9krIIjAZxUSipJUt3rOSSjiZaZN3/Kr20N
FUuJ1T0g/bQZgAy/i7+hBPLlHI/v8GvsK0S5cSaaZA0JGlsX/4Bihg9FkQ1EnLTk
WdsEEisLxxvzG0q9xZA6EfzI+PWkOOB/fExRXgBeFJBPkoBT6jJVFhg6+c4MstUn
7nJMBOGCpx1TydnYjLE19qukI5dxWeKbkoooyhQ2E2Mjd4JqSVxhjoM7QD5W/rXB
yQA3j/3Iyvq5rxd+l+4heKWHcCbRmge8vhMKN9/SunbbBJ9XY0642EY1Bw5q7L7C
uzo6ybWn4CNXXNBKjV2Ebc3JeEupKisoPYBYZWlONmqzDiRQUZ0/rUTCLmyLGgaM
2LLDo8tV0ors65lPTJdKRIH9M94Z7qtCimYBJBEM/keu+cq63LNpJGCyqK2JG6yP
gjeNoKblqdVPL0Vd1kyIHcNINBis7XVUssosCK1x5WIOpaDw81U3TC2CQw7VZzTk
nPXPuIH67vSVeDIyVweNJUx+54Iv5NmJM+JHfjB23d3muXDu1lMeIA0VMB0cv4h9
4gCIqXAw9e4HO5FSZ9vu62eK4Cc6VbbCRi/N3krlw1aaeuu+Xv8waOr+uznTw5EP
21ka8muK9q+UqGB24dJV/5OeJX+s2R6uWrkI+i/C7yFy2/F3UkdYfpIOiTuL7TKh
lbIXZE1UXAtmCihdeAeQPITgeMJ520/bIHw9UpMxwNqcnYmB6f2jebAsjwDL7s16
mbbn4jQAw3ChqhHLGNSg3jLwlP97bEvfShAUhRpgAF623QhI4XT6E9teSHc5pzKM
Ca1pi4eAJgKzq9iLNgEmBJDMfT7Fm0t1t4dSQsNx5TmRrpDc9KhrhtT/UsaWt9Nk
aS1G6V7AGZOHPb5qoYapSp7+1UzCqNYVJgKBHNeiKqJ3hH6jLhjkBNFEpoCfKvxC
U7jn0MK8eG42tbR4jAKbf0EANpdUWqw7xCUSehWN7AzNNxKqJHOdSjgsojrf/fRN
zzY0HyLTz4q3FSuz0nBNcFGCYUY4qcp/z7Qh0pL2afMUZsEHRtngGyFMOj9Alw8c
u+H5fp0Lo+FfhbtRgBbnqGirDgyArxa7QGhnd8yccfksT078rEH01qXjh0zdUjsH
UFIJwT/3assbGXN3hMehiIDJKepRdnM8B9Lo+hTpuCg+oY7Z/2uIZI3JO0wnYi8x
nsLNCQ9JAhKZog+5zOu7qElL8V2VcTp4Wd0f5HMUZMx7/B7j+WKfVJDzLYXqg3kV
nm7iI2CZ76MJcBBPFwNgukmc4U0nTexIY4s4j/Wx8UEuwl3nxFKyE+TPEiwgPOoX
wRdy9WBjk3H3m0j4LcVGgPkUtFDILbnb73Q0B54ScCSH6SAzA0n+d7EP43uhtzvi
FhMa1silpud/jR2m3OcXaxiC8IddVg977C67Mgxlgki65QiOiNiSerJ2K9YmL7gY
FYlfdxjiORFokSVHUs2DLG4V/kfA7JGQ8CsuNuCFRKYfQsJkZRtpfZeMHsfwuCPg
dKkVJvHrCVLayyVzYTOdxMy78R/+rKjYlRpDCEGiOz+YagGtT0ag+zoIUfSw3xDY
mwlI/0YegW9sOkqwZDfH7seEgRSWf/1QpCLAXlEWLPXtqqNg0GK3Q2DAPd6Bn/Xw
AIymIgTRuQYmMgOjqBL/sNzQSsLNuLKnI/2tf4KdLxCYhZ1WgpSnN3tzs3HCCbxl
4OHStRKaSasFuGmVpyw8YdpMF+icOJVnKHPpIFRdOxnq8LIHsFVQa0nW3vhbTaVb
xxCyEGTZNRFCOK+trMoSdCJ/Kvc+ksLnvupmJr4WyqDaVNiZqJfl7UW5Ak0Oc0va
i6RZlq/Iecx689Gzby3W36GxM/XsHlDygGyLcrYbVfapt+P7zrsJYjQXycBeG9uL
FWSIcGigTqkPVONqlrXZbgU+6s2JfPJL6rsda36xfo2X3apzlrsBKuy5AI9nSbIb
9snpOiKJ3+kNhVY/cMbx6R0tbIxMbTEmLHDbxUUxMlPN5rRdKRHI/NzNjTv5aujc
2hBEK/mYdPg/wBP0+viHZxhXMAayjxRVF1FZ9NY3KbTfeRH+fQtNSDdF7hm/Bg6A
pOPX0+GCrqqkgO5Oq6GbYTyr2LBSwMWHOzCiEI122Z5wFuVTokIVR6UqTF5+2f1H
oNJTmhwIt2aMTqfEVQstGZERwlMSFm/nNYwMsQFDFmu/gtrOwyYy9Zi7drVc5ms1
LPWZEWJOs6cXOu+6mk4Y6p9U1mhI/jcfr7GQpBk14QX67pFasjzdVRuVRnAuNiDy
ESAbMqSbObunaSOJBAj7bXy8gYZCbW6PGQS/yVuhvKWjuHZE6f6rlG41IGTGRcqc
qtS69ryxMPUbn9u1a6Krrou0Pfl/OD2Ubml7gC67OmjwKF9ODre2vVTPIKXwNy7F
EE7odItJG36X4BdEf8zz5XURByPWHEOVYn987J0jy3WDlpoI2Qk9ZiSwZNit9zNu
+KkZQlx+PH8Fi12VjI7bG0on4M4MTXoU6gErLMhVb7SxZlkTL1Ql9GQGQQbpftyV
yZA2XmfE0+2P48xIO3dR6ndlR6pB7dYXBCnpOh4lpkghUMrgI87FxPB75OgWvMQp
bgu5JdU/NR0EqM0iJigTWBdMmPYDqREw38VRQd02AseTxzFcIkYjMIBHiGpDUGkE
w0F7oAmXfd5DFTjbjokJe9HYdVwsj5Xit4WL/aF1nt0XQsDSyAPD3F0nRklNJiNk
kIP5Wj8vIJjgGT1xzs868JQhmoHs0eqavZ2EgSKH8TpucmP1K4xHzswk/Yzf6Itn
hBWM9maJE5nzF+LKk8Fu1l7tQ8DJo5je7QXIVASI6LRCe9osyIEyXMfIbTCk7meY
5hMcI3HSnj7AnXATo+eGrK45+4fkwdEhtGz2Qa6tz83+AdJU4rFfrUejO5qJJfeg
q9rusc1ImaegTTq7K9jZqrc8qElh4M7VDY7uVqeTOgbCkOFReyU0naCOZXLRBcbq
L225bXjXUiD9gUpW1mwg+U12q11XjVB+bXfLKaO6Gy5y6XZ9A7XhnTFW3jLsjTtA
GXXfcXVHTNXwenjT79A2fjqO+gZ5d8NBRBKvvNFJh2oRDOZfWXuOV3XU7J4nZlso
WFlH7VfXDwvAsULqBpesBdl3LQkEsxrTzdZjJcBN/SsvpyBousHNpsbeP5SvrqhP
qUGdWX/S0LFC2rhNdsA5Q5TPdzHDMHuIhuykJaeHy7MimOpa8lgz5i0MS0JDs0iw
phOIWcXrbEcB1LtOJWAJJFmYNjZPer5f0AcmmJ74i6KMGmtkExEHiMZotYQCz0Zq
vT2ofQ6PtL/qk1xDnKVbwMV9Ob3Tm+j6RUJ5k1QIDsdnGRuav3UsUAlTPxihrUu+
u4hqVos4xCDP5phLY+RpOUe2TgHoyS1LvuMdg3mwYbRhKqyfneX5bLGnQvjJ1QCo
uhO2QOxOjZJD5MmVzY7FWWo5MX4FQWmLantw48Lb8O7/3r4LGqBNIbTLVuHtbO8e
LTuzQNbquwh1xO5DBFszC/PgGbo+g+6dV0Zrhb6BOi32J6ODgRCvkn7LNby11fgX
QaUfIWVNv/N3NeTgRFT8vlMRiCK3RyMywM/aXao1WlZl3yrIpvmyFGa+KRA9Yq/P
7SzDUHN40vUQP/1fQ31+bZ6upe71Uk6qn3gmbLI0EFT9HuJOgbPx8+cqnO31WnU6
Q8ezVL0Uf2LBp3AVgtPrASRIob/ICCwy5Y64PEinxnAlAv79wqejNpjzmnVlIYci
dL3clAG3PeJ7n2bzKXE/L63mAuNoBzgfJViH1W1pDFb/embpJTlGRTG55J0dymxx
MeovzRrJUeY2dpUetHiG5UrGhrJGkMpMcRzkPxTTED1O1+iB3rWnk5r8HBG5YoKc
xASCALuJtqIN2OHFm9lKDwFKb6460DXbpjWdjVrtvWnDW0/mlWhRl7C1L3tnmhhl
/Jk+KvbSzNAqNBP7Ff5Wtmtd05R5Y9zXFYkNH/Z+bq92frTx88caS5EhWdj1vPkL
f2ziAwAxItrbaaFoJpcAqmDp/TzyR/QE3R3ewIYnq6pMWfTE6P+xYXy4147jP/xT
6uOnO2stkufK8a+oKUxtpywDB46ufqIEGvbHaCNwdD7z4IVJr3jN8lrBlsRNML7Y
iOz1NQYaDvV23lgGTpWcoMBiOEwnvWb6psCb/8xfCnMpsPQU+KuaV9i7eg2jVdF1
z8Pxm3x4PQV9kn+TekmUlXnqtp6qkWmn+5i3FPcczov1s6j4v55EDKGtySRGAqcO
6OTEHKlv8YcM2dxpsdRtPxdP5ytdwT0wa7gxWAw9qiKtTgh8m+RPgW0g7QavbgYE
WqBA2xgv/egudl0sP57jlZfTvhBLWTlBn4tS3LNsaR16iiyevfkX1H9TsSSTV5FO
gVL75/uuUf9RpIgGfWXReyKImi2nm6rPkJJNVKnZUWkzTtmKtW6EdC9FmuZah6Pd
NeNQp69lR/i7+lxAJ7tJIVw+ll+9S/xZ3vaifjkEEt4Uwb9RJ+EXXUWeLcyGLJn7
GoaHz7ekD93wIw0ekGvuEI/SRVZjpTxrpx2lZH0Zd1R/gl4u+zr0zRlJj35ly2vh
CLv/Ht/DHLFM3RGdK2MEh0hHUCvO2DuHVmPachCTHwKpsnCaXq/KTd2oRUkGxl5K
Q8csNp5KUznTADjmNzfny7YOYXc3zbo3/8G2IQZSg8toauvZ7t/HyOJszTjmbWjU
ssxX+xnWnQONzua1OifWUQqKMuelo87bN04ZAPKSXz9N9NuPlqlvTXqxDCar3wPs
nt5ub64AKFgQ/uzpkgY2a/MTLXJ4gqqtP7YLg5Dsus/pH+49Q2btkfQ6QvTsXCfH
RKHwWoEXu7zu1bf9ul4aCMGDMIEC4U1XHJe0I4GXvu1c/3XKpwMl/4glfl7Q3Vh1
fj6DSNysDATeATuPMMjCyIYF9ZhraXW0RLEvp7hDvpm3z1hnDCyBSGe+OJLXqKlf
sKrzwaIOg2cyu0ueERc3BnGt9Lb3NjRzkUspexOLxmgCSHtLm6mOrG5vyw51/yIr
UK1jCQ+z4pI9hqz0v683X4m3MVWTxjrToNk2AVgbU8G0Bk+6mJwhHyjTfetwq0wV
QyVimHytvVg1pDR640KTPb0eHj7HYEhL5/UGsgg75y2JwRSHtrBBEqyzhBymOaBw
kOyrkIL57w/VPnFFu38GDtbP9bcjK/wlYH2nAXWZQCcQK3Jx3ILBKtlTiJvVtaVE
74KzIY+DJawqOzFSpY7+9JPc4o5bfPngNb+Gl22Kn5o3NXMDFY58D3ZuE08YflyA
8wokjvtud5NtiJfcwR7Ka0Em44XbZMMl28gCsUmKYZr8kyfhmsb5mXx61I1YeuXh
uFV0sUNS8z5MzkhH88vdjvjjdPljFFVUZEYDyZS0CNq13GzM+64YIAw94LxNPDQr
1wEkOxMYSxZzN+EhUaF8EWUkjMKfPZxgcRLfFavD05OWdDFB8V29YcFARlzkJuiM
2LS03rVdckf2iRAJ5cnBmuL+Yr/9ZvoJisZfHjRl5Td9t9FexdndoUMQ5FA4+/Bm
HYDQKverGj9qirUjS5I8QmVXSpCCe9yCj6Jt5xt5FBsu1CJEhUPXPzuU/5l0CZ4D
FyOFbLCBBA6V1XeDGnaZmJdysOQFXKH8ztrAm5HUYVoASJwU1qDYPMr/VlP9sThQ
xz9pgQDn8iX4wsCmj+TENlIFU18FtBijEXMSZc8QqMAlNyX8/LPx0WTGB4w4/hfj
MTQ5ilv837zwoxwWexpr8Sds4g1DGthko+utn8cZvdtZhHF3AOINy+OPtpf3lhID
r/MjvTyz1Kb0gUaSGvnrFaQljVNWYzvDCPxL3sBD9hwct0t2138xtD2vIkhJfP0e
oiCKhIhwrg7GnqBPihIhXaAsc9Yi7bYC0Qdc1mwD3HgeIHP7v3NxqP7vxb17PW8Y
UgIUEdF1iCw8+lTOiPHAEZgWtyV19rh1b4ep0YldQMD/Fw9NJJ8miftomOZvhtQ6
8Rq0o/ACil2QCI2RhYPPE3vt1/vyVLPnKXWzrwv3vHx2JkXe5Qmx8x6YNzNDlpFQ
1+nnYJsLaniqoP7i60RaqMbD7Ea73M7z1+wMJ/wD1vQXj8FcxqeywJlxsCs6pBve
8DiOH0lKOukmcG2LfiXKB7Uyea/Kgt2xGk0g/oOrfyE8A5VqKoa/8ihFsNV0LCAV
HFLBgbdOoKwsTXdW+z3TN/nj/V7ETnWye4Uet0H6WZ8OpySPE+AGu2AugfN3rMSL
9MsV6UejFIDzfqk6y/m7JYc/L4+t2U0h09j47llDJQGU1UTJtBoYReTkSoRxphxj
6VcJEpXyN8Yf0P+LPMGfD/r85r6iuYNCxgMqWfBRjWUghb9AOhAYyI6cpdORc8sA
T+r5SD1NL2+l7bC1tomnnuoTXYZs6J5WEHqXWR9TgK3AvGN0ijoEmDelKDHJXdtO
x2J5x7xyt3MV+tvi+juUHIZgAKBYjGFXih4Lp2F4QVsSS0SlA3xsqTg4qzmvjH/1
BQAJhItqLOTltLwRs0vOfGR0+sxisp+O3nqpCoRssJWw+OGwIag2CkwW1R4twI6B
mM2vYKrJHKJg2zCGbYW+oFvHAspPg85UIJMuMIiagjhP19PnbkOgSPCv6Up4/E7c
pwMrTtgcmFONqDl2GxnWnOK9kfiIftW0OGSheIR44v7qI9F80/swwLwLFtkxBa7O
22zTKxBnmBh4uJNoXH31nsAOKHy35Lq89WXFMVhK5nk2xlpLTLAe+6noN32yGU/q
MZ9VjZKZGH48ZD7MQXK6pzKGPwXzXSQmDTVMAYTnF3lAsMYDis/bpcXMkx6vNyih
bjNg/j/12at9+ynZfRP6vWUmV7Zyg1lY6g4pD8s6jJfmRAnMX0sZcaNksgX/O4hs
TEUlRnAAYkAjqbcLIXQd6BmHMFQtssWrpGOe0PMfWtuW9I9UmLuH1SBFImgpawpH
P795zZQnPxXW9JW7J7fYSQjeGA2/wYV340bRDmjMXW8dtYBc2bdygTIQWmmQTY88
giSreuWoqH/UIzFRsThm02g9l76Ry/Lbq+KwxeaN3EK5Xzt3MIRKBtTufANL+R/Z
IpoOvNfWk3h1rU7hGV1qPaCCaMEsad/a3bxaS8DNPnuTgleUGPT3GOQTYOz/Nexd
vEq1ordFljx5O1wmvq0rOoSX+FcWHQvhJbusp1wcIuojo7WNUzjnTeoC1b2xADMC
LWlLyTBa0af8l5eDJENB9pjoA37zlpNAkKInzVTmSKO9DKB4E0zDjYOsD89eqrKV
qGb6/JeO1u6jMNk4pqdlVcIDcyww//gH4gx5VlQJAY0EN+nTei8I5GxXx5GSQ9i+
z6VArHV/p8dGEYBa2B+gvKJzrXnJnxCt20QGMDt8eve4gQ7/bakRM0DNuV/TH6P0
2miOBn5UQU24IxUwPD6TyjxuPlMPlL4Edm8hETpGcZPs2JitoF9oQWB9mbApE9J5
dD53OaehViBBmtaT59Fxhx2o5J5xexNsuiwrfJAV1dFdaguHt0KIzbaPTvrnXvmA
cW+h2RK8L+Tfk09X035VF5h93FrGaeRpL0ISxKP53DRxl92F5DUimMno6d6Et2hG
UgvZsCTVI69gncjL31sCxfdWmR0JkaCjvOPC55t+XsGSgMBEvHNnNftapn5mLbQ/
/TZ73+CQs1jTIMoOX5T/bIRnFCJuAlipaFsURydExIZWKojTYjrz6dP17sxpVKrb
9cLPVG3e5L/wkkW7x4uJVBA8BRkFUw2dLWeO8lkKUfP1tPhLiidlYE+lh39j3laH
tRL1i6e7a+vT0aHny+JLrZF3Cl82iH3Tp8qUC4wsfILcva10c5nJKK8et2ZPo0mi
2FmwxwyMaBhFx89qKQkC7X7H9vSvhgONd1fHBZxbQaVJP90/p0k9c7RA21F1iASA
xMH4uEq7bIj3dqdvoluiFJVxlH5/YFNwdOnYvo78USKDVRhfLWshhxyb5kgy+Siq
A7/3BI6j9LlJNi8fQwvUXxBfVWAu/3S2DmAT1yG/d7DxjWJVCAzBWr3zCv0pzi4c
J+nV8RYIjvnA0AbAfBg+aEaG83tLKjUeGS0D0k7dg+Pfsh+G4gL8mvNsla/yh8sz
RSq6nqOFokBM2xHJtBefXuPWmxII2BXcOWTZkDtQ1ECllLKm4uvOnx0xHCzWQcNn
l95a7nZwv6IJf4L2YoZ4ebmPuVmmOEnlFjxSmd33BozloWe/xYgrg51s4YlM/BD7
uY6M/i7AAZ0Pk9DaUTVvgN2odtsZF1jVBrER9enRI+rMFEg3qgdsuhe2jGnwIHOD
5jbaB1fQenYlr27zEs26OCJX22vxC+o5e4yr9FZjNT021w2lPAOUs0VgiUgbArht
faCHhUIQY+u/CQNMjQgIMiCAgL1ZBL9ZrYos8xdAih8lV7ByCMi/tmC3GN1h0+Mk
Rek1QDuIwz43kE3OnrYiAhg8TcMz1u1PO3AwD7z8DweRgOt/BMUeDvqo1qmAKCZh
WubTdaPb3C2G4t6Y+SArJn1c2mCbTjdbrWKAvK0xl5vM4HlCU6QqGXEYsoDynxWE
IfNI9liEZtJcstvpeDTnBfYSf6LPWDhJxKReMiUoFbo/sj634K0YM1G6+v+o2YXI
V1cZwefaFeUTSZCJhHUDc3sF+2t58X5ZaQGVMs5bgmXFx3aCP1ZIkhnEhjVQwoAk
KbdJMktPiOf+X3WB4KUIMzAazsiEUcA5z1A3roF1LTvlphDksethOQY4JUj9du+6
s+MzDpggOI/bhKwztYebmHitX0HJt8yMgWc29YDZZPVHUWVO5ZosHOYHwbdP2ULH
OEUfQCIYFKdO/LXRm0h1bXzFzEbV4QIHi+cdKlq0xPYm4u4GOGJJAGlhGGnL+WOw
rxh4Tjx8eeItDfR9NGLMoVp/gFVgGf6MNPih05sZoIeLVFfVdSlx/9WYz6Qmopwy
kedbqjp56EGdc/Z/k6J45Ky9eTQYevVuysGc9H6j/tLMiBeSL52X8IituWh7mfq7
MOf3NFDnxhm2FCVpHwiT6iNKVR/2fv0jKLmYRXUWHVuCZoTYL/mroudyfzkzU6JJ
L7w+Qd5K+lZ+VfI8Af47UT6LTUInCtp/l7MR4IKDDixHickvN+NceFSAeG2xjnMw
5faDB9JDi/xf3MKgdAdLSbO5wKlHbmpCVEa6EerTc8nrFPUHcIWPn68yJD1UsvzR
Y2C9zVsn2Ez0dtVqNYAMPxDLJgLo3SnkbFYuri9R5mLnVffqSLtoyx8ETVVP89SL
u8gFtAWbfh5fMedphqbQk57JmZbCJQazh8jrjvpb3A64J1FN5iUdkOIETk1QxUys
1tWEPuD0J/9jG9DkD+a+yKSECm/plSd8RAMUdzHyfvaL4+7rJ7yVhYkh/CrUziBd
b0868z/SIpfN6am1aH4NhbrA2pRAcJjqyhGIYrVLfZ8wEz/VF2ybSacd5ERy4E+S
y/ZZNYp+F33Z9BDp3YcLq6wT9PBsPkPceXDT/BEiLEJ1fHUjlIijdX95JvI5Ay/k
xBqwWlMHu3vqG9XDgm4ki0q6rWREsbUUzZDTWyzBcK9jDNxj6wvSf8oyZD73bBDE
QEht+6ttap5/tGoDhswhRg6H1Qj8B5pKizP7yU4/D5hkdAGirEtu1Y3IbP1+H/Yc
KzicDXubD+9949VvOuDbRo57MJyoOhle/qO+KSnYbezRor6Q3vrpFWtayJpDJfmT
FQ6Yd/RpsND4AVKXDRLv6Ea1u/fKLJmQ9+vEZIdirYTSYo3VBuueCkecbtwjGNe7
Gl0DYX3uu6V0QycRGPMd3bZpTtFpEWqLmpXO7pJe/L0JDefRru/7uQlsfH7DK3UM
xmXiQq6HKPxpBvOJUpGU6FyR6AV1jBRqPEgZ14wpqGYRBH5BvQXMovXMgnYOUvgd
Si7Yb67RqKVcimAVDHTEAzpSlYtM06jPw6Ce8lhgbSw9XGTgsnPpy34FV1Bg/DWt
mo36pEvTz6Z/dw0/OjYu3m1656Yaze/K+li0xIRei5aSZV9JuKMFmJr5/QCUJEvD
+gL9SeRCVqctbMJmMJIQFVI613+il9UdiJb7ZpOD0H65CFtK6N/EgFJohijMYshy
neVerXSiRuvI9ZDe0cWhhPVZphWpj3jrsuy6qxlbpGi9v92GC+FQ+J8IwF9A5ZrG
U0q1lrKc95mu1cOzgNzJQ2GqT7yWBCRdK7PtIvXO589RZe50c224X920z3Z3dBGK
FE7198qZ5RZZCa9xu3d9UNCLf5IIByTmTJ3vTf2f3d1ne2UP8QnHVFpSv0JcJ7xn
hg9y/WA+eR3+on+w0wiW0/H/LY46CgM5mvMPXUGzmSXmERe0BENnGmaHMFl9t553
Nbj6iSeqYAsBTHFDzYMsl0qQvvyH6pwX5PWnz/n3jZscQ3JgBuNIHddOv2zGDmIs
54kbLrfBTITma7PdYB3eT/UbGOPkUGtWClNXI2PtW+U6WYKwcosyrrYp6uAcfx3Y
tlvxpjmRmiyL025NhE4t7edufUYaIC8Gs3I/TbS5ATMIOKULEmO+ku1oZuu58aXc
yd5rJ8PNc7BGZUAsed0998Dy6avhutIsoJt5U9PHL1c35M7J2Hyh3WELAxluOfYE
BTTnuC8xHDW5/JZJ2Fiw9LePQB5ylq1GHdtU0M3r5MA6qK59bxwHLSHnOKOlsDwb
vAgq1xzTuUM3Oig9JZxzKKmxp8ZnWnB3uC/KmqSP/x06DID+fh79Cmip44Nmgauq
b9DMkAAPuvx7JPWkd9QXD3osgOPnVYiXiejUkDbNVGAraISXAuToM0ORsDdBOQyi
soTyFCJZTtNuT9k4Vlox4hAjD3jQMxTKgjlf10e+Ta4QZSHnf2A3qvD3XwY9sxY6
i/DFTUP11E5B4X0fIuMTZSzKct+xvIeSBV2HU+gBDsX8SwN7KXqqh8TtiZ3tu6Xj
e3P4Sns4ApQcvvj4dn0gOx9bQ4OTa8LG8ldnu7oneAZJh2cGOqxCmezUZ3sxqM+B
/8T14S7cdI366d+e3MxCFzgIPFuYoNGV3oWVJkaqcN6mmb28MsuIY2IrIStt/5IP
xgh8DIxzumEtZuXRJg6asTsL0quhLdDHNjOfjC4/Jl/Y7vZosEsLiDcE27mnezNX
jmdcXtsdNZ9Le4FKKYQQq4w54HKFNR8u8n3x1fX2kkFhZjU0DYvAhFoVSRKJKoyy
0K76J2qzIo/fK9oOHuei96IhVs78JQY7ShJKYsLMjJ2bsvOBKLsf9R0DtDJwRn17
Y7nSYGEt13suxiSNAB7zag5olvrokCcSNzhukZbEn9LwtXOPFuMzHkwcMQrSoVjy
jF3MgOmiKfCxqJc1maYo5cVlmnkIuCI5LPXoc18mREXfVjMfeQNwKRwMZJJb278M
pmcze7WHjepQToSPnHNm2wpn3MUAosYKSRBhrwB9xpMIh1+WODca2S8Byv+jjza7
u5ual2bUQdK1drLpnVnhaSlrlHDm5iRRI6YN0ENyplBpONiO9fsPqRMsF3An4mTX
dhtobIsP6Yy6s/GvqHv0V4vq+raGWVMr6G0O20reTGBXzz+SEBRWK/U8E8dDrAM3
Puj3vhRtCyQnDIJ/s9wtQ8HqkOjPinUMBrj6hJk99eADEd2BTzBPrxrS+8AM46j2
pLvifIciGFGWgWBRNj/RxP90DjhUEfepcilSsYwoDTBQU9tp577K9FQAcGESOg/O
Dd8Jikqlp00fsJ5TfncIQit+CYHBzsCLmyrED/b+sDTMz8apCwqH8ydeTX998Dep
UGdo7qRRVlRVe5GuvVPk76XpdRD5yqdT8gxXsbzLQ5sr4Wk9+6oR4Oyqwz5Sk7Yg
ORW+mzkRidop/qKJB0Z3aqnAMHcUMn96Y2hM2/ikyrgcN1BP9bnmtJup8LbF8c1o
001WgIawz81zZzldUJE28lqs96G5f1+SvxS3Z8mZ4tHowN0PYtySkDoWJX1ZXlyj
xP3dRIEoU0htScuPVwA48h0AejOXlqRvpb0SUcuIbFJ6cunaq/DiB8CJhv7UfW52
ZgdGoA0rX1FKDZ9wW70EoMjCdZSrFSdkSLlPtnkO56u7k0wkSwsEu1NOyE8CU20G
vxBpLPY4TN5FN6bq8vlT9XrQ8bYTIyfrkau8Qd+7xBuPOkft4WgLakhui3YqUQO0
n/fs9Y2c3OSXx8tG2gVn+sLesOKU68qi4oX14IKzLPkvZ9TquZjIMjXPdxVkBOfM
2RVEv/h3l94fQ6Sq/zHLJGtocK4TgY45FMKKPMXv9ssjEQLy+7ZDfZ4USWi2OsfE
fCRH9auNOpvRbrLlRjF01dtrWSl+M0ZQnDtjUmeG1zjiHE2ATu3IRPsHcyMMAn38
AtgEDJLXuzCGqZ6Qa59eypTwrgpH33U2Wfp8z2QF7HpMZ/YHjgi9TmoLm+FyBzNT
afAL5OeBe6ERC71pWsm2oWWZKUGGRvEV1guAXmrmemndNG+4sNGzn0vXZjzsmx6L
J6yqFLaU2ikF4PeAnMJ6n8YUV4pcfVtP039q/owqnBFWUjXbYlw4WSq6gaGKzWfi
pT+TrlSX169RhBOzDgRJ/hPpg1chOAIMbwtcQEL19n5EZYNBclhmwg8wc/skEewI
xx7V4RJMVI9PV3nsEMZEGBIDH/SHY2bTNqzD5ke+31aPQw/Tqq8btSoftELJ7GJx
eCBke4IiIa8KDzhow5eDZfOAVXHTJBZxue0R1MSnxUJq4rJi96KMZ26iySh/mBLd
nWu+u9x0fi1TTKRsbeQVBqHlgR9wuo5Up6PVIqZsd4JCILVe2ZTpRR/Z3FPHfqxP
Ar/D6wJ/9wDKcL7Um69TSUZ4sjB3W9z2KF6cJfnhPcvJ3BuoQ+rUNpz0zDa96Nb+
S85oaXW/uYXRzd6MsqGrXzGhJmo1P3G5/bg3TAntOckY5jqkFeNzf/9NCIbebAu3
3ixPtYRnNi6zvSCGX/E1VW3S39G/eBpb5vSFs02rRJkJ+gW+zHTiS3TbsN/FmIyl
OIpm4WW6FSpPUDllY8D/pD3NLyV1N8YYS1rmhsiPPzzLkBsTYeQ/2HH5BlWR4kR8
Z3IUG+xNc4WWtCRsxthDecxZUAWrKHX0vqbaoB7eAsWl1nDHmmbMpz1lroAPj5Mc
whMPz1C1981QSy2nwiCxRvl84CtpwEVFPi8My1h06S13y8sp739fUgieIN94vFrH
6SKPpJuPHjLBa9BwtmZ7heImKuxEErxOBOhsU7IrYdEpBaBXknSZomzoq76ZDw+F
t4No7tx5kR7spBHsz/kjn+pe2pvaA+cLSQXGTTVrdllQ6Oc04X5PDFCxAcK4ehbw
53aIC3GJUDloR76rxOx1SLEzzFVXXONdrwCh0xIEWF83tiuj/ohKdQcV11+zU8wi
Diu4+orY528IGv5oQaAFzBExx8P194FRscIPAUr+1BuGPc/xQVmmouuaT9NzvG3q
8BGJdZi2x/GmYu24RPjtprOdhhSB+FClcZu1vx5jolgbkmxkIRi46nKpTpu16TI7
5wPCP+Mzz9rtxiCJhv86vfGy1gKrDrN+oZ4M0oawwh63PJPzPg8MFNZ7T0ghTLQF
xAqUdnWqHaeMWsKQMhYKzX75w57h888eYcffG4X+518oj4rKjKOidkjgpLWOcOA9
y0S6mgG3kamAKWqsHUu1BC3BdUH9pPP/tlLfbcsFU7V0XPoz2h48Mit16oOOyCGO
0UANM05GKlB/L+zeSOhXXrjPPp39RyURzIeU+0nbk8BKJnAr4/CEekzoHCP/FAaZ
MQg72KYymTnN9UDHJEsahm68thczfditgLRtnLNtcONXbX5ZoS+f5PXB/7aqN1x7
ZOKmWB/Cxz/AHZBT+T6NXOWubTfyv66mAVNw2LNKtKTL9Lqx8GoIHVBFSFwckxrw
3lqm38SvpmjD0ygHZJLQnj3CViQW+yINX5Z+D4YJOoXRdmqeV9rJjXmAg9uihlCm
53DlHA5GZBUVU5tChotKIw/fLzGGEBv0venRrRZX4Kf5ZIY8quEIHmzHo80VBGKh
hjiVa1kCei9swIA7W9vvOfVT5xjW6LzaARHcnudwFsOo2a2zR9NNJLLNPlSPZmD8
GMVQunNkqaC/hd78D+iogEBVtCmRX09EJYreBgcfpHqzw78istN+6EL4i3XTV/Mw
mGD9MXUSWvQs8LcOXNPmHhJwYcRY3wUM3cOJuwJRbVIMYcLgwaIJwCsMAdla9tC9
2hUm7+ieW/cIWPAARBEHaSrfoaKcFoRY8z9s6STbGevlIbgAORxONXNncGe5nOQT
Y18e4vubxG4B3DUCFwoZZUvFIW/YClFa2IYmV9K4/FgmPwEqCcdZ3oy9XmgODVDd
PcnqPfq2uvVvByvBbwgsqL3ya70oAK9amBtfYIQOyiRiEi0+yc3Qg05bSL753SBh
a1fDiJwoYSGh9BvRQXyh7hWbeYQbz0FLq/FqwsESMjGyo95/X+xPiaNS1GHR1dQF
iHrGXiSEc1DrpymclUu3PXJE/MAPscjDLJTU1dlqVam9QyWIB6jlI7DDebJx03Sc
/wjILbw/o5z420XiGhtqnv2XDuqBIq69SWLUV1uT445B3shA2C8qdz8vpXmlw43x
VcVHK3+/sJa3lbQFH5VRCffNX+4VE0TsIMq01Mmb7A6gp0GC+dVgYiarxE+o218q
N/Pc4x1EvT3Ta9loss9GG5RzxSxJSsXKWMbESrDC3mfDfeQn8hB6XKKDQiY1Hx9G
rG96Av6qqTUg9A6JxZ1d0e+E6xQd6ZYPnl+8wPNxBuQKFt0veWbVBAc4h1bZj+Mz
dm7y0sOo4MTEEVnCdbSVQ3ZxAJqRaBPTk7H/V3DkT4emUXnO04ASwdGlT0kdPu2M
GzGs/ACgqJqwToIsKbvCefCVIg4ABCV4uxXy/SbfHFsnGZcCVxUO7yVqM5dqe23S
muhEAUIMgW51bHFHtir/3nmrrFIUFIKdKNX34bl21p1E1UynJRJvVdlMqBwIdL6i
hXPcwTY9IYK2ptlXve8pqlk6dktbhXZRBm+8nSyQGJ6jfqV//AIUSmrQMvhQXbZ0
S8nsO46sC1WMLEGVem9gqcrdVvM0NMlX4I1fXVZwdu84KtQhuBjpm3tJoGKNWp6F
+vce6laK1yPuerVnNIV/hBePB8+KwnEWbeh7+pLQv2TlhTaWgrPI4FzV0DzZlJlN
zkkeDe2FqTySM1hY+BF1istUKiX0m4QVR+abHXfJPTixCPrpuQWtt7ygOQidzclm
sEx5uqxzBxoUYecvJ4mkUp6xNYERPiHOEm8oZ0y4pANlPFJDRYM/q+OFkb8eIx+u
AXQjwcu7+52bHxNkh1YaXuP/lis12egJuP+N9/zjpP8x/aKdVAdZOUpC66z7hhkY
MNprMdOHBAABWD4TRDwJMKYgihsXKES4Gf+rqlnxq5nThGhOqYJJo+YF/zfdOK+j
zWGnNHwKHB1PRPLXX7x8FX7uNctiY5xk2j4NsivL61vhycRmk60Lz55NJoECZanL
ZJ+OisRneUSnjIsZc3ZNgvJy8tqHjEH7vlQ3VCkTAecinKqqEqgTfkAnrcMdThS1
SOaUX35rqB32CQmzCzQHRvfhYtzxxUX4gbAcXKt/JSJoiM2grBDH9YKbExUgXflj
w8YUbtR9ioKTexUdpxNZq+u1olyCXX6Ajm/3I20vAjG0+6w5uNPilYUm1bClF7lK
L/wP+rzlx/u8j3c6SZ4rc/TbRCiEt+fjnlrNH/YpXeI/uKz7eMfmoBL8+KT6tFdu
R/X12/JmCbuD4mxJ7J1FQvxY+a7T0HcvYeb0l7POTy0lrxKQ6Ev5KObC9IH6TpkP
BAWWa3kd6zRUmhO5XakJh9d/6+h/ONcDAM1GFplYnZ/dHwfz4JapBbWqNtNq93g1
hXmrfnvDT57Zjd6s8/x2lMlLeo8g2kblf3Sx7Uuz5G79vBcZiHskVOV6cUf6e180
yGVNVlFFGMCVIZ/pJ1hFxMTIYoOC03aSFgAn7jnXa3vdxdl0fcQk/xdxszmZns8Z
IfO2/x3iPeVTJ1I+tSHxEn5epv9St/1IR21aFZVfRU8tmDkaQyRsvUEKYccMC3tN
I//XAyM0+t6rKqKSNC/IVYgeaJnglmY4CpLTdrOyb/tL7qp5hD/lQFDQNfkOWIOB
//KmD7xoMkVojDuQBAHMBJPPj+sBBiMbVm5MmbM8MScz3W5DUkJUYJCgt4rQHw0d
seG2Xux1QnTEK/e8h0vu/E7qeme0KhGQHaFLfF7ofiw6fot4eSOOfpLRnTXHzkl3
f8ceHujbjLfkG74j6f+ssy9HI9hUeUYy97PeFpwlZBO5JnqmE6dofQMSKAY4kHWd
e0q1APzKZK5CceQ1bZ7gCA4J8eX9HzxUrQKZXvfBJkuQoSg939UtdGmPOAITDa/F
V2XIdy73FNNqkjh6pbTDDjNy1q3vHS6bwjfrZY+0rxQNQ8KgaR+T7Edf0XkNZ3fZ
zD9RRyEKq7FSAc7UpyJyZU1v0sVZnGcA4r7ogho8BeXGLZsGOro+jyIoPcs2ZTxu
4Itp93iutiHnoBPcng2rtrIKLzdOmfIBnYSWxi72/FptUxldoDrNJJB2EnFPjVQY
Lbp3/biPBvrgartAEsuyBv7fnJTIiBwAE3gBJGFYx4f0T3X2lC6xkQkUPm23MUtc
6VzbZYvbxXiffaojgwM1nVaPEJjCWYOld2tsgwDmkP0vxiGGyLtPwZo+KS8KOk0q
cH+BVvfGt86c8qx8DhI59bSrK9x7HitBDieo5D+Fc/4TUGxd7lQtPtVmu9YHQFkk
YaoHyENsFLi7E0IFX9pnwYB5r52/oydTg7YVgZCTUR/ew3JpHrJSrrfYlzXaa+Q1
SxB8Tnjbh2DUBw7zER9t945dmHBJa+i6vsEco2wwapHeNYcfFjjW1256p4izYGJ0
edYZGP1z9JU4XS48yuygkbFSFy9SY5EMjPJ7YXiONOIXV2t3Md/x1ivmYe3QfXHX
I8mpEmVmFab5c6Qju4SAEj/ztMQtg1L7G+kNfeYTo293Rwuqaa0JT5qLV+twnDXj
gD+8bqnYIZcjwd/HJSKWV2cvm20E25FlTbSMDrDpQ0+cn44phaNp9AIYU6AEYPP2
2/TuqF3f80CRDlGV2yvdk+Mhk6lWUSON41J5VmZTMB4xgUE+xjzVTwQ5yXvM10Hm
gqrO1Q2nDnmGNEDFAJXfZd2T+6RNz3AHJdg9Z6meLm55Hfs0usxAoU6kbmGm6Bua
AeEn7gjpQQ9pJVyEseqOznISHAdmrBzk5vDc7r65gt7pG/iEX+V8K1NoQWXgeMdn
QSuvTVpJ/Wm++tn4c4pgTND4ipxnsAszFwXSHFthm7fnz2on3d5gInyHW8cULdz1
Nq82s1nA0MD/Q6c0w+emRePb2sqc8D5L2aL6T7H1ZY6QsewngDr5NFi4E9A9dHdl
iSyf62JXCHsAis+nlFA+8LPw44Y79W035orq90tTDXoBRB1G6NXdrKLMYEdOlIn3
EoLVsh2FcqpwuPQmZC3MUqM/uYaPwFl5tPF60c/Mqw/XzN077imdsM8kUqNSUveZ
3792gKHJtOQUfINZEpOaftncXURsK9LTRsII9E3nDUSE7LkK3Dmxx7zPrqZfFZXv
/09OrR02lZMs+IhbCirJiQaaMkQkE/Kx/Y/qzalCinRnmy5VQeGJNKHSukagxmyA
CiUBJgUROMCY92B23UJfIo5Wcs36w0KkZf1hXTC4e5uISQ2Or/oG+XYkfeXWyCSl
Iiq2AIc0n+lqjg9FMVg7BO5a6gyRKrwLFmBIeslYv2hFouuYzJxUnpaBtpN4djW5
iUdqou78OwcH/2eBlISI/ux8+MXxSLrQY1KD8CY6vDDlzOh6XlaujZylMmdcJ/0R
dMcpl/tFQMAgACTPMuEPMvCyjA6TVnG8euHJ8tLjedLKfK4FijhAP1F03MVIBRkO
rE5mfiZAm/OhuB74YbqKLSfzlx4lMTg2crVSr7xn3WMUYeZlMtEdHiLpWshZDfl6
RKKCXnwiZyuBoeNqsHownTgEETIcggRIo2A1fLOvmeDrp46JfT26/9iD+z538xOa
KAyX9YfsKxfM8i6kjMqo8W71DiC+7+2M5GRimFL2Ef9NHeYoQ5LVHul9/UFnXeQK
Azs6hjGXIeZKVXvfil86LMvTWooRtqmperXS+z4tM61dKx+X7tSpLhyWNgqBDF2s
W5yLZ0/LcSr8opsHq1S2O45KBuo8jGUXdWy/LkW6ZRlbm0cO57vjMaDhtyMD2vPD
h+F6m1JjgaCvPy/Aq8um+JCtkXvCMP4HTyrrR3Wge5EtoQCNASnANNYV4Qt2YaTi
j3qdx/qmx7e+VHIcB/hSC+lI25DAa1lmQ0upsIrYv2BSd4j5tdv2xa9hI0DKHZl0
EUdyXo9ZOO4xyKpV0SL6Krd2CjnpUx4YCJBX3BDk93U5giUi/CZ3easygKBSzanY
vdZ+jD89NxnJm8z3BeMXPeZBSrVHi4kTS9Nc4C/AuxSyykmIvdQd97V2uEhtMmp2
ECHYjJuMluX97RAc3gCnVwiGCJ5C6uQuwdgjn0iwYn8FsYPM6EUMMqf6A1LWhygs
AysVzJDkF1e7WdWyWxrzdo/eJtltkID5PP/Ups/pSAb4vz78OJ9nWZGPMj4BFnmx
ij4GhcA/rk16pzu9k9Re193QDOaWyQgHueYQJLEWQ6I+mXTNdomUb8JbEb1H7zOQ
fVsvXMKvu2TkT78DX7zqkzDT8498kQ6cnuJKoOPXDvOhdUD9cvhfX7aPWBHLqPfx
OKqYZD6i340zhW++PFwpT5YAh+jETXeU6qqHXgOEGJsINnkvtl8tOtRiaQsXoMwZ
RiuD4p2Y6OVSJzy8Bxjs3xwsg2Sy4AEC9tOvJqULjzRd+bJ7ClFGOvUHQ9cmo6ph
G5zwkfrjaLPkE1VmvcSVRKUDBUdCs21dCOiQO7qN9qH9hF9fg0FtTJoqdLm5SMKj
lDTlpDvAZsPx5p/YfhMgF2Tx1OdxNp5k6QT/L6Gf/H29aPcW7N4C+8iU4ewX7IGa
/EKWSaqrC8TzmdK1CEYi9VHIrc66/56KHgYm8Mq/dUToTcaIeiQPb124z19yqTFt
U0KhMmXTa4aZAVuRXvuy+IWvU/U7YFXxdq0jlprTTSYEVOZ6PEvFVbod77jwZds+
bBgNgwjXK/WKO7WYxsMtIP0MCDC/xsx4iYTAVxFxNwuZVi91wNzXlye5gSVAOpc8
pGXj4zW9PIyv33X+5+ust1uemSJhWv7HlZyXrs6n12vuv1rWd7XbQGaiMTzIOuwz
1AX8iX5MBHdELhIQvdtRmMRQSEDNXePPuaWuhc+Ed1kquwhuAd5gBNScjyDK35UP
SvcbI8vuJweZUp2U5nEfBPWmP/wYPkh+D537WAYwyTW69R90q3z1vL56tB1f8Lel
5P6xtlLdf8+o9hzmCHHO2QZdO2f69FIj7kd9ZROFgI+QjKK/xH08QiRPAQZlgye+
X7UptYE+vr1wPaGYNYK3A4RMlRyViAhWbK/Z/ar35KiHLiHCUKUiVt0Z8WdFqt8l
MHcL8vlDAH+ai4LZtaW+hok5paVkjwyfHN8VWUfzN/IU3+YzkbxtckpBUdEuXLCu
0D3K2lXOZW1es1WjNRYamHokT8b3XhjsLZFe1lHojQGWFk1ml5sw/aKDannZYaSH
9C2VEAg9LXuXcOSrInkruN9mAjjzii+k68F6rY6xSsVGlIisqeYx1ZbR5dLp3L7V
c9hhCASWuVZPe/oBHptMBoJ9TB/BKU0sWZ2T7Zf5yJn9UFWeT7c2v64Z0FoylYvP
EjhRBILBeQHlPiNJ6aKga2kgvUjCiivISnPmypPh0XDGVGixqzI2KcycbbAxjxXh
LNrCurkd4YM+cbPbOu5e6E9W6eXgGlG5cbSVJqQGM1BwKIdBs9HGu5+hHHkSsWmU
HEBJVpwo8fzKU3QXNWgoG/OADV5pLa4RJZMTfcB0G8NkerRghGBnxnR3OreuUigd
rPiYtFjjdl0e50RbHCWktuVyBHcL6Z81IY0FvA+UjO2HvWcFOVdbC5owwoG1MUg3
+FqM/OtgqygB3O1fe8anDwJXUC3WKwbKEKq81eihy1JUzYeiHti6UR1Mm4SuK/XL
7m/huzsyw56gkI1KFo5rKWdP8BimJ8TpEAI7P7LN26QHaSUjmtT/MrQul0liw+46
5aAFRwMl5bEJB3koh7g0qEtGmQYfrfxJsDOPo2wjx5F/+ajGc6cOiCMk4v0MV9yA
GMrpFR6ib/KjoxVfoh5anLtroFF/VlYP4iCLqVbsBtPzqn+Lq9dCjGiuDvYHsL2N
RRMn1vIm0kZWo6A4pcPZvTt8l+Hatv0f9D18+wxLMt1ibJjxr034b+wXli+DIweW
urzfQHaA8trOdhjbk+3S9JyXYhyztAPGnPKt/p2+DmlwV4N1jOigqjYScEWtp1xI
DRaXLhp2pDalKorzU50kULXGymgLE7ATZ/F9d4Ulhv5fll4kFAImY3Z2z4qmBtlM
XkagD5ptxsl/Fq/m8fVHO+78gt/2c3B3p6mnqOZjHarJ/otYospMEseRIlNbhhpK
OWnCl2mIEmeLC0OddjBozubJACn64Pfb1aS5MTtVNmqnQJ39PUz5sLhbUD/v7lIS
AfB3939gxY6aQGsqMtlLUz53ivIRzYuhpexanR0C7h6IQy3e5rZ7NyfafYNsA1Rq
XFUbw4eMGFSyxptX6611mtd99TCSLuXMu6E1YuBufm8xEQ2rP4zR84Y3+SlNv8dn
ImVqrFpitO/eNZosC8ODCKOwiIz+7dUlaZZ9nt8NJU6R24ttUVZ88WyxZHTsp3UJ
whnBTswK53vxlNRCE2BQY0gZhotK1amKKspu0lpWTXz2vPHdwudqmP4mHdjRiCCs
FIYacmGCWbRQVNCYTVNmwIa907Wu6ggjuQDAI+tccHKsnKuiJK89LWoPpSMudr4N
CV1uAsznCwIYQ6wuv13FMhMVVh7fJTedrH82OVJm+BCThabJUZuMEh8nZqCiUbJf
Nw5eg5Zwr/mFNgC8ZyeXn/H6SmnYva6CIE13tlP5dctEXpDnFBSplxOY1eGlncHg
Hy5F/XF8kio2XUPcHFlaaIBU1z12+eES55QfKbSuRAMLbANuufo7rS1WXUQDn/sh
TlYBmXI6pE8iMkdNnCF9qMwePGdwvX5Ibpu6PvmQL+jjQfHxpgoqC23OO3TsddnO
fyRmvcegsUV8P+FRIWSc/+RST8XzIwsEDKcS+FQtGNaSgr95ZKonLPHliTO2MG0A
DuryZWKfO+Ia3YhNRUURJd239eRCflxD5oKwJbCpqhtIo6MQt8xD+1bSboJCRZDF
gp54DT7wSX/qd+FIe4cgA2XboIreeZBOOgF3qDg7EnSrc1hJKcsCO08iYn7Xcsft
K5Y2TCElgEvNtQRhkrt5K6UrlP1u800yYyOCZwwyXmyTqK/nPzojzkrroveRHwRt
a/m3kJKarbVwS3fxr8uLHPHDO9FsOhFPdV/o2LX0cWZBJX2TiG1/sbP0mGOh4IrS
of368GEY9J0t2b1vOQ5xETuotsOtmBJl7dZoxlcc8NAz53TlB/3WgpOAF3Xyqs59
enVcsREFifgLS8kHplaRuzOo19uDOHV7KvvZe81CCsf7LBewGqX+4C2gyQQ7E38n
eT+UYwyXHgaDQTENG8SqRMxU2yRg4Og+A7bcn9ItnJRliAsAuZfabp2Awi4giL1A
yddxaYHNoWnXmYgRYqX0PXhLlnZyniz5x8ZTQzNDxdb0pdlyA7Lk7sJxSCigu87w
dtXkKX/vnHyfEIjSuXPH9RI7uO0bbghwIXXyJOPNSG1uLCqnSqrXseIBuyx+69da
HbWIEwUiZrQ592MBHnQ1Z8o9ECFmXkNm0f7ZYbXG+Oycc/8Rr7EVrXqceeWcrYJq
7BXMp4TnjBudzdsFmZsS9NVv0Ej7QnN+/bmCyvODgBkBXorK0+eT2SuUgcjgELbL
bvTTf5H0Y/1rgGJ/guEXnAF1HuFvfvRZnwSH8KZlX7M40vr22nZYoVFFdGb7nQNY
Fir1rqHdkkD8LC7vh7OzTCWMkGEotz6nVe55NYMOnh58XEfh4zWStu+sYxxfWDwy
vnwF913FJrbZHEet7XqP9vBzw49JxWgoO6X5AT+Flh0tUenBi/jnxsz0S5Af8S4m
p/s0BLbowKwirDKxJMPKadNdgirCAsQuctRfQeE4FpavIrJQoQVORFxvUFH7uqLs
syxMEwu0/UMUdkpLvKFx8sAJIi4xwhyDkYm+42Y0dMCKJzwIJQlmIfMIHESNWGi/
XgHN2yLpCrPdyRT7fJBXRVSxF1fH1RQ4NFyzrBxwQTwMmrpg8WM6du0yk+Og/sgS
L9W44Um2UKDxtWpqkhoAJHCx1SkRon6EuL8lLuHW02L6jgd8JFjyxvjdKviIKvWM
g6ecZwtZ04iH6XJwFMcOEizxGfd+MZhrZqDj2Kuw4hPkvNI/PTinvbR3Xmcdv6+R
smV34m6bO9Qecm1TkQU1b2B8Iwl5l4MxDgy1ovGrxVCpyCxrco0Q6fJ5yY3/eODM
bhZkfFqQy1Zn5diAQcxYife4eUgDEfz6z3qpA8l3XEHKgwH8QvCZflPRWdaoia3q
bMDM5q3Fv8PrJVBVGk6FBip7tV/iynHfTIAYurYqfrhCUFel1ghf4C9wm3YjmIyZ
M2+LB46o5V4rOzkAgjBdQQkV8gOHDObAmGEdfyZ+FajZeN7OhF8QbEwj3tQ24HZj
NGvvyL4ZyCSc9JzxZqhS6CyRR4FugY7+mk5BPtET7dDP5RXh1DdNXNphuXDKNVsc
2oWug/XmDzjtaqIUEasBWgAMOMyCTewB12auA4v0InbZFf8fNQFZB3bGJVycCqfX
BIhiKce9z0tgmU/ujejB9knDPRfbD+8jfnZnElQn0siEebt+eEvTPkvZayW1maAt
srOxJHSJZAzfZ2J9K0sTff+7r+FOMQ95CIeyVpQvT2mxedW8zv++9cVPb8qlaxdT
3j/mHAHLk0kHoluL9CZB79+h2gq04j68p3bzjEFHbjs1S3TsC6CXsShnsBG1cPC6
WHEuhSOGb9020TuVsPf35FfnAJtUxhyJeamUBAICNGxlAPqB+XfIBvrKKmQ8CeFp
vu8g3sVscbWdb36pMN5NaDpOCB+AV4/solL4RVmsDkjT7sDM+cCnTUVfTdG+qM70
ICcWfB5xG5OyWqHTkCfHl9k3XOy04hr4vui5Ub2IqI8AO7QJMyEN+hjs29Toy4x8
9JkP9gSPcLatHV5XhPoZdBuUtV8aPHEBXDqWibY/pAibCle2ZpP+wO37mNopzlON
bb7U4PKVMBpddxslPNb8Xu0FZBU3Fk7+sKVzcgkD/wcWOoVHthQgwTDAaKQY0l+T
s1g45LlRMkkRoBvdG6XEMfcAK6eN4/BG8lAYhEVer9Dwi2LwvqQ71E4xI+iWAaTs
zAhL8NdHhIrXc77TzIujz+D2e71/BkgrICLv5K23jdJ75GzRESDsskC/AQXg6E/A
KrRU7gwr2YSn78nz4ZbKYItii8OI/oOG2YI3gusS3gwuNw7sFVoH4JsJuetobIRP
tHZCpdn8iZVuGrK0AvU1IR+vHde+lIEW15rNiTPDG3RT/YWFWxswwzhDypzMvmCj
3zOGy5/QzPaWxy/HHCwbe+NSefoBC/GMItkDbl8gZTl2l5kF9kS5+1tJrwyg9hNU
ZQlHLuezxUfjjfAvEeWYeeB24hqRzNpQ3zCqOeFdIPTQO3S0/3lpigoZuWwrUkfv
9KQ7VxG0rLWNxl9EP3+pLEFv5vi96svMmX3sNs2qmo3uKBr59Hkd5EsPDydNVEXZ
/pDygXC2jhrrW657ghGi7xfkZKvpFxZef0MnJHkp8u3H7Gdf9RZ0bz4TVo0OFrDH
vwrjytXmEj3Gz6NR0SZYrTcSrcTwPL+oO4MAIbd1DFh5x+kOxG3ER7IMJaA2he7V
k8dRbvgBKC6HZjXNzqJbBdqQjRTqF55XOFslZOzYEFwAhTelk57V+Wh5btf5Ag8u
dbesNbIDlRV6drZZpEBiB7wyo4jYddg2cSAlDOyNtSLeFLji+bYIXX5XxblvFDmX
NSQ3C8zat53TTJA8hqPLvuzdxLybnJMVZ0W6/TUhjz7HWhvIuOyLV49ZSXrrjMCw
Y1lUwae0J8h/awxr2EDhWntVRNmdBIWlsWywuaHw1WEwZgqGnp/CXC9TdyjP/m0f
hFSTXyCL2xxANiqSc0BblDzJwyMKs9AsVa4padCLk8qxt20mogwNseGp0udK9+XA
4wTc5y1TywWS2qn/2CJqboUzeTdemR4VSGK3qd6vcX4TXAJzgbPoHHbd0XcmboYu
+GKtyivjMcuhNC6sihelDeaKrkg6bUF823eAUgt7o9YHvy7vhvSd6CUWTi1DNJ57
OOOTwtkiQjCY4IXQvDWs1B0mD2Xg6qTgbM07yDH0c1zRf22q+b6MFYPSO02st0rZ
K9du9LaJQAgAXp0Ar4UPYP4psgVGE22ANd20wE02JW1CI1xeCW/eftvXHH1VdHW9
bHDiDDMtFWegO33eOpHHmNKYq9JdLMR3JiLFzVI1cBcR8VQRLVwo8YkBICJAMY/B
Yfg0AOyjX2BzT3Ry6bU2JsH3L8vGPcl6mKRxsFzNqKNcAE0iTuecNPxJBHeTxL5c
glt53cumKjTT19VT9zIeTnWzJGFsw7tuiUdwCHQ/6buDG6Q2S5F8hlCGMFe6huzC
3ZJx0wpM8u2Nk1nuVbnO/FsLneZoYB/GaaDvHG6nESMVOrgOaIE01Vdv5mRwUr72
I+hCxRZDZu19cLncDdL7FlHA78YagN1InRd7kEhK93cAobyxsNaJpTkkJ+lkUfWq
86L3PW2OTCuvXxLFGfqf4z0sX+qHsdRP2CB8xvElcm6vesBNqo/8iYhbk1MvwaJi
MtjPegjbtqgRiUlYmFWeM8fep6zktkpLEVu/DeN8ww9MrU83C4D3ljixQtir3SCO
0lOjiMbeJPTKGSooBrzSl+VUA+IuvsmnII4wMua/VZfHHo0KOXKzcFx/T5jMgxwo
lMFT/4zW2XNnvlioZE097DyhcCZUKil6WWxUNpgN1g62tR0FhwSIJzwoQFX+amW0
w4gCT69tqgYV25jM4E6ashByemb6zS5p9PuMOIUpWYRkiepPPMjA8lNOVwftqWif
8s56irtrEFdjjPIuYnrslTgZZFtNxn8/39wCqsZ4f9dTw6nrPie3059qM8I8cBdM
B1qh7ohmYA3VoP2IsCyivNkCYhz27QqoXzcHSO1xUbQ9OI88J5FvR+T6/W9Q64Wl
gunzxqS+l7dXq435TI2ze0unOg+zcH2x7eXtnaFU+YJIBx3dHmq98qtZqKk9GGXS
XRtXzqV+dQeQC/gVwGBiGUr9Ut+8OqWsXBIVaCmykICLrJytTiKGFGA0lCWv9wwP
dD2tSUvAJJW0pZ4uW1JmfGPsh8DzeJpaGinAERZ8+1wbjhGN3X4UF+yETsf3IvSN
TsCGPwV55eSNtP437AGqA/FVXqRn5HwBQw57bfO+IMW67XH9k9KpGJC0DBA5zasK
c/71U0G4+k0hTpqKDQ2ZeO6Ubh+/z6rPklVepq3hydbMXkkMDD/KfMQ+cM1vITyx
Lq1h3MrQPJ2HCHtd2jZrLBZs8z/WvPzgMC5PfakOogLRxkTV+RoSjkbStzDUEmBn
NjgpBuR+zlF5tp52lITXkxifQKaIv7kz3gxQJsRbFZiEXSfc45ybQszISv21dFQ8
UVIcmAmijG2uy4SW5p06YynKLI3A6vWiT4vzEKpwL+qikFKshYOPMQ5CF4XurwSG
OBe6SCfODbRk6/VDDiSwCM4YQDYu+bcuSPRQQKOs/UzksHNdsCzVUu+0BLHhRt7H
wIKMqjivUsiy/U+Me6cvVzlQx7wxF8ohKYaPnpa4YPs6BavXtB8BNjjG3ogRDcI/
oA1T+DK4EoYD7L8yM1I5CyYl/oErWScOA7Rn1zHkRkLaSLHDLy3ZOVUnGxDDCrcs
6goOdpiwLH55hjeZPHhizfGEnVNQQ+yoH6+0hZrnnsE4up6HQBo2GB/OLawCPfp/
r7NxxuhUfVumkzLvhofQSZ9Sr6t7fcJtsWmjCl8J+JqJtEYC5xjrDxHPSLfx1DJI
9Sx7wBKrImupzD0GGwAqDXI1oq8TiDQ9MEPVmIVS2hIXkmUPT5rRudYVKtcUeu9N
WjYMgSt0w3ylxSKMrzqoXgf13rWUe/dzC0meXw6Q5eDM06v2mqJYRQlEMMySoMI0
sDoPVsLM1phmz3sVtuJxYWFaXtwDi2rUFiacvlNWFN04v+A1cig+29MD+u3B+X8i
hcRUBt47hM72LNcVmHEAD65Ay2UmnQppp6fsW3SjIENG7XSMuvIOgBMW8wCE3aug
ro16kY9kXKvYMfHT06SoWb1s8nlVvpbBnYbUMN93xHFSEBjPQi3IrqTKqOxqpaqB
ojnbjqXD6LwcW9nVwime9L0Sy5LmjUNQwZgIG1SerjJmZheygm4NLyrbxDSlR1cn
kx5//DDNzFIMwiUCbqsUL/VPqOZPakvxpOGi9ylRwLYgdUX208eXGJ7iK4RsQDC0
qY1Zrf26OCXabNT/VS43EGa2nuLjrDzezek8JfS+6NKQsczdgBhyNPCwM/5EQt1d
BPp7U6or5f8gsB6N7cqOIPN/+oZ1SJQrgqoYyjB+Mdio7zY4The399tIns59QW36
fLxMWIkL6Qq0qKc5Pm8+gSO3vX3Tnm8by4zQiv6xXratLg70a2J2LeEB1FZVmvFc
w/EBhLOd4DTgfqCbYZgrud8F4prw15iOvuPMO9QXyzbTBVVyleNGXIrY/qmF7GpE
noYpbMM/WcIorYrzBUL99+orL7hJt+vcWzE7xOSs+smbakAZYie+A4VGcJxe61Zi
jcr8jOnjaNy9zHHF+1Cij60JZXFDtGmsjOFw6IALMFE4pVq8NfAUgjycjcj3u1Zc
gfmwSbIh13txY5TTHOsGhdiKlAGRyDS4W8TGUtUI5kvoIL3lTExaAdIkLb+fnG53
/eNkPJwJNPoA4r3mPZ8UBci2cLLZ7kA4Mdsea47tSkXC/g6K4OvvHfV6p7MLUi3X
LS2JiOqfAr8wXBMWfmMjsdRBDVFF+Y3cFN8Ph+9HIpec14JQLjxlsx1EzYKy1/jZ
JxOqejM5fZHmuegKorU3k0BfoJTUnQJGAh8/x9+rcftt/9/LvETutnSAyr72fImO
gpd6to7id7pHLw2+1JNLAIXV7h93CERSBsPaOFG+7+dw/Wmn5croPnM6u68u2q9D
uYdWqk2ZXVAb4TjvDYWprg6xsW0WhZ+Nh+9gvtLYJF82YtBvuTiC2/d6PhX9B4c0
6YE0NHmLwqT3WvftaJqSSwrBXbLUMQSYnfa7hxP0x32N9RYwQgsaBqOczXxNYi2A
Jy9I5G1QZdR2TmemzGLHHu/0PAYrDgtqQEJOQyxhPizT9JHBnkBFpMtauchjaTNL
KOBZKnERumGbfe4444byRhLNyTKTQzhEbVSXWG/3Wi16XFFu586VYz+ONHLuvVAp
8p3P7+f5029YAPntQJzB8fM4rEoP3Qi7Ow0YudpFxICc9EpTU4gHf04AZPD63b/e
P9vNirjhJBblEgRJU8zM+uGiWqolEQPR5403L/5IE7nzAk1wrbri19vIjkq8b0q3
EOT7RfOgaEOiUkNaJeosI8lH5vjJSTdB/fwHsCbTsS9r/zOz+QyP6lIk+apLGVyt
d8e6z4QNcygRgKkV3645utZwJBUnjSr9w9wQpOXRatLIaAV0++2QHLdHX6hd4AwY
qhWKMwtdQZj/yt8QCWP2TsSJkea2saP6El7EUTemvlT4QhPU3sTB4O2h3kKmp7Gg
LbvgTRyjlWsnAR5C9AX4oEIQpjiCzMlLBYzjg9FLXOUzqzdVGHycugIy+g7LkE0o
Qhx0LksI7bK4sLs8nRcXDU7UQAMkomG05peOiBx4oRHOlRih5EW/RynKH8qWNkXL
NwFt2pBHLRRcUem1ty7y128mk2Gm5C2YdwUDbuhNjdP3EOsflfUjGdefF2tyNmYc
dr+ta54BGVip9yqW9UlO4a6cFUMatpNT9EvytJT549mqBh9c+rCMKe3i+RoNYxHh
M5ImXVnocDhl7zb83HeCsbwrG3KQxoJFvQvAi5g/SG1GLHPme0pDi4XOCFDAoEnh
zrJz3wmuJ9krp0yNwnrIgnHu6BEk9VTJwgfZoULAFksY6Cxn7+gonYxpEfKXL5G3
HCWIb9rYuGWluv09p4B7f9cc0nALGHqp0VqROwRqhlXIVtIoJv7nBjbEvhU484g7
+xpy56JnGqCS2Xpx9UhdRQYFUdI45VdcA4URc0EqwXQ2N787SRslSk34WPTnPNtL
Nz4y4HaXMNbO3Qrz2AH01Qs7PMTfW7OFGo8Cuxtz4K7HZfH1lcssP+jmrjJkxchi
Dtmo4YrKbnNVftGoOuY9WUA+WWeE7DLmotpSYeMS8zz5T2338RknqUOWpjdmxXGB
ktQWAstu18b/Th32ujfGv88ltVrq8EIoKvxNutg4fSkQSutSnAmPfgK3nBOQkW9+
LN5QTqY/tsakXMJ8TYbXZIuxpyGf04SyBtWEfhKPiOPfNWN8J5x5P7me67AI7sH5
Fr8P5MTngasARdK6R19HHVLN7VjHaIk/CWH3zHoMW/aTE4bkxo6IoNt5XoSq/y0e
xTG1XM61SNUqZSzXbaDGEtytBarEFs5HnnF5ikFlk5v6zsoigXbVARVjlJfL1LRP
bQyTjqFER471CFSTZn9KuzO9JhaKRbS0B7D8zfO7xggX1zTvbR/ByW9yygvM0Sh8
vqpTlyqKlAi5tcu5deusNYm8bTzf/LBKoyOx6fav7sYLlPITnNx2S85akx7P7JXN
eezPnq3qZw9i3+Z8npLonb4lLKgXCEnZu3F7xoWUvu0o5Qo6bsi/yTDqkLm+/zx7
/t1lfA15o8FGDzfq+Spj4GNnT1tGowQQzNyVRlHyPJsBwGTXeLM0xse8QFk1OgYh
f3keS6VfC2wQo2TmBNSu9ps0Dj5SiRkDqnO7BC7JgrznOcnfq0j7DWSY1W/XHwKD
7UKdsJ/w1r1SPhQfp7ZG8RThiJubqFsy4hQav5JW8Ps4bp8LjTsNzHWbQI9LIULl
npLGJ3+SAgFinGTmXznu5MbwcuN+2JKPo2cjEkGvdGVgfv1wQdEOqlj4HKHomOsZ
F73CweuTtLEcbZE5uwJ2uDwicgxgNIKTyjfBeAWDH0xIH8dWA03taCkQ0/Eh+get
tbXnbaDNQeuEVDHN9Oi2MOEImRqMN1Mi+qNBDFYthHP1NMQm5WAuX9y+/3oyhNag
NM9acRgtcwZ4Cr11jataMrF2mARzpZ0RQ1TndsZZkzQtGMzrm+VXF2ColiOcJPoj
5qua4oQ6B8o0Z9bQxOvX4iCLf7ExCrs4sIZKpBZh04wBaPTfwucR/S47IHdeYpe/
9GbSDjzpgJuu0DLs3GbL3d0aI6kxSOedR2UOKqtwLOesyGfygyw0GElgB4v2xlL0
we4YATPGbpMoI3EWNXkKjN94PzP6o51U3uWwJv8W1fgr4QWBRthbrjx7y0yivd4E
GZErSO9VbpTUZTTHJ04x6qD0rD1cz/3UUWQp/3w7XHqExOziuI0ApR3eTQ4LdHvz
GipboAE7R91tbSB2xjFX4To5LWXXF8BwcF93D2mTZBX+5i+VStPZH5rjtYHt0RoX
Ax3o86w2MpMcKzAVGxAlCEbFsfi2NAS541ZdOnYUIXxbywxVFNTXsrQrfObQj6FU
cw7DApEi6PciYh2jY7okfh1DLw48JV5ECOTMUZSsNMk9++pJB63OcF5wpmtfvtn7
P6bVNbFA7MgMql8spMBP+TCRmzYlJmL88gTO8Fb66qwNq7H2i8FM66EmzWZkfTkO
BrQprXqEGC/TA4B3fogZHmayMsRNp4Uca9NVvYULTWwGjBZ1uFQy/K0z6zxIHw3q
fEZcoVxl2F4jmkKnPqUdlBOQ379/1DGUmqeLUHbvaqAeE4KX8o0bpta9qDmMVCYV
xZ/s1faFxZS57ES4v+ldmbEIXD2iwHyorQM0Dk77dwXTRWfO59b7eT2FbEWOWeyX
ZP2p2LJzOdpaXR+JGSAlIX1bO/j+Ha08JMo9GZgC1ZQ99b4CVe1d3MPAGtAGCfo1
11LzoAXB4rjqeeW12aCM6AOs65I47L5gAUYMUAomaSJ11U+/M241HNyT2EvG/UAc
nVvZt/Mu9BYxrPlIttdQsiUdAGJwqTc5YdXZX2q3WGRMrMppsGhE2VGCX37dE8uI
CU664hrDbFNuIWlKrevYLK/7cTlvdXN0GxHtIla/l/v+tKmGieQ6WNvnTCza7Gh+
HKSsdVKd/zQEzUjaGEuPFcd1nRfzv5JJtlhkDVK7CErmhhGwadOGpZMcrgznV5la
pYXvIGRi1C5PdEbTSh0Qp4W9gExpDpcxYumY6Kzbavo76w41zwFOxhNTxkk/uHfF
xJhK+dt2rKwhAVT++GH5JZmZDpcljLnIpZCZ8z6ctgWkYRRDJ9QCn7YVcR9SOnCZ
xgK8cF+m8Wu2CujyBHUw7G8KZ0n0UVv7FLlaFg2YLZ8Vv0VTEzlg9IXzRHC7SnQ3
D1siCegz89vctl2GV0CfyBm+uh0lGwrbxe4VaijjsfwLVtDXwCYB5h6xZql+IALZ
9lGlLdvGH/XJhS04EPPG6ItL7UlquLTy4PgkEIaVgYciruf9WhUi0dN+gNUXIGZ3
Pf8x6n3IwCvqP7rA0BJvWwogvmjHiyJ4HYegHbQ2W1fmcrp0lBDNzXOGlHlH4YCe
JYCMASECbbnrhoI60gxzc+qPamlug0Ssp2nnCeOddT3KmyvfJuR2y2qXiMKmGiR4
S5EEd/Adv5uowU8ycsxkhaZp4J7mGvzd8Fsi89yXUdi6R8V52YQpVUmJjchyJvG1
Gdy9r8yZUjX09KYEK7t0WNIiJKysyirxMbgrfHDK37MtNi6HRu9f+ISEdMKxaCrm
avHPwbhFihsRgp6jMhLtzLUZ8ucILN7Rkq7b1yYEwG+StBAYoNHU2M9yLC4w92hk
3arMISbGvgIez70nvc34vNwdt9x3KDF2Z6+lmhdbx2L34lJUOw3KRm49dUK5u6GV
3/9IZICgPLKaVtF9cdo6luae3M//YoMefvctW1xW4ujLxW5BwYVmBQRJuzxFAGfu
fd+NrT4CAotl0FSTAAWrfKl9mkc5qZxfrgJ60DFS34HKbfuJ3stkiYowOmfqWdhR
HB3KGDYp332ke57Cn4Wq75WrNlsKYvrn9zmKopoPnFZmHHCOfu68BWttTrW9LvRY
u5ru3xzZDxb74mfFaultfVF8c0SoygtZ0e/pKJ4kwMeNmwnosHfBTyMNKbAeTCaH
H191RfZBFMB8RmuiytyGXfb+Qi4YL8bherCFWi1A3H+mZOfcxX0j2F44WBzh6bwB
3tF0HkTwc1e9xxHIRAIn1NQJA+ao1qF1qUK16zQe+7VSmY9iV4SA6LFPPznetj5x
akzpb8k+DPjzZzGcV1ZB8Pc+qFPYmJOtUrK6yRGmP0GY/DNZiMYY0dHdTVD5wLpO
P/urjonog5a49bLHfvaBQLpnUAqgq87gnbBrED6JHcFYPd6EeFSW9TYFBCwjpEED
OXhHxqA4/ibfNMn9JMb8uRlUhVOEZPxbT8GQ4QltKs06oQMPP3h1Hgt5EMv8TCdw
q76x5sZhw6P+nST629YpUtc5GxESFrYeFRSeb7WnNmBWDVA5hMw1dU08VsUaQXWq
4CttKHbbXa2bYdpb/aMZsGBGeFz2eaTACT2KQfxgLuNFQi9HtfFS+2fUm/AwhvS4
fNrhojWgCs1fOpArNXs4FvpROMlkH2QC4Tb0MicAF66M9uXQJ+3tg+/OOqf8IZVV
OvQVsKYPKJEHp7tTxcaBDCoyvYFqg37I3WZAfyFlKhM+n+CKL6VSl3tvmycdKv9l
7bPFQXp+wpvXWs36lNKHQmKmp7Qg9+lDL9fwddUSZdBh7lbqSNdfAssI9o7akCNS
2EYnxkGFR+UpQeob2hBIn7JcqIMrr34MuEfWZxGxp1Y1jorCrYy8WYZEEDP+JDHl
zfH9YZr/RpvajF1gGo4bP3jRV+aqQuBrOMDwgtvETe1CS+NwGjUcKo4Tep5fkGTA
GCBWKMfzUoFDklgAs9LVgWJ6rcAIQLVJrALd8e0tEuKcJzlb01779h+LqrwsFrxF
HtNkxYYpJoHtl4z8kAfcHSNSfbe0vdKfrCzra2lI3X+RZk9l+1z6G3MlsnXAHyVA
LquwTBm8ziftEK7m6AjFdb65M1uItrIecIkYvYOBYvlq9SjDPosFy+p0faMHuP9U
6T35yfVehXNd9UGifOolSJ/myNZD9IWLRLIywgf8tEIGgyQrxiuxR/DbSZTqt+fP
rwu9x6fCSpuJlwCFWCpGlZrwemy3Puk/hW7ZbAy6vIhy8JXudOish5RPEev2hExc
ceC4n8ElG8NUjAbS/8RKK5h66U7hPgj7mJWzxRZf9YLNrWhvtHgBO5duFaGH/AH4
PzLoszu+eAW7OXc4FdGCJBBXPXiKqsiQ0aEXXDQ+z6A4vCC5paRCcf+FgrKCF8bQ
Zkt8Z4WpJpjOFHtqfJdAlK+30BKZdz63RX4rkUzEm67PgTjNQQpjNRVs3rruhLY4
7TJYPOTn7/beVAxacjof3LZjF23pEuPAnKWAHcFn1izNBUJysAB++rrXOV0KVJ4p
kRZ9XOcJvJXIcfKTeXmF+rJdQrAFi4wf/gXgIpX8abOGc282eDZgs4smjWPYq+RW
LaTQ+ajzSloEK48nKqXGLGGCNmRt+x+VtzdzSmQu0pn2UeWnG/A1ea/xqPKQTVuB
H7AH6bxkVDzNf05VaSMcgetfMOtbFT6gNNkZrKMooasLR/O247hJ88B6031CrQI6
xJ2RqWX3eM+cGF6fjn6CNQ8wcseRHN8E5X9+PrdvCh3lMFzAzvp4WWev+Z9B3kwl
L3e+VG+0G0M/rRGiP1pA2JLtygb5sBpj8LLbgokAFsMNFudRp+K04LblEkosAjL5
Nn4GgjnT7ZeYIETxM1x8enz9co/zmUU9CCTw6ljgqbyTUwe6BBilyoLJ4Z2nUGc0
yNUyrQnLN87RsMLJqZ+1Wf7vr7RZgCoAqN491bk6Nq2Jt5EzGtphF8zpOd9z3FoB
FC25Sn6qD3WY7yLjhgXCx8C71rDm2UXYQk2kuF3JO5dDsI7YqmAnfSA4FGlVg4yn
hi8DUwMlMY271Hiwp945OMcgHj5/2j6VzzdyEZalyuIEVceDs9VaGldDukxcXPRl
L6lE46u2/kIbp6vK2kyiOzJoGrAdnN5EVKvRgtiFceysB9Ax+Z9d2T0ibNbf5pBw
/uZidMDesxMV2L3lbe/Hb5qCjfZVo0q6PiGZw8rmWGqPeD0Du5GAvDFLgjUJeYOh
dQzU0U2bmAfWNjRNXr/cv5m4ZJGn1vHY3Tse2C+DZPLwyIjCswAxFQEJDmvou8cA
0aiK4vwUU9BTXhCBq9q/fa3Dh3kVGtlUx/WNGFtG8I5FRE7egsZG/cWrHVXtXq/F
lb904CULizzd3vTKjOcO2EamlOxa80iCLz5kHjDMIiD/1hv0nDjUjDP3ILXio+K6
2iebdpV8QSYGY00eRQdhx7lVxwdz6/9ktX9TDGVEAvEie2rxPS9OnEfxaqbnuFWn
zQlzWlc/0+aCKla/w/k5NkzR5OtA8AOpq8i58kuoaB2BQz8TPp1jECLjogWB00rZ
TcWeWSoigdZm8pITNVeKBgGyNeCNe4AMnDZgJLI1560mNqBAwPGaFOGSa2zZGn7V
xk5jxlE53Cie9RvUOaPAn8lTLe1+SdjrHRMo2TTP1tOk1yqNai+f/iLs6mbI2eGP
ObzFi35Zf8mvGMOoHe2wYNUkcENmesSYxBkd9irvL3dV6FqP6fn5aRiKUnc0aBX/
D3M1LRVQ8IWYTee5ZnkYCSG3y7OJsPO1RTp6quZ73ay0JS0yx2DsnCW/Aq4uLSdQ
m3b1+sQjXdxCVve5/5KfP//OiJVqgStwUEQu1BjCrFxLtP/L3NMn1s4Q36uVmqJw
k4TeqwiSG0Fr1CYsolZN9v+YYtwsLSYVt4WucjOaTQ1yhRFpmvmfzTWhDJambDD3
SM5cu9ZR0qpGBoaRgoKA2vdLMKSfRPkldcraO7cTe5LAeBKp9eWxdSdZpzVCVNbs
XDEFlzi3ytjByEgvsqMNobN8IqEeDWMy9gKqCoRAHnmgFAD1HZa0HslCKu96amFy
ESRcvFzzVzJfgR1yoWvGBKfLrynV7jdKmARRnHbpqatzVIFObAsBJyWutQlkRWCO
A82yzsHwio17Vy8ZAEkf8kAKRjHPVpwz5xSOV96Jjp0E5HKHoBsnV/dWmEc/bQI8
PxFW5wXo7Zq48gFAMxHuIDTqfLK+FLzXZVgBzbl3AAXniGaUKPravWUUWR+4GA7i
r1OZ5gkiO/k99U6oUg8faX7fmhZZ3WoOHMwps7AOBYoX6/qbx0hjSIKA7ANLGif8
QRKsLcAkg8WZNHYxaArdNpWCXErJ/sWgtWtnGqt8WHr/zuYHctW0Aeos/Mqwgfg0
9ecyovFWjnwnQvNYU/IYjh5wpJXk+9XeJ81UJa3+r1HXVAlBPCQcedaI9V0vYG4g
HeGJV7f/64oO7rf35V5ZYAG1wt5ZFaYCzz42/b6RyMoutlmbOVt4gXyTKK5QnCCN
drcP2OThV5nY4aQJ9+vo2GlIKYPbevjAEcq5fqVDYYK1oCs2Qt3VnmTyRbq1hxGI
7jWUIUDf8KFanuAEN878BIkz66ScOFXTDJR2IlYys0ixXq/WAKB2AWNZweKZG15d
Vv6hz7TDbS7VcCSS2H4KUgQBENrqWNA9RniK9BF7rITVpSX8Zp6rDa3bDurrBovv
3M2aav+8k8vbYmzKEvVdVsU5n8L3zrjKYFKZAoHczV9IHnOZHLEy1OfzXYNZRZ3T
e72iOZisIVmN06pP5KXIzJkdWN6qRh7Qb8Iq30djLhYjamtfC02MJNDHsvNxE8Wn
/0Kdy7r4W3n63LhiIjiMopFvgRwTqJvDPMgZXgDoI+4DfQXS6C6L+62HylIpFMV6
Y2nyvYUi74Z0YoRyqzax4qRxzAJealawlbrcj2cO3gRaUeCV3oU2qCRXmXz2gQzi
kED0mBUeUV9gI9ThqOsZXFuOLvqNDu2eQUDx4juKRL2bH02mgxhcNYM7lSEgEUC2
ytRNFKMUi1NGc6WgBtxI8xNcRox5UJOD+IcMaz8f6zCBMmHmQNGQZB8macLNp9LH
tujwnBN7HvGgYoBwyomzrxI9Rt9fkkjtCQZzQrU2+3DtEtkQKlAcJYtY1hq5nwun
sp6Ua+PeR891wC2PXKIjCoYAgIzHh+s7nc7DQFHDgfd1UF7GCDhGipqqQDjSJnSG
cKczlguaSNRVyC5ZwRgTo4UsdCvR9ubJ/VN0c2E9aJR5KL2xBWbYfDAIE3NUa+vd
PpSPbcFuavF9ILt/zE/eHe+Pb4CFWa1YvMR7FU6KVjHR/jXsWsAS05QX5EnnR+cG
UAke8ukaC46Mu7fZELVk9Pd48V83aPPAxOLhFP2O3EIe6PafrfQ+JCcnNSDTRE5Y
1jcXZKQZ/0MS5BUJc3NBGfxtXz6oz4LS5Rv91i9P5VyPtGMlrbgN3sjlCKDfjEXT
8P5p0pZLVyJwKut5akirvVeJKWremv5bkSRbmhnSlWdkmrWMWcGzjCJXSp8fiGg2
UmMS/yBGoXoY0R5WciFJTVZnDkmHComCPJ46ovvsXiTAUwB5eOg0hdZXNthqwHEU
6yap7e9gosrQaYPruo98Xz91R9A32YDFq2HMlP79mVExrTTLVAW4u9BcizGffMx1
giXYELS4YaDdjy5H5P12OcJDg9EYHTcnjBInbubiJT1u1dPM7qJj7I5Mwi7+vbIZ
bZGTfEoXyjsrz6+QG3kTuMOyjrLM283/bPUgd+YypsbGv76ohWiNBY8FcaPZeoL1
uzevFYmXMsiC+cTlq84TaTusNEnmjmWvZubvzGvgH5qEQdZEooqBqkVyzSmcTjnk
REMjElGGBUgnJgX9EovuWZsGJrHUoUoCKffZ4eqrb+WHL0ZxVcSrDF1NgE9jMbwV
8BdZ2M2YGHHe6xdfvDGruqKidodWCZlCOo0DCqDttcBMlncHpvlmfqtjUlzfjGmV
MFbvEsn1gMVoWj915XmQ0oCr5sG7H/SGxYEn3bHZiXEXmAsMew/0/q9kIBrD8SYm
cSs3RYf9kgXGzt9ZyvLQ+RcUdeAVcedI5FY96CdEBkjzVFD6/jfm2QGBxGk55USq
PKnneskSAP0ku5/dnZAGNj+ZkBXWNjkm6DWPmoE5B1eXJ7yAplzIt1e7Utdnw+Aa
yi8EzCZKgFA8Tk8HLnYOxIpDxmK12PpGlTbbCpB1plGaKGXGXInhuykKwd1sRkGo
ht6mvrlGmFSgABA6zdwWXVdl+DiNYlgASi8ZRzzZxB45Zp47E+Hj+Vy/puzOAk9A
q7uWXkh8lFfunwozkNReeDi8XKsfKB1XOtst+QSDHzNwZronFGJJSiNKb3hizAX0
qQPrQ7CtKHBaL5gt9adAUsPLcu7Amkd4WeHecx6fXxJOCQQTm36coibbfSHpkUnf
O/hNyJ9DLK7H8gw1ygp25BhR/2Uc14jYk+YIWrcq/ilQu5U7yLnPZkdFpDJSARkg
vHvqpV4XeHcu2Og6r9Y2w2uUJqxW8CTD8qLEivgheQqCNj+xq5MmODbDRp+2UcEL
QVrxNzLmyswKLDbHG9oTGkykhFckJUJU4KBpDazZ1U+t6zMC3MvBaeeB7WDG+k71
npNGPcbfcrX0stSmFaTnNausIMiLqFSCPv5IQvA8LYTrstqxeUpLAqqGv5qHHWB9
eGhFllQinEGhO6d5uriR4Hru/mYvlwzbEOn86OFiCwqzXxzshRLF+cIAQRK8uPNG
8e6SU1Xv+IwhJ4fGXAsB/m1QpNUS2wcVbk/NDtnm5WXOzJK5bdU9vNuIdl53svXw
Lfj8f7gFzWPS1/FRR4+omXJOSZDBxkR1R+SKBdZ3hkDQ8gOMfaBZ6NO/DVzDW1EP
x0zan+AKBw/axYIFooTrqz1FnhuukNw8rY/bmjruxrqQa0WwBjvQWkloYdP+gqyS
zaZtSR7Tg2/w2VLCGZWs43R20FiUKyN4PaD24j0Fy1hqCwMVX7EmUP8B6y2yz72u
UCMdYTPk9CwZFQDcpCVcJSwQAREqu7cL2qEOGCScr7c1sLun7938Jv504CxAmPwX
diZ5/DcSOvhKbNHqfKvkztd6ofWde5Guiulx8bCXNMpsQG42IwpUSaJCA/6d3wh9
on1Q2tazHT4sI8ELoZJvRdkyvLobBEBsbR0J71Lkm/xxGC4IjWec9Dw3UsXGZ2WU
SwfoJ7IrEj0wOSOyvsPd0+bjzqG834ULeOc0xpPh7nClJ6bq5iQ3k+q/mUWN4Kdl
ieCErup/la1Msw5ENcUqToLu5ZXU2daHjNwsDbg+8HSONke5GVXHhFDf3zUzrOE7
hV3gWrnL7DHFwxnIpuhj2TJ9vxbcZCycV90uzQ4C2tfhqU+ngOFV/k9QTa8evzYR
u4nXQO9eKy1smjBPNrtelu4Z40mlnsESP58katIO278Xb7p+TFDfHZgC4SCL7eGI
AAsoIBp42uojaqhzGjIgQmxqaXRB1Ob6QO++Uh7oQjrh6sfrguyoZS8oEH3T831f
DC3b+vdL5xvm0YbXKBbep8PUcgJgfQI8S3MeixQGtnx47/X+ovH1kaWr2o1Q35sL
ItW2NgqT1l0qidCXuwTjCEtH+oN9bJvFEnZ1mGX0phh2Yt09UvjQIOPXIIIg2Y1g
oOfo1nFQrLnmhX+/ANgPHT4mgv/Yse8hOJ/j69aDDhAoCK2B15jN7xnuvojokpW3
76pnMFEdAzjHETN/BHrACTPEe7ktVMYqHGxGeYR5R1BpqoTGivzAFfENVWTAD/4Q
ogfJ3MPR4lis1xsMIUh026tsdoOpVonjEcJHP0GkTNgxdMFIlnxKTofXCyhI2mLT
zLhs6Ad8j5xzljoDqXv2cANQfDsj7RjTnePNqScqyHFnT3NhswU9YTCyRXuW2ssc
K61lv8En4blQ4ZLLTTcz5Ix7YDFtkNQSxAMeNjcTNRGPOCzkdKly8qFskaSPKTYx
QlrNjuN3sqST7B5q2o2DqFNlm6vua5BHPtSW5wFBliZjmCFDdphIwiYXR0fgth5E
1f+F6Q0eGuHAQhaCcWsxWoNQxL3qhMfJtdBwhbiKt7BRWUxRQMEcv4fHWT6XrS6/
u2aGuLezYsTAmK3bdUmjZvd+0wlYGIjyC9/tcvLTdqL2667ryyL87hWnAKkjYs/3
jwE4OKtv3mNIAhtotAqO1noc6LlaCc9K2cz6NrhHXmejK0Mh3v0hEGNZGDbKvB0O
Pj/0EJ8oUVOkXmON4tnlttpI4pz+lqJB8h/NWlhzU76IaHYByi5YzN/2pgw3nuB+
t1m7TPjoygbSyHOwSWnyE/4JmAB+a9imxPt2hlJrsyE0yMx5aJUpYmobxkxH3QKm
3xjh13Tg3thuH8ymzUQdhlqhQr1PB0vfnzIRvXheDkO3YKOJdbBjQS5Zn+ExKVU4
SoIdK6eBf4CBuVO+E8isiff/qE/vQ8D+8PSVt+Ll+1Kvs2aY9j0HFcGFA3eVhvez
GondZ14YKS+E4JVMLsapZDYOi89pQfVu5YWg2JczTZov2LsZAV+TEzp8lvbxKQRg
ZjBQSJ884fRi7Mo1ejXPHSfjPHZOFIyfB7Sa34y+49STS1fLIf9t0IbnkTykKf0v
Im+1+otcNEIMXzjXCOKrNnXU4ahVhsh+7J9mPI8jWrEnAHcaEkmDe3PC7zIWZMMS
99iNQldWFgLThMJSHA5HqR2tFCuximg0MwOX7tfnehHZgyNFEF4stcAkqMhtUeZs
JmWtHRb0gxlULNRo1LlZbP/L6a/Lbtiat6eeUebiHFVqBI7/Eb1CsMK+c0hLtfOY
5sSYLgEW979tU8KeK4tC02jBfelYO7ms39qk+M2n3uXh5Rw4QO6hLWcbSjtjTdmb
YXhnb1+gLx57rWCe83HhOJrlf8WBTpC/d9bjnpduB4ydwJObv7vJEGu14N8m3Rj0
5+7jCdewpXASqB84W5SOjbqqQYANtUYXp6/zAcxZ/A5m1qI27jTeh151r3bsEgQI
bUDew4IfQ9o8A7v6oH4GblkgvEEpQJee1Z6D0WrFKkz7SDUcihVHgJQXuRwDuu45
fmqnWcnONqw65Vczu5YuqBhAX5gJUsCZRqkSPhfxrQV8iY78cJjHH82Alb35PVLo
XDJ264xQY5sIZe/U8QmRO/A535Is+LqA58s1HJWyq5IIp+w8w2ngku6dx/0vkUDU
xyqc9m8uDvQW/uOBIF1VmkztBmzk83fNUijlbdz19FB0kzo3e29VeVgbO7djzQn/
/7WhJipFhqp/cIkpAxpr5JLGTThXxPaHSB9qL2zTsclNVHs3Yf9BCrPjDSH6xlMO
KdbGxD1PAApcQjh1cufSbk1CFacjZOM5seL4OfiDhA3EcYfu95Ne8HCLFQ977sFL
+9vFa+B1J5c/320MiTL6j09S3YhQFhNO/R+enYxjZpqWsQAOUkMDLVfmLvEUOqvl
ptn16udAcC3qb2NQ1er+S2zIrRglBSGJ6BHPa/2+T+vNHGr2hMRl3lLRMn4Adr0E
9lhWmOuu33CmpVMCPtg761RuELbv+YvaRhgrlCrE72h91GUKFFrK7ACXZbCqW5S1
WuaJXJL5RpH3wYzIkalBeQRtRN/y/WETgwo2oC6lUOBdGMTFVpcbbwid5f0aWNXf
/VdARGQ2Xy9rzHHwWt8nFT6pPSXeHZUTTDE86zW7Q8fadMPbaPGlz9J2WJioqf7I
dCmxg8+IXkaa9zV5svd2PXBevbCVksIYOCqHbgIQpWon3F08wddvj3GQ+7syYppl
nlb066hEpf0KHkh6khBRU0smVybyqQjUarfqT3F5oaVtNwl4mQHNHblACpHIEko4
Nl4ptNFEoxktYPAc9ndIqzmwboop/eFeFwWHpZA7RGRJvAo47QTGKJrig4lLA8w+
IN9/89qjtBrBi8Ea7AtzxNw0IFogEfbpq2IMnBccvCk40iC1/YuUWaOQZYQ8L04b
RtXOYSmITVt+2uQMpx0AfGXQHPof4TDJiY5SAH6FPWGd93AnljdLuiCFj2/gia9t
dN+Ynv7fw2gbIPR3MU6In5sWDXT3OqYKnZ8tLqQwr5V1PYe7Ab5jXQV3gjBb4v3j
ZrWZWVoZQEtqXAyZVAhAlODfo2Ea2EQNcu+W32GnejInJ/eEzMh7d3gKabm4sJXe
aJ/cI5TLYz78oQSdmCHHuY93H6A0Gyg/efjs2B45NvsEAVkW/3md9j0kPT5Nw2SG
GuvjJJzTcX77kp5q3nIJdsKWg1KwR6nOrgB7frQoVfzslYiXO0efrL3YRHWfvfNz
FPiv1obT6Pm3WsVKKv8DifcMIoQRBs4OC6juATleeBhc9rpMNqHIHZTXLap+nauV
wIqVnFWZt9klgMoCt6VjKD8ka4X9XmEOsLTTDGjbEYIWeclfqZYSHQtvK0H0qfq1
yWYymvi0NTov1MrgOkEIBo7HuqlAqlL96SF4l3MmzVyNA8gavbsYZH1ZAhI0B5g4
StqexiE5Wis5bDz6JZVo/B2qsTsHEwUmbY8i9xg8jr/xhAn4n7bYZAbzd4t1UIhg
CIkkCPF922/Pty1ri54o+GNUzxVMngPRWsATgCvsRj/0THsfbB+JxxMlJU/deoBZ
6Q64GGEMsh3gKihtPOuavBsChpGZuHgVj1baadpovwdwRmF+b6RwsOiLaU+jGHQE
GKLENs/mvaFmWVnmfTUtwOE4UpxkBXKLn/duikbPr59L5hTGcrZfDbEtqBJ+Y7Bj
CQoitM+QoqALjsaIuwCZfrMOqyxymYPhXI3NA+uBOply2IwNNYiPyTd1My7yJeSf
JzFaPM5WpHevcUweL55Qg+thYSbmMY2mKauTmSBV8VmDx9Au6wDTmdWXfAwZ1FGf
F+m6ekjFbrSRZr8npuGSn0v3B9S6TK56Fc0iJTaEMoeM7fvdTq0dHi/GZ66pPh3+
TjhW0e+y44XEYGywtjOm5kjZW3rHm90eeWD2LwICx57V1u97m43Vwi6LPqbjn38n
ScZYaphagjNuydINR/EWNFrA9jXrV5TBshJBAi8ybrPzKodB90+mQnFk5H+6Kdw1
zyPi0YzeB2fJlTKIFuJ3cBHHrhW5yZ0ibe3Hz3LtPlp0UIso7bEVH25itJLAljAc
DOh100WthLVAlIkzorkB1xErbSB/peNkK0nX886KXgD7bPEhhikE/qpOJFljVrKL
hqQ6hsNzJtDo1IC3bajagoW0rwvot8X5aaWyWtLegIernObDkUukOXpgUwwfcZv1
lDemYB2ac/FCvskBXLG/4M0Pgwxi+b90YO4Tl7F07onRQKkAhtMPlvrDoOUD86Wo
YLD1RNNcnmE59t4Bk1WQHStaK40YBky/N2Te9E9sdx91fi6evIIeb6RLXtR7mRaD
Lm7LRyPAIzwJr0rpHQcO8V4NPnibgDOworSxxskf6PjbBASzGUICAUUKFjVMyh6y
U1Hy8F6EOmEaGJAALrqau0TnbVZXPhWsF5DxmqfvOwH3/HIefCpMW0YcGtCcxIxH
1oM/c7ZPfgdfuDUAv8Z4szdO359b3x2tR2+QohthauvQcf0u3sY1oO6NM3V4mp+M
n5i7bl8Xr7mgioG5LEGLuhtZexTs1AbjtZr+bb3bsixKY9f4BdG2PG9kesvJ2vuX
izMir53DBF0ndTdelNLkaj2XtVk/Q+Igf8cZpHwYzgT3Vvg1Gu6LELCHA0tPNY9K
GU2VZJcbZoq/ae2hfcPDc+pK1+KqADNK7SU/EKKz34d1gYsKTLB0ADSFd7XIXz67
H4ip0OjXaZ75PQLRj81437uRW2s6n/FPyoktO8iwmd+Jyzb+3hw2jF7vF06+IgTP
Rojo+z2o2dUsU20awCGAvBZcH6kqL3veOl1d1SPnqWlix9JFIHvcklhIVd+XjLO0
y0p2HkX1tfeP52tpOKqlyHiaeB9u8W9zA9uMHIPm7S9uWR1r2zl1b3uJwwQDYKY5
ZgmbRBgXgi0/RS5fTFxwrKqfmdN0Wny4ngxtNJ2RICCTMqpgcpl8y58WCOL1+Zdz
tJBH0sdomor9xlf9XPdg+ncOMi6legBeLuPl0MCk4w5pBu7cjQFGNqXmLZz1j1zC
mb9Txi2bDn15cvrwZ9MTR5DxVtCwPO9RtZkTm9YPUo6GVmLQ14IT37GqguVOCQro
gTEVDv2149IVHh1CCZLJZEHvloossUrkqPgSVa9fNltV1rtThnfcy8QhEoP/0EHh
RkTQZI/V+imyo0DIC+AR9Ud7daQq7ivDKIyCibdZAQK7IDSvRxcwg1gXBQCnYkmC
6eIF+eSdAy80oadtqli+/dGX7IHLf7NkXS/MX2ttgMJKpeQLHfcBn7MxwsyTLQpT
IWIDpz6+aNQClGevLbpnD8J7jw1IpQeHYd6o29wqwYyCBTIoorUWL/gjQQ6iUjVq
PEolt4YcH51T08yvDZ+JsmdPa6Jk6PSrQZ8rc/G2/27mYn+wbAiP2we8Ug5/KK6L
/kjp9PuYobnPcEgrsLrP9G3a+zDJuioWcxRb15U0mSouugzcju127Ky8Doo+qIBI
9M/mK/qBPZc3TA2Z54R8hEA6CevjnlLlZ0BQqfCwyh/3BUCNrwTxN04Zwfdp4Bvs
ebFkVzOk+5ITsRuFVQeC3hsV/6FILFb/7y6NtRS0AdoYv3kQBfM2p+kYKybrbws4
UA19rZwplPrORrPQqRwBaSjwaTSJOMuehdqfedrkjkLOMeCxHFbGeXU0cMKzI+c0
f+aXwHWHqTjKsWAIR9JZ2pO1Gv8RRhX/cDqDj5JmbAgdKxsujpXrJWp3vSV136JL
aTlB04uzsg8pbTuAbcfvxARuzdER06Toxb7l/nGxymkHke3M+u2caT02j65XbE17
6k19GVhzInv6Za5MikeiZlCsWbn9PfOwRiqfndH3dhDU2ltjdAONZ66vL6eQdaS+
qQ3K1DoUVG2UpZP4PLKNQwco6KrOvIMlUTkm0x1D2a7j31apHPEIUPkkbrbnaOF+
bskJmVL9741hYXwIYbar/CbuFLMLC/Bef6ysBLSCRl20UG1ZrcliLSOzMDJwVy3p
3cfnFHRYt2U4s+NTtwiofRX09nfLHfw4Vuo3OF9VsMU+V1H/TB6IeUANQVm6GkWV
IlmQl2CwX7N6EsuhtQvfeb2Iirt0HnH4j51BcJ2tA33HR4fEZRPBlXO49zNXR5cY
PAPOuoMiE2y3AqQgsSIBImDoSGlGWOpAuormGGySh2/51O2EsX254E6DDlXjWmXE
d2w5ZZS83TpNpt/x7/08ijG079m6JOy405n3QBxgs55ELvrHY+irZcWkgrlo/sLt
deS+s9/iELNxPMTRs1zKjupb81c2jrE72w5kMTXjtYlK6i4pjHZFuNiqojpZNtxW
2xVLvz/P4PsZeqMdW+47kqIPQoWMSBsyK2blTyf/GMCLle2cIFtNOs0H4hSOdmBr
uQBmThTCPblLQ/cSOSgd3++dwsgK12PTdlZlVFPEm0Q1tbAqnSwi8MswAZH1NBO5
HsnlNW/82D4HdveBI6LsWB2iuTKj2yS6Y7zl4+pc1Ei2GbPal5IxVdnt8KylCUZ+
qC38eGaxGx5TO7Riy+m2K8Jlr0CS7Uvl1r+YDVjYoFV2ABXm9djKdUO7/sHmvIxY
Qa3H5ymnFHWq+70H/f8+sk2alAy5Kd3fVfiaB4ONEfPN5b6TB90nACltpxGspA8W
G9FYow14YCkQZR1azFRmrfmR2g8+B1mGS3tpxppFE0VU0r0QXqTYsOtnWH+Ubi3H
YZw3hOYV5V4yYNoV8xU0rkKVet1guM8tr+aHdi52xMbhGXr9aye/iatIyHs8Q0rz
TKKyHIi9ifTqD+UspHY2NkMKCU2onpPiMLImic59Bd0yOrw+sqhsDjRbPTkegiMl
am76gucU4kYgMv7bF9Xo/fBs4WvKIPKP2fiClLCTksQpRfhLzDv8bhCGtMkLNc0P
SCldTVjTplRMCX6YumnkyMTmeUCxDavU67UPpFjkzY8NC5RWGfdKl0XsK7fygcoF
KJrSzEphLelBDUeuuQ2F9ZTmOnHdi6ZVnESe5qhW7WOIjN+Oc7l9ku55y2qJDL+2
1YlccmEVXQeKM1JnHnfwmHddhS6ZUI/FxJ26iGpBa6R0Fq4VLTBwsZdjDzYQkku3
e26hIW8DTWLfwzaGUd82qV/y9NSsQu3gxqDOyUd1OZWey8FsZEWgWPm7UOm2ZumN
38chikHmP1hxDugkqMUVMtTFLPi9kN6HyUblp/9tVmqNkPFEoAabs+7WWMtbj5Hu
pjOt6pIaE1bfMN+2fOj+sNgZWpLnbIizgorOtYm4abdwvyF2qUIkoLAxtSJfIRVG
sIitM2/5n1OLZYQDenaSw6jQa1jVEj4PoJeZq+LgqYK5D5dmiDw2cGS1ZuaO6dkW
GeLNo+GyRYf1PkFkv9JJySFBqq+8awgk2gmTrqJl2bRAR0QoUttVmsgK8LbRGofg
DHVwXfakxP/YPvRwDtXMb+7TjOve/HvQbXvOAvUyAm5eAnqzIiG95JReJjjY28uw
EPtBRSxRn2Sx000MhgFuOCWs0FtdV/tTNJbJ+eQGax4HmPWvQIYJI1OG0Hypa4Y1
6J7PWw+in965+sqAHWZ/KBYIQKz+1BJ1PHly6m1DvuBr0dK9WgNA2lrcOvEcjHuk
hWH6BYcPBUNNkGHWgjGwksylmwB1ORHRLDM6KiD2GnstQQNcTwI/jUQUhbKuxmGk
NN/9aA2rWy2Nio+/RPoYrzzhmUu5pazaUFZPKwasS3a2ty7yQKYdF9N9gW5UDE5x
Bsmrg2EHKQ08dJBjcl+GCkI4YOl/hTiS0i9kQi3rnjYMDVJfd3k52vj6PuJ9VvlO
/xT4XVgYmPPsBTKhj7HrwXF5CHBBtR1AcR73X9VViEJzpHiuRheA5XC38TLWUyHK
AvG1SBIilMFVslHdRvLfadVBNyIdRVT2f7nzRryMwD6BVcjDALhc73KNmjxyNeuI
YYmhPJ+Nd0GinqGUKVI2fL2YLSqNYtxkRkbtMC9216CFmHcCEWWiHxTAWpPduvZQ
+MNWd2DnVLVY/Vw4/rMyMAx0ii1qfpUvbEydKQzbrDGx4N6huH1cKOqXjvG8/fON
FFOmjheGf/GGlMOoKLg07R/Iavp7bxl1yMI9iJoqjaRkfGBe5J5tCLQNaqycLh9G
bmHdbQk4vPjJwLA7nXuUnM+6LygSpFV8i6fHSeXJN86OMJTapwpIcrDVr2WueSt4
2NL5AvfYU2q0NDOlx3RA/AHCHbvHbvjhFuMXjxOnYGubJeTgPp7hLhd8myibhq6h
dmVcNnYPlluSwWCv0Xom00Qzdg0R6M2AadrioXUmNCy6eA5QL0xp7Y57xnCOMbkG
FI7tzWKKyfjli69XAUgl9SPxg+C9uqM6r7WGkJDkSstcv5oVQbrG2JSn5HrrYLOw
XRzaIwT3oVj2OgQJ33JwrTROl0/1e9HzDsZWVR/HoVbFHntlUvn+oZYHjz3c9uxH
TMdlgUhJgOPPekEXGtkfR3K9jgb0iFpCSD08XJksDd5H5+Pbwq5NJTx91sKGzE4e
rqbxFhxjAG98x2kBtQtfAkqQfODf1XxPa3SEDWKNrOMecHqaRRbR+LxoCZuQurAV
NQNKVoSrAyQJlZl3qMtT0lJ91iJmd5kbE4i8OR5R54kHPDV9HtQBREcqh1Tj/gJM
xXGt9lElgefRXuCf7YxuoYErn9rnLCjr8awmWBVlAelcZvYRRYtQqGoU7tWNrX4U
omlrwk03MnxUeMCe6FfJFs1mHiZ/BwTD+6uO/YUBsDB1d/iG37G7a1eYAJ4yT9r3
/uTYVZ0bz0xvp52jsNNA+cy6GIxTMmyVOX9h7N8C8GzHWci1JisiQxRNoD99Vn7v
jVa5X6d+XGqy4PN6AbnK66NfBD6T2f6uPiufjniRcGn9tHMCDNpb0oFRaax/mORy
x6RvvsBDHqYBoNWTSSlECx3KJBIVenm5ktJaIocW+hVLdD5sF+eUPVVh4mwyFX+F
FA8iNvOdf4aJZztD1CwBSTCCCfgZasKcwtI4JK8VkpKHbB3Z6OB3bZhFq6wjGBKY
vnbu9MYTq0aXMEAgE0D4QI46rSYnwugXVDT7yfMlJcs0kNoiPj7ZYezPD9mcDwFq
Px5jMyON4WK2GtZ/rNVT9lZ52sBJ9lO32oxjouy6tJcgo8hHX8Gwhp/aXuY0gvTw
mGrZdtbJgd4cuH3C15hvEPMacIrCiRpULM7PISFtGrO+03W4pxFP4gaXvvroefiG
yrenl7fuQkyuwrxqz4o4bhgcg8p/aAEUjUV2CFKLQiwCkWLRcU0i0dHW/tfTo7g0
9cDgzZ4U22R67sQoMwvlxA/G1Sz7WHS3CyQIX9gY/9pAoj1ZpQ5L7VXFuO03hrb9
OnC+zWLN18uZo32Jzw8jQADARk0PIW6CRdZbJkyFqiRdPTnzQuc4shR+b8I7ZduE
Bm5ZpqypxSjwq895nPzRmDrNqYEtxLeySap4rYPyq1C7tDocdUYwKo09ogj7NeUJ
TNSrLJ61SDddETlaZ6fcvKqYScdNOLcxLfOUqvF4sAC9OBYHDW5OJpsIbt59p2Ps
RJsXQIsKlObva8QsJbtwfUZOOt7WtOrazGZ1t7gI5IW309qD/y2bJlaI7HyrJJsA
o2tiaaflzyLVM9FzINDowaHVvBt2p5gAlQUoG4QQgXq2KfrV7U3pVvii3qICwCV9
dO4KVX23/Q/FjzYrsXQP6xaief5a3tzhJBbUDmCNA2R+8q+HenaN00g3xFYo7cMd
15xga1sZkmtnzMTfFgcFGxZ2LXa+P1HdnqFKPgU2CSBU65+jZv+53ntdHOu91P3p
INHLKiTNKQzI6IsMHYTqeoVb+qsj5ldV/7rVGWrpHN/Omzh9J3sA/GEa8X8qyWPu
1AtplUVqhpniDZfW2tZGz37mCeE1yvNm442wuZdHz5VSMHZnmMeQbkVMTuI9uJAj
UyaXTyJothONKQUJbOcc4E07RsqmjVOIDtMAJTccyBbDuTTk/wXQgVLf3PWxVWOD
Q6sQbvQ2pr8zWIESrCtKFDt4a1+CcXjMkPDvo6d7vrAufrBp/nfZOHnxoZXHrkGO
VZkX58K8cvedBC5pLU5QlioIfb7um4zDX+OWTABbZzYQCJJ/DMDJDQIeTZOd7YSG
atnTEKef8ez/x6+AKTpml4uSE+lEqSlPbOL3C09nFnUqiTvg39kL+qMFxd6CQuPL
6Okoir3pcXyrq2w3Cv18UKtDhGHp5oiU5+31qN6063JRCy3bq1WN6hZRyb6NHSYg
RigLVszodRcQxOp+Zfwurf31BHXlCS5V4PHf39ms84+K7uL+i9sw+cNlmVVmieQs
bRxKrFb4EhtoL5/zV9qT+1P6jrH5hwmirfRGKZjfpO7RH7eDAEkKFt4XJnMGkIiD
unTtHTZ7qUs/lse9VmcueBqvwNrB7LlwOLEMldA4+97Ptcece4RPac/E+2chXkSa
fnR43tJ1AuFlG2TmIGC/JI4d+Qi/6hR0wmemJPpPqbEqy6bt9AucCIg/yoShesLl
4zMttheox+dXnb+50MV+CiD/fm5GyQGCHqIrhUtYvEB++w2TDNkMN5Ob3fkX5xHv
3Br/2ZP/7+XbZtsU1w1o/nb/4RmHCdGK4BIz6DkWrZ7Vd9lEczDpJkvWEiWd6mvG
DLYc+lOukQUEMDkAMHa7R8aP02HZdF0hIzXlgcPPYt3cfJ9Fv26iE1yWdrTi6rZU
Wv0w95B+MAward/NdtPP7zvWR/sc9khaQAgVUVMsEbyJWyDDBtpjw8Jj1sn7cZZ6
1jg1Tubr1EKfiutMln8fCnxJLQVcC7AictUwCyoV6K/pN3+jfOj64NviTqpfcWYC
2cM9rTCumruWesGIT6Yo76ot7w0MaKjCmi02fJUxbauIS9lvrQxqvIEg1vetpeQm
vqHSlP3HxzFOxnKvz1b1vt5K5/jX2qf1kT0PayNX+69Y0LVabx8uxLDq7vSggVBf
Wo6fVB//+PCI4RWFIWqp8qQ8jUYj+lpF1eliIqA4Tk6G6/yretCWFSNL1XJe4gns
/M4Vm1q9rXKz2GLKUjdy66V/jWoIjMtB3wfCOMF9PKghC4aI64pg/vbTt2d5498E
MLvgrppgdovtPJEW/0iGFlxwdBWCQVYRFO4pxe8UHIZOjaC4GLiRaf+pG+FNuf63
cdR7Ce3rQBslD6Tx6vIH1SinVltAe2lGJJxMdAqD5VMzbcbSRouNTV0+v8Jcer68
WNEHQwjXk8LRtJzzwIaTjv5YGFC6yN8MlMjRuH+0oGF7NnG1mjWgg6LB8Qn9WMUQ
5c0P/KEMch7KEkQ0TV0QdTklmRB/+NJkkALQOQwPqglfyJv6tYmRw1wRd4lP1LAG
aN6jHWBubHEdB6ZpJwVTiPIEaoiu9jvqPjzzlwq5/CVUeVhbsACpAECldFsdpdr4
uEr7DPFWK/2rpAYBzex4iMOcU/vkG7+6DOKCghqGNRgQuQKyC9G26bddQ5sLk0r0
PikzvakDhFN7OtwvPpHvVeAq7vb9KzqfbG8boJ5TUTLbVtS4fJUYrr2POsXVyi6y
xXjuAzXvwMiDEPX7R94E2e6vUxytkRLPtIe767cN7xFU98AUsNnDD1rczeTtI44u
J2WfyXP0mn0KxVbKA6JV/zorC6cPrucM6gmRB7qCVZ4E69SDzAHQO10fE3BttafU
EzJ8z1YRYWgV9vJhSyudvPHAFFwdJqAybkFb15bhMfh9JuIHaaMOf8KP4Cly3MjE
vopdWT2bPZRNlNEPEMrxE1YGMbByyydHPJdNIvW+E0gaiVmicIlzFlmUh1vhvOXt
MoCWAFWhYiZXJPX1UFh1A4eAGMzQJht2Z1ukP4xJNet24RmxXKUG0jyb8YUgJ96J
sEccYzLDmENBneK9W3IM+kJE6g29gjabUai/8mrYptoO55dfKQRq1FNUKS0DrMnf
EVEOtzFPSzI616mutFwUxyA7C68qXCkPy/JmZkbE6wruzvJgVkTJyoYdWVAqvkSC
mAargcfctDpS0iQG/jqEMzfyuvPXjWyo4XmROwhU5zmrN3zzCnA+Wyx++BTmH+H7
Tjn+a/pwy/C8XgPjcOh/OUo0qNOBrE8wQO8fScMW6DsvwAyda9l9GcyN9csuZvpz
Uh9rNNk2y6LrZ7rz/+IIcK3wzjjpMTJbckOYTRrjMlCLzjEjzUrZjBWrHQ8uGQYW
LTGP9Yas6AOq8nngzUBV8za/5Dy2EabWChoX62pbt3FoI26mn9qM9N3B9kaieDsH
I26w2KZNfQyZ6JU01PxP5MozDFbETVyIEBOWC7bSmXnAfOPPK/VjK9Udv+2pTeRY
I9ColbaCYuxitm+uv4IiFIvpqb+e/oRAbrL/SqvhuZQyZawxSXWlCQgzORTR87UC
JfxSrUy779UO2CgKt9huvRANZ+JRr9x/6Sr5D4MpydIalZo1jKw4QavvSbCCVnfU
QzpS/rPJvz8h0q3Rgf0NCJ23zB8A8dsKbJIJC5aNjdPZX3OLiF8GAZMS/sgFfd/r
xbFsMjSaFaHAzGyX7ZUV410dKAshHeGEvAQqLYRUJfB5NitGm+swOpk3GnIk8oGX
i1h7o/NgPHJGbQQSLIYm6dt8efjjp6ftFBtOBJ/9XmlFRiCOLMJvycHKEkzjKsKQ
F69zmJMq5Djj+2dVzt4m9gHS6Yke4E6evX9WSS8NvfckWLnk1JuqlZj6V4YAMU2U
9F3i1o/KFmt7XCKELkB/byMTEDU8cmChgdADWJy1tsfEzy0x+2x2rr0Zb6Yyd9ut
BWElM8CCMGQ+VtAxiB3ZjhzgHLflQwnuB7lKrOVDe0OLBTg6zRD1y2e0HHv0m28S
XmABduwKt37Obdv9ZrYHEFkM6Htc53tQKfUwPVdOdNxSH0o2/0gbsaWzKsos5E43
BSHI6Bt/DQnsb+X3q7fhZf2QzJlbL69KSid+gE5+8p7+PMuNVYJUFv61FJIdEftL
BIpge61ZAw5Lwps91Ocf3rguAgh6KQeRzKsyzxRc79KrGpQvaM4yPLxNNTXLm+DR
Qp/uXcNu2NBJ7MxTBt7BbgdHqIkVFs/f8ocnS/sAcfNF5G9UJB9Z9l3pxDUmbcih
GNZ2CExcgMxcW1wYHZqKkSPShWxpqawdB97lSSv9VeRhV/1wMAIBzZ4iyii8hUHb
W/QhdmaikyFG7BkLqwY15mowGzVVdGOKZ1kCV6t4NUkIBuC1WmPFmRPZnIvoK892
3hxf8bXJdTkvr2n3owliTzDlsMlonqYKrPT/B+GFDphi1WvTw6nx8JKrbqdcC8Im
ImhmS7DLjXQ9takPTXS30ESufP7YfTVald7+EeV+FBV0DqG9oSiIqLVf1LCfZ9Z9
GyIU3XHXPMd4n/dpvLYKNeLstEDBqHRJ160+tFdQeLdugr+Gg5CpG7wTktbgj0Kv
BYIjEBoEWtn8nX/9ZjGxErzj9UrisSvLICVVciMixZSi1AHlP0YFwRJqwL3HLdlk
psfJBsqEvHP4jN1+SLoBwnz12ckDh6eowsihVodfXQr1JHBfFHK3MK69BZDBov38
vdqeFTobINsGLenDGpEU6ZE/jBe/pX5FQYsbvTq0NJ1zxZeM9lxBxQCFx22emRrr
1PEypsr5XCgdW3V91ncDTJFRHxge4JUC6NuWX9NqR9qB48ZVzR7375wphe5Vn/aO
WP3ZHRcSHrlRRFW4ltf8fllG6X5nxasQ4xGWnlYZyxp8SjFh6Ev5USlzXi10JiSz
7Y1E1rsWHiKOJGqDPQyEbCLKqbsa1X6wbWXdN/CtQcjrUfyblNzmu34axqB7oTvo
yG69zFZUImzLVgxx6278jAM+DLYtZXR3+euPOm4bCFIZbvaMwivr8zFBbfgLABzo
Fm+LaYz4uynyyv/hiEcZvwgBGQG9+9R6eZ4UI0N36CZY72js1WQf9jv2GR673ZNi
BLudSqyqaU8VHt0A71M+mdoxewdSzsLRgpg2y7vEnxmaFzQ2YcyZraKt7J7RwL/s
/Le9HS+nERGqNE81pRfYspffSnkTBfeKaTXD4S9kdrCkizt2M4ONj9gWtmp4tY3h
pHsjA55F6yU7qiEGG2EmYomlGFRQRWqbsaA4gUFuZOmR87orcoTOOQcNlMy/MPHk
+3p3XNqv5laW54wo/U/Pth3mZ/vSwZwZqYQ9Ror3R1g3xouQ+/KD8qc7SNHkzYHb
lTjjvsHB6qXV4DHFa0tZGobbTl9H/6AlVdlI4N+zQRSBrFeJUSjRGgI1dQ7jZ+P1
u1isJmClL0lu1CbBAhW61n81VyTvZPpBUGVAAMWe+OTQ1SdBk+wgPWeIeVS7YZf3
QlMZf93eW44kuueQohOd5qZ39yIpi3m0KhVwKGK5M3o440LcVX3zL0U1FiHeMCyq
t99GTI2EzZbAREi6nQlLxyrEEZuAu3qZTCA9TctuCMDNpPUD93oyiIMtzJz3eaQw
z9vQJxbXCfuzqMr+GJmTWQelzWWpapHu3K3rdsEKfGGAGsz74TGdtf6NJ/72nqbg
z7lHBs/MSz6j8bFAh750m8wFJkfb1CXeJzSc0LA12QyVCvvwvX4nRLuyMwHmP7uA
N1tVHujt9OcL4uRCgSr6b4LtfqZ9cWaty68Fkbg03dNSIRJx6/zWX3UcNsM9XnkB
gc8cB25CXdUGDkgInBR7bB6nc7yr/3Gct/dPUHbfNfO6+wFKYb78Qxz02iHhZoIO
ktv4fFRU/HDsYytd+q9sgs5PECN4xoH+J6/kKvLjoUOMutrSdiY9hPjHvkE7QxWj
8Kcgu8YDMiec4sCAJTf2cbqEAp5Cevrw6vooVCRSM2eCqgTaOvrohK2JrSNVBmUB
kvAZcWIrp8tHF9Me9HktJvC2LHXl9lr1QCZjxEI0LuRMbeP+BS8lgCT0yNGAlmDA
VoMACiyraLnySbshuiMiCPRAY7W1WbljN2QiRkRnkrRCiwIPmVPt52MhsOCXVyT3
3FMSdjzhB7dn4rGCFVCdn52JLbvNZhwgVYFby7Ldsqq2IikveFYDxZBDnIQ0IxQk
I8A0/RxAH8XwKnhkZ9xzJBg4t69+w1K6aG8pbVkrePymEK6/BmWHQqtYZrqj9qCV
gL+7O/n9iDEmGZ7eHUJwL2ve5Dn64kc6+7Ikmy9F98RfmFz601zVwZtMUZbvEpmd
VwdzkPXKbEohAbb1PHU91genC0JV/qPdrKe2y8bqxdxm+cgDYSAUq55v9WoZzCo2
9IyvW4D6154hjm5zezpSLg2oM3Jsl+FYW6rDBCO2seH9edVjeSrFLJMshGncSepJ
HPlK7ys1w83Jdbbps4CWzNOLx0llNgAp0tbT9t4kYQmnqY+vXUuQPyknuEXMeSIj
CE5d8s1OBmHhs2X+7xAYX7UZl+W6qT7gY2igbyWUdj9JMhfYc4oQ2TTRyNhLpqOO
l+3LrPmU0i7hp+OhEy6hqXwEBiIUOQAinFNBQdZDPUrtIU5dZ88XsU/xpvNH+P3j
kHhB679Dl9Ww7yKV7sO+ZqXOQD0GvACGX3qTwLy4fYP5oMRj/SUxrdGiEzrMVeB8
MWSLhVJgGjhOhmTAjV2JUvDmc7hz7s5j6xEjFcU+8837CUJiCYuPSbNYkGh5/Ec3
LAtRILIFgibNTLEAfXoKD1hdph/V9g166FLGcv+klrsvcaLdoIn6XRtXzWzORvOJ
YImi84tKfBaEMQQS+2kVB7JcbxaAfmGoX3OKcwiS01aQEJfxyq6WGw83qr7ikfLx
/O7Ql+i3hHF7b2brvweEQOHrg27mWIUZHE4aaiOHdwkQFKfMh2S+T67VUsfopycd
jUDF++RxihGoAhn+dTkh4FmTvgj21hLVLlZ1YVnqeiNji006awFVnK0Y5DSxv19t
5MRA4qEo+8u2e+dA6xeog+xDsYFv25Uh23XCWxW7DIA08Hrr6LrTDqJcjB/CfEyt
qC+3xaor2uYQ1fsFfjQZ8jEj7UT9XbHbKqKrfAcaWonpO1SkfXf7HZB+VzlGpEpy
15uei7Fj5oy90UmY1ntorVhjyZLNG+3gnK6DryDijz/g8PAm0v3P7CmY8Mzn7CDz
SVZkXcmOKv0aqb3UAD+XP6uMkYqPWWKAjAh+c1lOvIutqx9ewftkFCe4n6A9PXYP
DO++TTxMpBoejIYOfBVSuAM2NgB19+f2uCruP2XmkL3l/E/+MxZKTv5w2IafCAkV
t3h7w6sBipLZQpUXi0mbp4qto6rOwhd8/QX/gTeALkz5GAT0liYKQEeODiCSsNaX
Bo/ovkx3WhpB9fQV+kNjrDxZ0qmKb4CkLauthCksbcYy9/hAXwTq0Rpz78t0nS93
OIRGyVNIbZ5lirftrWzcp4nSHpqYj0CA+bIIbLc46+cqTpl/PrBwUpPU0RevYSdQ
mYkf+oavoR+XPhz3F/g2mZvsb1PWlH0yB+JXsGQHO8exLhqt49cQz0P3BsKr/ktq
TFchYjI04SUVwYPYrC/9qO3l1YEPG1ualkCGIeiZkTicxJsgxDW+xCxgiZciWm9J
IDZzDrAkwLtdth1AnUZj15KtpL2EXDUN/fanNcFYRU+Nh+DaavZrvDCly88MwIjd
5wnuRlDa4TXbUWzdV4J0yyJuCS1c1NsxIv8qVFpeUPsmb1q+jT5Isnz7kTeID4Q5
9bSNIhn0vcjM4BW8ZI37gcDamgp/BI9ngaoDkKcUSdgQ5dW/lQOz9b1fstEMmzJj
OTOIr1cEMo1+siYYZLMUzcDcDNKElBuApfRwSrf6K3/K/Tzw0iCPmUTbQKCYDKNd
EGZqlK+2rbHBeEUUmCeCEU42RH++/w0BHShrHn8Yux+aXTw532q0PlY5UB2qb8dj
5l/mzoByas1RYUgGp3vZM7TxqFdBc7kyaIBz1/R0hHnxjdjJ0JDC9NGqDTeqc4aC
lOwXxyOGiRnhapdDY81mseQnnILAOO4RS7szWfDOQc77mhk1wzlRe68eQb/fgWlC
qDN4jqLqabCEttGNcxHMEMdCVwiE7Njcc8Merkmq39/TwGJwZzLoll8zC/eZQUb3
/2UVYZsnwrUSissmsws50T1csm4waoAOPP8JOhItlsQEC3a7+FRJoOWXJqVrPitN
ZjOOCVJdI0g5c3545EVMoU6m30d/sF4pCjC8CVbxAtTlMHrPA9XvsHUNzFBIf1M6
7ZiSx6sA/QKAqTu+to0QLRGRqBRsdww7SXI3SBbbHL31w5mUcqRy3JyH9FFuJH69
W3SoZqaLgtyudSP554UPUh4kE5UHdgdcRBAJL7tQD8G0ww9PCoz09bv320zH6gYw
E07wuZtTehod9XaI1b0Nt18SZEXzdBqrcBt/1rBVH2Mx3Hpubu36N2l5g8Vd1w6V
rRKmDh8+HX9r/Si2s8n9Y8bTjSiXmxI7hjjfvIisdRgHbrr4rNGZsabxMtOo3ORm
U5ilF/sNzEXoCAp9VFCyqdIC+I7uKjWw4SFR8yP99K6CL6aV3ieWh7QMyzBSAY3n
NPTrggmur1Zdp5ReV/RKMB/+DCw48LSKNzlbXHf53jSxrOuiy0aE6Le0jznj2Ufj
C1Zf9fMx0F74hjFaxsb+NNPGMz6qt6n7wW+oaO44Ti6zjeT2GHI/9bUv38Y3y7dZ
IzdMeRiEUt/vtAX36cMq6T0HIMWO3uQLkilvtHZjucdoLeqmycciIAWjX6lVALGc
W5PUrpOZZpBx/YTL9j35wYSyrHLb0xJIGW5P3tUJR/sH5ILEeft9VJJCFxrEl2Xm
2QYDedlTxCE+ZTMOI8fXa07NKuZMlUaw6O14blpUpM4cTAOt8UDE/Eke4mH2AY7S
lFiRqdaJc//Z3o0wqoFMXeAdKpvsZc4NcMSeVRVFiAUj6xnpCVU/A2KFuUvuBEeO
y0pW9Gka4o6sY31+whArDs0ccOts54RVLd16dgrsUs/VCc4d62/oertZA4IrZy8T
bW+gLfY4CEayq5+v9xSl7gesv7dcmP+7QjMSPO157KvVMCaKIZEwmZTk1QJbvxwv
n2+q3/zHEDsxpa2Rx6k5J7UbmLFASdztSht5g/RDkf+OEX3Yhfu7r7l9wkdMMn/K
2cKY0Fmuqm+NJWXDtl23rlYrXuNBHF0VfgU845yUATGxSUT2R9AJXXJ3enGKozuW
cJKXI6ik1sJqYX2oDNth2quy1OaNpDwJOs/J0P9avDFJEB6YLgFbPnRPiQPMNysi
w/Nit48iupkuycqlUiRoiXBGzLlpHy3ZcMjjMqN7CDZw/BV25zVJXPj0h2XUMQvu
P5JVzGS6zos7JHp1fTnWZiuu6F35mEQ3qee+vBUlvB0Sbs7lUdX5L3j+/NPSB93X
NJjLliFHPV/oWvKMc04uqmCiSpaV59hHaxhZZQLIpneaGfozdLOW3ng9ertbwXAH
lx7oeA5lxaMl7FBMT96f6adFOpDmVZpiDb+YZlRn1ZBdk4hAr8tXmmVUPgIzbJkE
8ts143mtMNcjrnVTZFrD253rRan5mWxRlu2D9yGV0PnFquYtzzRt66bgzyGtQCEs
/3CMtzkSpGxMhKwox9e8qx9dn8fbzcXxp74uZgbAKhsF+SbQ6NSmfj58iK9Z23at
VcaWZcRuWg9iUbFaNaOdW1gV5+ObYxIk1C55mAVNK9dSTQIzyJBEuQC0+1ll3sAK
cVdH+eKnpIiOmq+TkhNMSkrl6K+ysv8Z+E8upS3JeohxLSgGeKRPu2gf76yGN5dp
rymly/S+UTZjPe1dLhLmtgvbW1fVityDZniPXi7EcpmGSSgB+B8iany8TW7hk0cR
sq8KSpmm2eyHMROiKZURBhHNrW0+xOID25vb44c6+LXEBC3FFSC8yyCqxFlUc8EY
5vhSu/ixCqH+QX+qtFwpvBfjktU29wta/3n+bbSchuwLu3kuKhVEvKIfMy0iI/f/
TqQLsjBuyJhCb2ICn7SOJeoXOSJ7bHBWHRmUX/oExjU+JoKf7LZP34/H4tHBr0so
XrrQTpXVc/m+bIbCkCJxgcUXXmhqIXinPYgRXr/NICoxxIf0u5FohtjjeOSTf729
uuX4dHaX5b4BsPD6HxqfwWRRsOzA3Znyh6eziiXlFCHHAiNaatw3/JKgkw8XG7Qv
A8jBVU4g5/fvrHZ8Gt2k7YV4ycHENDBro3aE1Jrlb5dFuVlbGc97MfS8yHb7JLBx
qFvySKn3WHVn5ALWxHovcwoBCglawL8/FI3r6JK0KtLZQ/yawVS1SdaYkM3iJDn1
cg70Cdbk2+lID3qpSUOaNpH4OfMvE5vVyyz2enC7d5oEVddVh6kKR3fwf83/UTC3
rZnKhCGpGz/81nloff4Wok/YguX/raI7Et7uOv3rghKQwxBmiYacBLMwl9K+qgDV
ZDOYjDdFFcd36mQ0hwEpKNN/24p33/szPGMPNsY2MhgKF5bjNb+crefrw57qWyF3
hj9BMUxTYcrXq24PFhJ3VaVXnOjYdPvwZyewDVj2R00LJ4yikfbRI3Pdak4aY1Sz
PrY7IcjyqvwcRR6OZ1cPa2JkxAxfibsMdYFf+t4jpIiJQzwIKOpASb0Dml76frxS
wA0yJYww/hL78oIfLPv6FqLxUdriGZQiaUJceqiYqp62vM19CKO/svSSdG8aWdPD
KRdIp9Q1JKMWeePBov20Cg7rV5OM9rjnnmspwcE+/gUwL6TsLmfWlla0W8Zpn1i4
EHXPoUQYdQbZz1/Qm8RWck9EV8+tYtLlFNUo2INBLklKS6DOfPYWbLJpE1pL1/Gj
B5vZ7PbI497F4NO97FJPoT+TKDSQk3qpE9F0+4xWR1sp91zCRAK/bynQRhSWR2XY
tvUJriysX9E6TKxc73cfvmSNBhXzMpnGX/cNQW99GAh9SWp3fvGhGJik4A1kD/e3
l7s3mT5mK2BNnxpPS95cGOCqhwaPMzcaKfcDhDsvEgOQwxY5Ip5THQtJSNDMgkxg
X7V5YGn55I4cINvUlYas1clYf8KgoLYXLzAzYCPk+DQDNszE/LZH6kAH77DpRWjH
AZHikGMR8hQCZA5CoHDkZ5OsJj1MtxOfeDpOhhGlSFcOtC+6d4PuMba1vhg81EFn
oq0HNBNZCUA6Na9ZYiMlOGEP81sqzO1XdsbJIDGiH0b+HfgInMrsbV1iJ7oK55l2
9j9zxHNPsXFTg5c91wxjHyy9sDVEsKMYDXm8eFgaKyNHsyFuw1TGZ+Q0xEgQA1Nf
RV3FbTEzXgq0hif+xt4zxTenIp1aWIVzrOXF7gEd5GJSH+kl3SEVxrPwlGG/Qi+F
xriwP3mVDWvhopUdr9wNpA5Jq7DE1K4yC3EzuoCFlT7Nkc+90Zq77r7av7HLss6p
7/JY882O/nJnoi+GCoQVA8sAkpu5il88sapmuX7AXHrbVUgdPZsV8Nk6pT9d4L4s
LvMdZbax46dXHJKSIqh484O8ovP4JAE/y873uox+fzOqMWx2kNtcRTRBr7zkw/rt
JBWUAp9FFJlBJ2/C7VFKPicIynRccydDCkxaP8oSd5wPzB8Xv5kkwvyxJ0aE2k0p
G6AQHHkLBf+LEsE4VRRSaTKW/tnmVxq/o/VfI2yNaXHtWZeVq3EvHQ2b4jqFxBKE
jlYdtmsoE+kv9WMp/Lt97poX5vISB+KPp+bf/TMgbmeKlTTNAe2nOrzVfNkJjWzC
elcLrqKDRF2x28JciVIltTm0cmeYm/yMju9NRJ0+Qcn6oVgCmaDWLVNy50doI/+A
n2icxg9EgchwQIzOmGbDOutdUN181luuypNEE678EAnGNohzuAM7oTPj+t1pBVEm
hHPbwrzzmpc3Wtph/DVWoAdCBXF0fYU6lx+AicKfwPgCY73CSaa9owgOSUyQCcxO
3IvAjS+BrGXOhz/20BSRus2DNqRBvBZAmKuYXZvjvUGmkwwe0lPk7eghbIyHsRDI
9zMfyNUWev3IVWoDgksZmrlH88iyAUOliCqpIIwKjb37lV86ML2I1a6TbzHC8yKM
VPnE3RmJu5+5exqyvmHtfOCoZ4nAi45itCej0nSpM8+hnX4KSBoChGbWZkq6ue5A
Dabw9eZshyPZ/CPXZ1sT1p3oxa8VZnx0RTaknq+Pt7JJvDpUisl2JA9HbvR7fib0
lLdrc+YDlnDCv5zbYifTTcU5uIXL6cV9bFQR8WL0HALxRMi0LSlz9Dysyol2xevm
O0IovwPeY1di4/9Qbyc0EIbRCb7xMl6/3mgMCnV99jHxOPS8TGu3sj7kOCBxTdRG
gwluvKxqfzUHzbIZiYyHNUMVDFIAm07Xfn/jvyZbpjz+lPVnNtnSCdARzwVQH6H/
k7XIcyaQlwCIuL1L2NGYviCfuUAJn4L35a36loghkLbCWCdfdNkZuzImYZR3cBSY
3VD+yYBj9Ab5ADsjTxgM8UT7JZsp6Rf2Eb4w8t8Rx8gFvp2QpKvDDWspoeBHNXrr
Y5bhgX+k9yr4IgMdbM2is8LFUJwuRd0PaG9Wdtv171famj2ZwMnK8G3fsWiaTUkR
4vRs2PdQY8FbBQuXt5Uo7nv3m+x5eSd0YzU0ae86ytiGA3F8l5grDzWwn6OScY5b
GRal01F8EQYwk+756ay3oEl3lGqtLDDyuvj8mUionsbqp3OpEL6N/G3rYNUoCpND
KO8JseVHQp+SVVwFzOSU9y7coASGYwR/Bi7r8ayAfxitsddO4i2cZtvo4x+yRRDr
JZvsy0yiCs+AY18XtTKTOs9sJERmpZWthsVGAp8RQjt1Xp1eIXSAZ8OlnAqsu1Hc
dT5AF3hUS7ikoezuI1tUkpyAwCL/zV7pB1sd+KUdo7ka26+H2k+km0dQVqp4rtUf
hFzX+eKWg7JFh6bv609JDDNxpN86lkke5+qCWFQ53QqkoaV5URcS5w5rG6ARNSqy
lg51kPlDXdKPYJm7ndp3nH1aJH0LLdt4fPU4AkAOLpPCW2plQr2M7EeR1+zx6xq0
DPh2LSjh6KqJxAkR6i/xg2CkRK4Ys2ApwuNFQ0CSVd8abuNOss7mo1Zbg9Mmc6RF
OZ2s528h5s+7XFP+2eKmL7jr88/8NCocc4D9Wv1MVHBkC1jMidkAFOz09jA1IlpQ
mu//9bb2UvTn4EvemElXP1p57Y6eN/M7ArWW8jiMCvVdB/aiZ9dDeuTpCWb3I3gh
qudCbDhdXVX+QpxLu9dkg3Y9u1lo2Y5+psSRj4i3zVd/hGzFXQ32SedTlr7g/nVK
f2IsnGDze/lCpZW+SwAIVM92bK/DoW94VXCh6kvWzUgteTCAS5o3zR1T9SuMDCx1
DNfd7d+RAXEFeF7nqknovt/217yaCOVrh2rOoVAh7xtvCJlD9GCvc2aiRaJnfIRW
HahkyLlokjjhujuMh7ppVmoylIkWfqSaCV0chNxKXaz9dNtqu+8hduo6WDULvO/a
xwCQnYOX5Ky5+8OMIkmwPz5q+v4RsP+16nc/CU5PeZ5PWksnHjwcIO9JMYbMpaxp
DaegPZe+Gq3wW9PbxzFMxO9ZRtGiVE3wSJHE9NZkYYZWZTNVUzXv9dhcNhb5XChn
hZoeSXfC6F2LtBTKKqduM2wzwgFHuNZzmvQxgukGXJgDsmBHgTW9q0pT/3qBjYv6
IwPOub4Mcu4C/4UIOqueo6w9NEaUetX8sddu+cs92Oz++Kqw+c5cQ6Zuo835x9NR
69pcpJTRhqx4qI2MV5ZheG1Jg0gpRFOIbc5jnLM6bliBMOtlGu+BN5ZkDf9NCeXJ
ZtwSMwIqfwCqXeXulkY0nxjxpWlVSPLsWf5PEoQ6mOoV0FeJIF6YSIdB8jTHUuOb
X8/EuTiiH/JW0GnqePV7ZWgko+FnveYpxbaq3pG4fgg0oEgLE+BEXa85mTY9T/LN
7b8cW37YCFad0QItq9GIub8yrEzc6a4mMaZXxaeBduFnEZpmjeWM+W3cuppHSKho
c1UZDa/BAT5Tf9YkfSMyXrb8B2w1henqVv/z83UwNb+Jh+ddjeyUyEz0a6thVdOD
5KJRHWkPWwYTSbIEQbYFvG9oRj3IrrFWQjAJ4s2yTJmkJf3+wBkWRW1cvb/ViAzC
klKBl/5TAdPGv6Sqio+v2IA7dKCgOaXEzs1accFW9u/5AcDSVwiCEgBalWMGioB7
kKolRVbq0mnM8uxocA+JWiBNm75bl57uTbNY3ziAOaJj/cS7vnZ0r5zf6pFnxjFI
iCEBpr0k0LDrx3AfUaORxTa+xD974Z8sbk3sqbRt8qa7Rj6yQfR0JyK6szao5PG2
IhnRNp8TfasY6ux98e7lJPqqaLRah9B5rmqe+Mk/yT4Zxx5gQZPlaS5ogj6PhmmU
VhgNjT3Y11lDbLxlLdOnoAlgvyJfdWvi0Tscar0ytZ5yxBDXapiaQfFdxeo2KrxW
dADDw6i4NZctBGgOq6Cd6YS81nB/yLuwp06gRKoxNO6oLjg8JeJrQ4aXeyOSGJHm
SUmTFhMMSZuiJjcY9/xcoDaxs9r0w0UDCLBfKm/2A5ovlmG9qIVQqkHFVWcCRfKU
4vZkzuJq/31lhXwMXV3GVwuOZLqrpgaE35AuHKSwqsLKo+un3Vg13ULCOHz6N70G
dzrGOocSq+vMZGSsKeR1HPdC/xQ4n5lMlKDquKmghZyBPGWnu7dbljBrHXh5kzls
zOdGp+/CL7HkJJd5Hin19i3bY8agi7RWyXatKUqRydBIqG8KaRcjE+MO74iyBGmj
qHtU2P9pLlZSDMtyA0ZDufxwMWgPxbq2ZrbfbXJ/5Nu2YjcSbtL1NKenGJGZr4i+
2nL1LQQOSHjRapMhEKOQ/RqgQecmWM6Jy5fGVyQTPo70uqK6xaAQaxl5oDiRLQ/I
bFbwJhUIju7TRz9dgrQOZLs/rZG5M0CHAcO2LPkkKDXHQ1S25Y7GQ6VmQWnpdxfV
G9wxP3MNpV2lxtDpdlCwuw/3/yF8R7fSQL2E9XNfDrxhpcdp9LLmTftG5q3QKqQk
hwfGxRxbQWUzJyqLia5NvmZjowke3ElF9oIcsIDEjIxy7OtCBniZFpd4IQeWcKna
r2IobEYyfYokk0tCV2yLswBPRTzt0LYTDzo5lz/GLe0zSURwcH0PR44gmPJm5EgF
EyzPucUDMZAhFUkDxzcAlM9fiFOikoDtSNtP7WapHVLF5Tss7VoFmjwFVbVkH4MU
Ox8+8ge92Kf/90uHnqDKHKNqeP00p41mlmpDcbntCXrl8jKWRLaBMRZ13YoF7ou3
THTWZfZ4ZIJwd1bzoIuIpbhbwfutViQd6D/2IAXOcxpWFdcFp4QM1Hzk7bIo6SF6
3oBD7GBfE7hhm28hXGMkEBV/n3xY4PEk1gkr4nd+qVaY3623sTPE4gwmxQ1RO18g
VO/9xXhd98LeCC1D4glHtl7SmqCuhYNgaRNljJUCKpe9czEH+ZFu2YFiLeis8eRW
bkgGm1ukBSle5THcs2UbpNI2V+ygFpwXtMu1WSBjWbTus+w7bYwzJ3OWHULpQtUI
3RpxchFfy17z5hQzxGHgX94nc6SQJrjWZ2ZpvudNii9wl3SfyQUCTIOrwN9scmq+
QlYgs8jyh4+AreNLZ1YdP1urSTvZGIFsBCKoZo3ETxKYjsXLYMuOo3Sys00CDI9/
w4fXBz1kAjsqzhXFyxFjM2HvzzrAI4CRnoTbuu4nfZcfY/7QDwt/CdX3rfsLAhni
lhAoAS2jSVQizbEqcsLDJzqjUn2K2e4v03KuAEyThnwh6xSOHQhohACPqIPNfcov
s0c9HxJHXiBUsievFiJqTTIfEKyY65IJbTh3C7RAF5Qo7UKoC7W3AAJjtXZ0rKeF
EtYUD5UR5xEnewbzmhgaTscLpdP6wCA9DZhxgg0liaGpG3kbrrxaAGN3Oyud1vkf
ZHELQjd41W/LxGMTMrKjJDmc50h43gbj2swxR7rXy3nWy7kguSS1K/nRZOgAfsGY
mcaZY3fmciGbvwhvSF3BgPPvshs3JGcxY4Y8hBFObxaKiduyJ23l8uLVL5abua2Z
CFlFVaPrtnCYrx0blNrKgpGK7V0kKLli4Tx/QakG6m9XOi3qDJX1k3XipgmLi0nc
w2d3gY5NkdQAxIUkkmYJ6MLpQVtOVyqbggDG/IbLfZQgCMeOnzO52Q7W4fKy93eq
TM+J1H93Y2MHhAUGSJkSI0VQgksGP/7orJoAHUHrfj1ltzN6xWg+lHVlqk0NlolQ
LgNGlaU8bI/MW6u2csK3vG5H2tA223ajDsMnCuKlLh40zzezF2Wj1BBHfY/mXKhX
yfiT4YZubS2g3UzQCMH7u0xQXOjsorf9rYwwJJdmBhE4JOdqkUIdBvd6q8dAlOPd
/D6kuC5NVTBoVjXfh2MjL6VPBwU7aqwDSMQyHpIrz3eCywfVm4aY5PxaIAgQeRlK
ivBfnTsxlVTbflAvdidI4XjxiU/xjmeUQEMcSN5EddS28fk08ehSXlknkFLEdS+h
RpVmwufbSDTtFsNgLLan7ZuzdKARbHMk63XM0Op3IoV9tpyIrSfjkC01F335llfi
O0m2tPnWsKcSEUq/m1bQjC3Fu0DjXxIX8G7GKYY9qPMps/ZyorlKn52g4xf5/UzI
IZ+sXGuVZH7fF7yoEfSnWlza2CEavkGEB1OM5fZqpuLhsk6bDONEio1yuXme0zto
Mt9ZzRaLfErpV7cBUBPUTiloLSLcJmcdYZh2KUdJDFXfMNBgJMEgRE1AFwHrVtCO
EY5vstRhvKlNydJ4mLRdDE+WUty7KK5OP2ZKAuJ4bB7kzywUcQLhugTawIsegGuy
iB/2LtKdSLJHWoDLdHSRZj/GVgG2GhhDPicMedAZTjz8TleFpsLiGpzckP/L8DdO
d0IKag4LAI8R0s+nV2RLZm3YGcHIy8oefcLXtAxc4ws9HJU+xNKMBDLpyCTF5qgz
9SUeHZ+XBGv8q9h35XXzDIjUhEPsYwcLAYugTQ8SylPFKm6FEmTKEyt3IEjiy3VG
1fWXw0cCWYN3O7UrPrId4buYjtBJEoaXoopSahYztv3qH8eNgbHzLw8WnaJlG9It
upz/fVoBeC8WbAm2EJfCD/ZixseF2Pc8k86Xn+Xqw7XkNBhr5MQlo7gqqlyRzHc9
8w5AhTJrSH57+vo8ukMiJ8+59UAFGMHwD6W8qNwtYrlZi8BMW0wOVS/M6FrOELcp
cE7XSzFpT9wTmhPYXqJsG8xVVr9kAS1ojGBpxOV5g3jIkWKY2p0/VDhhDP8X0D9m
MbmQz3XlOv19GZxDneOqZzVVkPe9l2JUxjG+25FA1QUoxHECRmMBwQi/V9NFOO0l
/xT3CrT9eGX7ikUgirWuVAN7zLYBJc1vGKxbmBbwPiPoiWNinRwm419gxNJLE/of
imzS8HN4m8tRa6dY/8qwFzbN5diDR6EJerAY4r8GDv6x9RB0YhfeRu4Jg04+0BEy
aRXUyC9xrPO3wYBit6ry4dHuor/xR4/l4Vi4sc0bG+jlQPpyR2DiNu/Ggs7gCQva
K4Rm0O5XwWe+9G/X+noZU+9UsWYj7CQmWk7wqtSIGX9FblM0cZc0VLbaQ/dEMHZC
yBSguEhwMF0TnJz22ROmrFDREaXaY6AkHogU7rCFAliHjIQ7WUAi26mX0tMY+ND1
2T7q45g52UJE9JVxG+IBtBClo1agkH99fjXU2XCPoSfkZAtY6oqh67aj/QYHIpb+
Q6+OFMa8vKYt0JvfGlgssDx08GbmZXgDoHhhlOVvXzwysfVc0W9E6KBKzMN+Lese
wX9JLJEBbsLlrtKYFycrpsMy+d+GGSOwxd3uDCMA6x+f+3wXPVwUukCkjw4+QZax
Y6f5jTf4cy4bj7pH1cOJN3QkvsAlXw1AOAydN7QvIhbjjeWFOT9YNoH17WL63Itw
SDrRQH412OYDIbDyTB/7cNoETSg9MiQvqaX1ljh9k75FskSL1SImy2m4Jja2ZP0y
FrjgePrdb98amxo4gsevZdBgzdSHy2U1/X+dYcNwqpgE4CJCvkFk6wdiQs4EHyqf
VK+rOEQH15bxc70s1G229T6pEWNLYLrVOSza9Lpfo1wrh+aUeMKeBvmK+67k03Ls
qF5cVM0RBlVUjIU2X/Lr1vKQw889tsaGtwIrwQ+dvhbH1s5owLmISN8cqolZvej3
EUjHutXkdMjCS8XswIMKsg5FEqOVnoBf1YBl+rjnPDcwQoKFrtwooI0cSyncH1xq
pFheLWQH8C0LRpFQZ3FICoGNG0rJ/K/fr8GIpcZasLOf1aWSM6SkNApxWYjnj+Yc
4GSwV7Se66k0eupa2UETG1ZTm06yLUlKkgDQ32ADcBZkLQ8YbzdX/1yTD7zGIzup
c3NI9DRbhZLOSxa4Jh3boMa0yOWmTstJF57VG1g+K1EtTLWntMK7wdz+n0ebstab
ng8GAWV54OueJDtm/rk64wupWFLy5qKi5H6Sf025urzCXEY/SFLU6bJnqqe7UfMw
8UPjSS0DUnBJkDZNHY7IBx+Ajyrg84X+dcBQxqpYqGhncFmvBkBztoKard3IqEqP
8uaa68LO+g6w+P9vfhTtnD+pOmOx6BApNws+XGh2KBGYXUQML9MVeIFoyJltzYG5
0waDZp9Z0eVEicidgtykAieyXNevn4wXSGauk7NhuT/Nx42MFu6PEpsW+xEll8O+
52J/V+XU4PjL8KaTiFfVWtQ6Cqo8Gt4H+/FMJT4R4ULjsv/lKzsjL+xPs0WTusnD
tNSql1VyKYhcBw8BKi7bkGLtgj4+O5mv+XtNdzkZZAp9lIv5VUGPlijyiaZyNTOC
vq1Cgk7G/xKBctZRyROrs2yVVONgs1pEDaAjpGJ0Dj8iBmc16DdVdQv4PNimaxlO
kGI6LEZI9/Z7qTVP7yYi5khPIhTlOXOmdFiIIdPxdrGCjll0N6aDmAOJ7n/26nG9
sc6x9H5vY5myIIcBD5M0t/lAWFwSVz4TQMHOTtkxlVLwCO6rdt/prtMSXdLiz2CJ
a7n+5U3ouPxGVMxkHNrdVruOjO1Mar0AAzTbA7YXLM17bS10yoUuSrt5Z+nGijjC
6qbds/B37TzeKaBVdFsS47yNgp+1AEZSN7sYuELJzA8dvrzKk3zOcxFLvYTV0wLm
6Q3s6zzynAALy+uFou9VhPjfeqI9dPtNTEsKqPEG2GgihRJL7omfSWsEdzEouNQn
W4SwigHm7A7PmLZ1H8XWfFsdGAIKnClbHvxomWbIPAhlw4Kse6N7qwduOgOzQq8V
vqEDBVBGRD32BMIi8efqzlr4+Yl79c10oPI+a5nuQBSJwND7fkq6l6PhCoTlqGvZ
3UF/p5XoyCbHVgsQhkdc9iwmK4wuGzKe1TVKKSPQhQ3iNLCG9V2SfWOpVc5orEWJ
Z+DaV/bXEXf9YFuf4WTZhltWs5bTcXe17Y77zNx/vokFOoXQDzeNUqU+uArohduP
Q2uWjNLTgf10SlNvw0ybSDUS3iPuBvHiY4CRW+cSSl+h52M0TVqf9BZ6u1eM7f2o
OlooBL7uvDeoPLk+Y22NK6acbfFMiYoVczu222W6pHf1cfNKY5+sbOzRrOK7gweH
EPNR1BktCdCsnUPSUXnHCmTC3J4hBT/Tl9K7EciygIo3xCec/9uSDuRfTypwOwIu
2dVoHlk+z/tX+LYK/bHfFKOklndO6v2EjoC5CLtDb8HaVBfJRVOK63Qn5Cd8SPVX
E098Crvz30dGtl6oL+khCAvFt0t/05+3O9MJps4QMrqGxAPS8O3/Jd713HIUoKvl
+NxFGKcFDxmAWFUgVMrSUTxa35Ed0oO+BGKxtES/xcGaJ/AA0Ff7+iWAA+9WA9hk
gXwlxcPcT76JPb99XThpwomvZVVLSkQOYQ5QsbMg4D0ZdsZckTtBH1Wlah5PjRU7
RDGljp0ttiFCHpamwlrmpGm2oRQ/OnL3W+MTpFpZlEnuBrM4CPPLKXJKb/IQB7dd
GAYZeGgiORiETPpI1BfInmb0fbTb41IywZ+j2llzhPLAy3wYsFfgmRq5zoYbUCsk
leyLbxWIJ3O/QaPtlBQg4XogscT3yh6WTEEozp+V3DBDZj1ES7Y1YcfIKm1jHG57
7S5UaNql3eDGvwKB8Q02I+hdopo8g38LXUdBQMoZK/aBkSaQAOD5hKD4DZhpl4MC
2wrO13U9/gZzC9qJ+dFWw8L3qdsuAqw0y0mxn89bn1pMTGO2Z4HTWJsDjttzUesl
iKBTg6NtUY0ek3nmNc2Gj75gyzS7mj73ZWdmJg9aLGBH169GT3dRZd1tx1y5Txmq
PzPYZPZ2kvWJ3gLcRr0EvsvFTU+NA4ZnJD5WuQG3Ybr9jUEe9aznmoKbqLdK0dVb
Z0Fp7c/hoKtvH43Sf8zqLW0LTZdkTLk9755L7d5G7HEQSOhJAfsTtJKS5Dsrbso+
iW10loWLGNhfm1XRk1ZQtlAkBnHBS3W9cL0+DHhmnIg7LwD1SlcK6AcXMlQOo3wM
ElUppweFxS6h/AiboxrmBiSNSkhnhA7izNjPNEw/3gMdtzgtURemuZndzUYBpSCO
ua8/wf2FtPxuoom0k4nKTVoB2aewi9z1aRQWeEUTIewQHJPpQEJogEd8u3KgT/le
+ncTt857maFmdQv5AMk7kvciXortIp7br1TllnWV8rsPhY2BORUiDjAYWn7UAll8
XDycCSsLai+gyEazRZS0FDtingRjj49rZ3dBSAOvachpBzduZgEncI/EkvNhOOA5
fE1JdeJBT72D+hBHCsHGfw1mxnWUqGnkwBmyzYU/dUwJo2X5OTh9s1Vek5kaXsCI
k1p0W42c+UxUNi5mwGmhJiWxcpKbETjRDskWGDYGRfEJCu2Nd/W/GyJFf2k1eKoR
DgeL0GtkQm33ZSHc97++CpRfaubvZkUsrF7NYpbuOd29x3gbSgY/FMF9JfzSj7bR
dTHaxSXjVOhl8ic5NO4ss3FimIBGH9Ug8x9ah/MI0WpwpsOLAQ+y1Meyq0deD4J5
RAxvtS8Uf28BQq0sApdelB3mbtISYY3Tw83cwYXa6IpTlFhKDzJArNRr1WJ/P/in
dQZ/R9NKyCG4I+wbSMpjC6/NBY5m/AUi9EQtT2G/8f+ugd+UjAiN+2uhJgYpcraV
ddIOcOc+S+AtCb3CZf8wU1OgHgEBnHIkfISsTOgHziFJ2Y9t6rYNJAO6OwU2GmPO
bdYIIqCO7ICACaauU/NDsvBqw+53JRgvJAZJZRUCA+5nj9y3/RvYtVDTerGvqxUW
mIXYIYPqNVLjWst4sHMuMh74T6jiwnPOtVaxSmrAnGo/89E5OeVNWfLA22Ne95Zh
/NGle0Ej+sbUZDSeZwiC98CgmI+Lf38EGaImDd/IE4d7qK3erXocKtJc+1NuDTYb
FdiY6qlzCamj+YgNYiBve0q7npGAc/nYt/M0ZGOKkBzYQJ5WkuZ+auSPjjQZxsZ4
QgGmthVWN71N6peneJrTER5f5vrMU3U4tS0ioUq/gr65t1pNLd1Y1BSP1bwOTcTf
FpnlqRaUR0K8R6vxt7Qf4GmY4vmn72Uvt7+8Y9nim5KkoxEpzv7C/paPYek8bokL
90YfvZH4IFqHG8yBg0gfuZ1CiKvP7Tt1fE7SI8rbsoD+qUJYVOmpfJCtLfLHiEAa
eMKxECftJiy3pg8fVG2JKOxoxv2E6BHRELwarmFIV5fPF5PvFdSrk2EPQVCe8Vtn
EpBP1E2COKNXTvfsSdkgaJoBaguRgFm/yYiibZWaAxPCrkLmhIzcUf6d+b7ql+yQ
pMrv4Kt8KmzsiNGrpGzc862UCO+yBEOGBpl6VbDQCKLi832cM/+Okqjzz1eHbTea
5rlWabg49SY6+sor4LIjO6tOPtNit0yGWeBYYCrYdSRFvOh4CplojiYDNYovGJha
VFQYVrLX16Sf1vJQPaR+F7VALsMSKPB4auQxhVPMz306hdJIDEf8yzlIWMf7Xo9j
NxNEEBId/2zBNnKLQRFQuoRDTaZAu2GMFZs8HAFN/tahjdk8LGfo7zYIALmrvGZP
qPzIimjSh3ek824qzdXAS2NV7VkxTxSiy/jZzzsG6Q8AjZRiZqZf7DE+R3ATOVjC
Ye5We7x6jKsTOQIXpbY4VLU3ln9MWM+12MLjcRyX1053KHY7zgi9Av4FbngHdL20
y8zVjVaZvUkV/3uPUr8SyHMmLye5XVCcZSlZBov7OWYOnZc84MotTkLu/NbvM9VQ
kLcH4L/4sYEsv/sFstzpo+UdIGC9OWcxsWIHvbcGRt9bMQL3gvptne0ZuBd64uuU
hV1neumcU5FDY7CUUrQ3ESPw2d6ZR/trkJaGe05Eu7tliqv/knNpiQkib0lgem4f
z7PK6jAJf1DqpLvWcXkbYvuxT0dc2RwTLYBG/Mp1RBWqZnQaETgMWOHum+S+8zKP
V/vHAfBLWAQMkX7842xEnfS/rCG3kF8u67meJPh0ujbrmJD/AF4cPHTviUEwhci/
hgYSAti6oBVnXeBN0xtQkbbGol+S8JKIrib258d55iHr/KXrFKp/sb5m4rLCkLdB
0YOExLI/2IJH23m2+ylD0c8kdW1cx0yccvWtigVDil1Hr0eyzWkIYZQ2rclwgHhj
/rLxjSnMna2SuuRrzQUu9x5YLFq4K7+wUJ1vb6STcFQe+BSshjKFb9l3CA1F0lVJ
MkT+/FTFDu+MDCqPU4d1Ks4MNRMhn+bMDsTKe/FFCKXfAS4oebrBiHp+OtzR+zwr
FJYrmHeYUGFHALSkdpmOt1R1Ly9tmUQB9LxR6s8hDRL79W3xOhZYtgNYZrvUgHDK
wYAW8m0acgqzjIuQ44w2K8FOJQDru8QTSFEqGRHfA3HA/kkMAi3SWr6L31SN8KSu
Z9wHPYS+Y3esu6Z9e5602bA+b54d7i3QLuxtVmAZ1nvJ7afXQl6lXAuQvwnGozcs
MxWZ0b4uZoV//K8UxIqSddan3Ps1bAtwuW0QUvsdVWYEFc8uzJFQjoUZJYfPdw5Z
Upy+lbGZC5TiJU6sbi2fnfoaw/Yd4IMDCcMLDf1Y0imeobVeGOKGNtgNZekhHabw
au4chYX623UUB6Q3u11SL9q+MDEbOa1KRhAdi9+zhqeRJMHfROz+GtxWV2xXSS0z
8cq7hENdSoI/+Aup4O05wHnJWP/9aupTmR2NF13F+dTGJRZFSpnWlasgbhq0H67c
tgCo93f82xhbqv3z8+1KuUJS5+Q3UVJcNU6uRozCN8f6e2q2lf8tor5hEfU0wnLz
b7WLO75slKSe/ofzIhAruBBe5KpwEnoGH9EQ0wEU3egEUU2IYw061odsxzaMotBK
AEAzbbtrBh3Rlk7dNOOpBdKuT9bLToJpbMQLejRaanc2PH7/1IonlRnEtZYItTkO
9nEytQ9Q33ffJbN+8r32sXweI5CQU/2CKZJuvJTxTOiEma3j9Qw51tKl1WHcBZi7
UTl02LKiHDMGGPyLi7YDafDkoOIqJe5BA812+tf/QVV15oG5illtO0mwE3dfY4Iw
7JzhpxskvSGLYClc5ustvzO6K50Shfh2wnI75M228+fteShb4kGpNbQrLXlkU+u5
HGApfo6NHUPhpFW6+X5CIpdVmT76cWv6nCua6zEk9P1+jRnEnotjx17CoqdDWioR
Wg4cX2G8/O55r0PBtGHFPzQkahKj3MYVRmWiFN1wsxfeics4NQYG/WE6LRb6gCxd
VnTa6lK3V9PncgPvHdqUPDn2mjOpv+HfJyowKRxh5Cc/FRywAmZM4WCC0UULBD5Q
eO/RDN/ELD9W2OhLrJjZ1qVlO/4N0somxhQLxrWy4KEn4M+tWWjbxO6i8nk4u8SB
4GU5CXnC9Rg4ag3j9f02SqXDGdi8YCFW5KWPfb637lM1n6R2CY50qP7fd0a8M8JU
sdJ9dv1VdTOCIlnDn+j+sWw7fKucze+RGEYof5JrddYh1qZT9c7TwGyEQyd52fa/
Es+R6FO10kAtmbEsCsjOmXFTbIviLGisL+iEuFF5aIP3mk7JGElMA+FQg4OHcTBq
xpAxXKlPEZL7RdmiInbwZC6vuFnUEL+95i3LQzhKlYkDVzK1+7J5d2jcqTUzHSlY
RvGtQOPFOPeHKi6cavPMc1+mpOLtsBkuvbT5Jqqq3eCVmY1luZIUaKHC69Y5WDCy
4s86iBbnCIjbG2LsGe+qy+YhrXhegDVmwCWfSVW7g6duVkuN9crOd05htIabk0uf
jdb5JH7YucJ8+N1biyNZ+9o9nTePkwMG+Xe0y+Fq0L9pJAfCQPGcxPf3nHvN1iZx
reSCNyMowiMdMKpSu2aMTHQVeXDYrl3kaiRJoXM/kYZyAOLwjEjrtpkKz9JK5YWV
41zUkf5ixEvKizczpKUVUvLaHmbOl2C3/YTn8Ek4NniZA8hJb/K0ZBKLIJWoxzQ0
uW1Gn0JgkgB8vuVybPOyPI6yFGo75KX/ik2rgGl6DMDbtyRJpyFtdBWZZXoATsc7
wkn+uT0VPhWHjNow2RPTbufTMvG3yxlqpgngsWLJ5i+JhjrRbM70ZCvkuQMKDUKe
qhOjYgfFvwd63onmCyU/HsY7Cn9YgzX2ek8nM1P6yOig8NCbZYfygwhDmqEoTgKi
Qqye3ye+Cy3/N1g8VfmMhpHpK9MZpd+G4fBf4xy8NIXGP6UFu7LQro7bEyzh0j7t
uXHlu+5f9XFnYl4J405sZQuHzSJ0tDQpQX/Gxc6s5FjBsIjmyptki9Ql3ysORP5a
xhwJSYPOgjWPbB0SWJEmu80bDah3JquCgqMDMgNmtcT/YcNQzXKiT+T4R+vQMXyR
U4G8j47widEUMmnld+YgP3T1MUXvZ0rJpM+ZQFHG9PQ4j+uu9qMoOfg6r6p3Q1U7
kUc+0/oVuzk2nGkrjuoCWChkQCIFgWBIBJu3NPfqQFMD7olJXuXtrtLa9Jbwu1Xu
gohm1/2zEPUWJBTIH4k1eRGQCugL4NXh/Wu3soHxk/JI8o4Tr8snRHpk3s6bQh4B
eKN+eED4eO9okpocNCTDiE1SrS0lzwCHVu8lla4Df7V/Xe5UrFVSYPajUWsVguee
lQOHPymYhQSxAhdUYEHFA1Ogx3u8Mm5FtIVvJeiWrtWsxBwr4PcgQ4bzNa4jPuBY
/sTaqv370NhCcq9EdEWvUbnFLbuOHyiZDBdBgz4RGisu4KB1n63pahG8NollXt5+
gSTUVknNg10iF+FDIox8f4kOasxLODgvtGgHvPmT/2gRZiqEaj70nKIhxCmwP4a7
vJim24Qko6Ml5vKqq2jXQWHFm6IyDShAZ0IY4xyrfqDzw0lGo5C/YyQ4FXxp0EbU
xu3lxSvG2o2EORLuKbaDzIhCfIbVvvqYvIIPTiFlBzxnNYGw3zaxprRXLe6oqjuT
HS8AmzG4gjf8koiSaiXYhz8CL0o7txtSIqPYVUpvV8N+Wn/AKEFU0klol87Qbttp
mjAxwD4vDIqOiij7Rdm8iN78IL62+2Vt8wgQEu99O6l0ZC8IcEGKbVH/q14bzNy6
j8LNDPCmr+fUQxtw0GQx+NwjMwd77NJuIt+TeM8wtlU6YI/xnlYLu0RsAx83NYZG
EDgk6ETILCPBPzVHg4CRavMsVmenKSKMBl0Fnl1ItcIlWnaERfJr0PnH+xhPS8Ap
ajwP63GVYx2dUtV0kYPbV6eahwHtZZVZ/Mf/VYmdYq0I9sfUcDtfPYHmqJ7Bo+pw
AZbtDa4Fi4USWEq+sArR7anXLeIM1qk4YltJX8Ia2/OUaOLRnQ2O+UpqP+Z1iNRU
92dDQRHPDQ+v2dh8zgWyOftOf9l8iYweTBhSixkRzFSOuplygdH3k/5tPNoTqQSf
jU0mHcKgiQauNi4H/fZ8JbkyYzJ2i5q1O6gOI4Uk8EKYPcDl00wtgW6rxgH+7Kxf
2xreuAAFvDrTefWkeLkJaAFVucJG9B7KAnLMcFoZ+v6l5Wlys3pIEE9F95zzGroB
Z049cxtodQZFyIQP/Wz0kv5e1FfUrE2UxBUOKGk+FQjBDq5keof40Ep42VT4jFOQ
lT1anK9yAeoDItmDZvofDDE8GVRgPvgoDCI7B1QojRFL/hJPE357J6xekiPcVkzo
ugM/ZD7rcSnQp5SsCgFFQ1Mz2/HJ5mksS2Enqed3ZA7RBaEpEPnx4BsErjgpWHyj
R/f0t4bloKwVJEQAnBeuySXQcKJJwf9Eu7eYnecZYFXWVCX/nW1cBnufmfDail0W
9PvB+0tDV4L5qVLialHf/aQMP7ZcVnKl/gGqQ5TzcTI+TIoGf7c/DqT+3ruHZCRP
VFpPh8h3/qsVFUkSBqRe8JjDhiqoTWwKhqpVqJ4xysN18FObBxO2++17dd/OXnaX
7prlXOqvkHLhEozNp4iMmC0Xt6ESPjf1Nh+JTBt6opP68hh6EWgLqZxcmWX5MULR
U+9iX7FFKAI5J/eu9+NzhwH62ju7ptryT3SVyHi9mKLAg/ZMQpL7LolWYQqdmLIC
N6vq3x6ykpxCx+/NAwDd/MNy30ARkmjjhpIemfepyGaPxBt+XHmmK7NxiyLVBp3i
xClAFnVhgBULnA3uXyA1Vs5i53CP87W6FNTgydVqQ5hPBm0xaJmkuro4ObUSg3tl
O+W/Twa6fVflfrwmRj9cf++VTZtVD90rkcaSTSYUKRwCFMgVnBnMZzg3Z3y+Imvh
pmC2g6d62pbNGyneLMKBPm/N2YYNy+ediO6m7fiCtmm9uA0wu1ic4VxLHsOcJn4l
80t0BmVlbHrUIzPEekbacmwvzZsTh7wGoNqn/uKe8kp0YVnJwbJ3Pt2YPflEqht6
ckjZvmM/efJBbS5UAZczaIJ0Oeo1tUIS3OGUwaebDC6omeeN8OV9iOvsxJQY2d4R
+/z+CQJ3gj1f7buOmnf5hBSWOWAkUIzlmnxS5s2CCst8o5zSljHVh631mOClOLaK
CNhqbDw9/O4py7OOWXfMCRjJqE+jE5GcYJ+oG9J+lZUdCoIOPE7/xqDszfFC8+n0
0rXtzkoIQUY0D4liuZAUxv6DZ9IdG4M6ktRUPatKiihq2jpFpav7lOam8VPXcIvQ
8kvTkCPGPRjUfH6BBz0/alHKITaUXuFshCTyA6Io7sYfJqJhncLGsWMz7x+6C0i2
w7eN0xOY6V8m3hLQQb1fZl130AKOTTx1XoaSSHFUQBwUmghMeHF5TGzpJwMU1HDG
WSEA22Av2nYNcCWlnb7YD09tGGbwYU5PvFnKdsQLXHlF+WnzecdK0Iyunb6V3g5L
jl9tjOZP/B77muM0E24qyRcsB08/t1HpX54VQfpKmWsAUyO80Q2zR0SNGrbxKvhW
UtCtoiyvRpycHkGtS5HvxdkEpmKod/N5jR7i+sMQJWmTN2csTNdI0qqXhoRlJ2hp
4+fAaSXTNRz3Ix3ZQBnWQjgc6pP6IfX4q2KNj/o2QFAGkj4BU+V0gRszRTvcraHs
8rhyK1t4H6n1hQyALmj/ddj09AGqYd6yBklrf3MmZXaTlm+f6ZYyKV57uuDci8oZ
srkPH8foxG/aX3Ezv56+l4pccEZpAj3sK4PFeaM1xdqqZ8//XCxSei7OJUGAepu3
1oI+IadNV7cJBP5fKSL3TdQjnUDw18GnYc+lMeo248lI3EvZeS5M8nI+ujAUsJ01
sn2r0/9THOh79Dafazv7AhTdkguUazgifGVJodsTPiX5W4+6jrmqnVOtm+tilQCf
m1T5K2eBb3lLPqJYoFV8jnafxoWLSM1NaRe6HBsU8CbQzeCufDxtY4na/u9Y9bYy
t4l4qixziXhh4E1MZDn0FGHVuIYWiiJAUg5ZgYAfHW1CgzMGMSO6TUVmwr6op3kb
QOC4jr3VmymYFg2qLoLZJA15hCEuNVEgFGAMdT6AwVIVep+JSlnx/QzF/e152Up0
BQP9ONVE1dRUMjThU9QtbhGhMPtbkpucpmJ6hlZntlLY//oI1iB3U7NZVoA7CMi+
6JBXfEdXeZAv7+Ku0SpdIWiyD69VMqvQ5LGkUv6rkRIZRZWShnBZnMUSTOM8wMn3
ffHecEzEU7mt7iSRNqyP+pmhdu0i/wwX0rUQXv8rAsW1DuhDInUkG26gY8Uu7Xf1
JHn1+yw9MNb4qpD1CMOYYtFrY0zrxPgMtbqNt31Dyi3GSCTy1bCqW+lSdU0Drme7
bxpwPTolPJnHzH+WmVkyOzl87SC7KVLswse5IIzcCuhARA0FQO3T8HidprnvRGJO
K4dmKYPLG5FlxoB5fAKtHL1fqJDvfwWSN6YNWv0kjCgZWgPCuxZcqNR0n7plzJEr
vx3YzNLGLCOyupENFIUub73GnhwaHfi0FrDWUSpemhBM7RLY0WaPWMIt2GwAC6B6
2Mg6ljDPqob3gXreWO2MtpgPjU84SFJLGRtndbjJI4S/h33DnNrfV3AAPh5ail0X
z98BUNvOng/b+VE+065NnBI/Go/re0oGKcnPdXsVXDfnXEANRMLIGYh0jwEeNsfd
tE84P3GpSj0HhxwpEI3uYVEpGwGAXmxPLvAHAejDcOLfP2eazIfvjJ1Cw6pOAoMD
svTqLP+8iDVfFtMEzlLIH6PgtIQveLJNayunlLcIE45euDlYTJzas5qQRC8GJrRI
e70KeoOSZP1Pf1VcjjkO8BWz/dUvJlmdOu9pAgPAWwfhBU8gC5VaTt5+JmCdeI9N
0W+7xGHwLF4h0X3hf6L3rEfQlpWeOjiZAm2pS5YctClYSR/Jhx4jW3qBFCU+uyAV
ZcTPhcRDNzFerMbLfWwJwzdym/mCd3YDZCldYONpV21NFLhB7FQF0lB5Be3Z7z77
HVW7erq1za+3XhKj4ku1Mhwsu+2jGZWwOh8oo0pTbZktguLVt+TSknHNAql5FbxO
LH9e/LQwiUCeEwxFl4W3ZZR1RVSo1ueNRXNf0N2/QpdPE/g/yXA/hf0Ta8OPL8pL
H3j7sM4Fz7cRNieJ88ykvJjSCgdOx7VHzYyZLbXLUCUmA+diWgHD9bkPNJ1CTbiz
rnvGP3iblY5FoeBCczD5HRKIeXl24cemwp5jamCLwLl5fjtTb8qY1KEflxBF5h9B
Bav/dj4Qoe8OawHg7UDYfI3eQ7DyNuPounwUbJ4eH3sIAA805lLzqYBf1FTHbcjR
Hr/ppNqFSiHyOa+XC45i3djtjHAuE7Ecq2o0NrBRU1J+cFaJf5iv3VeVr8sGPocX
1SIXNLJRoYlBrxxq0yUkvl9NIOJJIWb7GL2rymsqTJA9Zy6eNpN0TcvsJVXLfWEW
LbbNqLIgF99XgyVuMJUyism/0wEEbsn37YnnmCEf40iXXVgYPOMG0hov5UExOfI8
hJ09fyuNhawoCYFSyEITANEY2FOjlTbZah6FVEQT6CoAO3VU61BY+dLu+gCtFiZA
UqxsQ5szn5xiBZor1Dl0CGYyUFERyfZd0iemLybAryaFTwTzTgfHj38zh9CeMxEM
TOoxP/5RFk5bs4NNAMMF/RDdi53Ku5XWHNQLhlym3JTdklP+R3oh7Jqw+VJ0s1G6
dzXX5WXxhcBzEb0bRGnU8qRi2a2wkhNz8T2zJJQN2btsOyitug8u9O4NF+aEM4WY
6sLpxfsJEa+jQka2Jjo1YkR/UCWxDlLiAbr18RmAMQ7OntLbeAXlKPFP7ruaqe+L
4Yb/gwgAD8GQIV3upwogmPKJisXfqheEhNQYqWaaPkAUL03x321+0z+9Hrt92gMs
OsnW0MTsUUvP2Uui5loFZR9yZWO1bwFGsFkvkOGjk+qnWkB+/JoZu/yAamMViuFA
ErOWuhlJmqNzpdmXA3jwbIrAb5bhLYZ/ssgsT82AJc0QiSSydBlZ/X4poAD0aEip
u/O5/wBTvh2ukcAmh4EHgbMHxnPShxo0W+NE232Nm0xTbKRlfg4xbMyhCaU+wox3
50fByfq1x2g1wTcurU7+jCNenbsCky4+YHgANuX5FmqjTRMvNLp4LG4vNKk9jyd7
m9M6k6y20fRQ8FtqpFSH84NNs/RrEXwXFAOwT+jg2SG+BEW8jQbK9lLE/+LiYjud
3u5RE7uG+COZi3uwU47QOrMB4mC1o1oAvLgzUecO9z3uPlNbL3cdBkbkrmm6cle9
ebkZJRwqEqhQoKpvw1qwHOshB1S5mobYEptFvo6LAcshHg0JttN570uBkVFmxogV
qIixessLSxWSBY4JkL663cW5WHJcl1RkpB27OVa0nAAaXy6Xe3K97PAKRIoBsSwb
HN2nZN4pTEbv1TBcB7FjT/jJ6y1uimAvyY2NxFcc/suJJRx5GCvHG2D/Gqlx4oHk
Yupgl76ZSErfvcmZDY11semOtvGxFz3xp4FQ1zQgGQU2Onu6ApgrLnYv3AwMQ6jB
Q0Am+oMfzc1dY00uSt321iMw4V61KIzUpjWDubM9gZn1h+A/ir3LCKXkVAoj5ipV
hMLPOX3sNFALHIyT3/n+H1ZbcGtCJ9bpJlgdNqXUCf1n+45S9839PVvwWPO4ScA5
4cayG8twPpnzukBwPhAKG1jJTkOa+BaRb4P1ufIrBLQk8ONxBv0P1SrmlE4i5CDP
dCQxsS/eTY2sAgIzzxRRfLH/bwlQOV8vQTGPN+DbnYcvIKoHESQLj3bFKrB8NgCC
n4HBhV3vi+sVnaovA1G1G+Fcv/AC4PQWTrgbGUWNzFVUMQ2Fe5KAwtE4qS2CKKDH
2aRm3nz60niFQxmrcs+Pe94v9CBEIAU10hGyoYsbvP4F66WwnSWWog1SNWNewoIM
Z9hdHnUjwVQqCMykUTbx5GMW5B8OdYgAsNxz09kOxAfGcNyPK4nmS0FS1LzfffYb
AzdIiJRR2/NbkwwTVk9nKAKvx5gLS2FdKdmK38wuD2j5XUMe1get+6b5/BAUlNMt
0pOKRdgrDiBcnbcpnsBhlGcx3YN2ZQ9M73zh9982Ac/LvVBydeeew1/qhQCrwz/L
VvLDs1bF1ovLSVphjguRN5SxaCUsaIlauLa348mxA01FVo/SNm5DOHJ6sRufWFjl
d0AxS0hjmtG1DZR62t+KDPomLyHTcK3nmjYTc9AIBI20Etd+NMMAyTsAWxlOuqgn
HvSdJkD4MA0dCEFfNjM++3JO9wRHPQiOXrQdKu+73MY/Rcbl1p6EO+6t6amaIWUD
INfKNofj/DH8dj8pigspONFJIoW1RV6zX5kbPp4RtYp0qqVj/c5BCEzI2nvMaSlK
YhGyBkbWAG7M+hj1wrg8DQ9F7jcd/r7w4q8Xb7x0sSN3Y1ODKhfL+qReEdWurOMd
uMMlFKzprDj+ITGzP/9zXsfB+G5B3sH0D8P4km0dUTMl6+nOHvddnOdECY/sgFef
m9rWdmk1oEAYPZlLaJg2YxCtKBsVWsRoP+RX9ZX15bcSlwBrNpnYniGH367tFtF+
FCVSioTKfumvMgcgaGuJqmgtJEoGHSj6+liAHKBa/j0gIYG2S5ZnU39kc6r55mQy
ZFTFPDnrcagyWwKw6VaXS+vokWtFZ2MieO+XxeXsVALa5QJsu5OY2a7p3aGTKZX4
gvkn21MsMGTL/1PGZNU2muZ+/Icoqrhx8L2LHFH8mggfyzbMzHpCgGnP/kHkpFbc
8Dl0RiTVOxLGXnV7/qXsMadLY7VPMhRE/jV10A89n4YYdRImsrddMSCdredhwry3
4adKwNVq4nY3XBsk3pVAoeoixfF+sbhfOn2CXeqqib3jnceaoOfje+RGDqXdwbyJ
FsLz4SGEgTpG5g/N7kZEe/6ycmA05qr1oWLvu4DZHzG4JXJGkadxZhO5HpIZxd8g
SWbpM8lQUIqP70cHjzWJwQogMlGS5VvsjxqteuX3GFyf5vBn+UipjbEdmJWfWgS3
/f1jHEq0gKn7etRRPqRlVmaTo0kU1ZWvz9MaFGyvY0K8yhFZcjMtaCvQ+tY3N+cv
/DPQSYe/OZCchFROBN+lXSKCy5ncAQD5rkZWbV11LUDtKeiR04+yNkqfi6fVLPvQ
aOCexVC1WWQ5DpCRJYw386WNLZd98M1lo/TcSd0MhuGCTB43J0+SlAzv+de1KdTI
C/9LZpcy0mO2es+d5nRab2BndKmtzP7Xk7Cz8Wizi5SdXpJFQLg8ivH6JNAG9KRT
mNprq6r519a0tveDr1GdFkGb6F3/rWztafcBVi+IDUVMTiLpMtiYpYpm3OOzMnem
blmSECJarbffsD8alMh6rayn/ZgyQ7EBN+U4B/o2SFbPjc+i9+KiBypYUNDSffcc
aHZdFM5SWbEq0bTDVVKmyKe5ZMRXUYWu6W2ucdd970siwZNH7A7mSBcmTDNlhVAh
xp3uK4sm+2yQkoumNQE/3Fy5Bb2muCRuM4MVcAUzH3FNF8klheuOqHg6qC3Nh52O
e4fM6IYzYFjg8EZmpecx6Qb+w2XeEMuA1tUymhcMFJIJgfclI4LjUMVG9oG8E9Sa
v5tb3JrIOCI6f9t5uEnoEt12ywDF6WB4Xx0RiBOw5hBm6LtQnppwdPd6eiyGDNM5
q3Ol7hHgjYvx0H4vxjkuHcQ1a+yyb1shZ7jeyff53X9av0ecTU70AFR3LmAAy0j0
KeKGCu5mQTivC+LOAUmiwsUpUkF30g1MEyAIXwsrrQGr/528U4e5njyikRp2PDxs
yOPcwqZFyAKpmgRBY5J0FxBFxYfUhX5nOm5DjEJ5UvbGZbfBy7S/BgA/ZK55Be2r
lfKQXlT804AM9jz9Xc3035eLy9pI8sJSyxMx427pRZ3QcqUYEk4AsTnEJjNn8kAH
1rdHohXL/FKR+nMLfGcCgEwxBw3/7JECqI2SVGHddlSp/MjPo7Y8SSCC+oZmQNLn
JPo0CgebwV/cWW8GWEwuGgvbeidDV25gnSCESh6YeEwxQYZR0Cmrzg1MYX6F5Rr7
ukVhrK5HatVGCUAYEAPLVgrW38JaVwycjeqcJHDJIjzZAplwt0n4iPAmDopzABxF
OA1ku5kC5bf0prCzVcnwr7VJ3jaz1gLpZ+ww3D26bvRbUN9zmcYzjkQ3SY8eV21L
AmSsGsfX48YiNpbU+SAFFl25cid8GvRSZhSnuKko95iZboXn4yJ/XBeP8zopNd9c
OLMWVOrxCWfnBpedlWznQY2JHAU4+UtFB08xnZfIg3pDjelxFgwhxpBG7FYRuI72
/7nFtMJDPhQ1J22gz2pHba3hGhtBcRUfxQFzjmWP7joO+4Ci1eHhlBWZuudC/Wal
YXiKRK3+15GyZX+Zo+zSZYWOAJLvQqAeocbmYvya7GVCwvqnXnycYWLmfR+RuAjd
FRXVn60mFrLWTPszmQar+xgMFZZm3ZnCZaeG4gvdbkJbyW+uJGYVWApFX2P1ov94
exEf7pxu84FFdsHccXn+NJmn7jAojws1fInlIPPhKffqepllLVrLh1Mip5+uILBg
NOYc96RxtWeOqnQ3p6lO4IEybxupQBHBAP6ul43AbgWEurqQY7TQA4NY0ksUCAX+
6TkGAtNR9+DPVM4wDlrBUgVaNCjgDCCWHVnbxHEWMB++MhEzISARHiSZtvWhdGaA
bjNmTb+laSvbHiWJcAS1EpM/kjkjwsVEKY3xIfswF6oxjRtllwOhvIsGE06A3zxt
lBa/8VTX93J3uon0SbkXhXURgl47aD+Rltfkrd2kvDOHhDndImiJV0CjplJ/24tf
4+IGvGR2F/3sZgt2jQ9ZHQhS8sONQT1hFVkOG2uMD994Md2HXQQkBRna9D49a6AR
LC6OBSmwVg7VRUwM6NqqBXwuOCkAN/9qmRSEuLyEcZfh0CnnB/w0luqCKgW3VOZf
V6sWnfgaQOOTJNsiLq5MHx6JzohJjGAdzAkQKDR0RVbiXaJvC4z2nnEOiIghQpN8
fsIlq2vqY2dd6R4Zdkqomzj60G6N2+bGSUPZ2nPZFXRi9f32NN9X8KA2dyd35Hfm
/uB+k4Iq9R2ZsAhKjm9htttzNWPm/gK80A3CfqOCUJBdsGhDxreMQ3JURIxLn5fc
IgxfUeSM1OAleuxhPBTOsTfEBYkd7owit7QcHXRh3dSJt5BDtQGgziIokx2QHiFD
QxDPj2kG9PG/QOq3bd5kmwlt5TjXq4cilRduCnBZJ4twhQiHEc7OpjC1gbEzyXRc
aQ/5CatDHKAveiacrZ9cv+rR1b3EKF68/JuSQscwTW2IqOP4cmNJ4hN3HeoPTwwm
OW3qMVtBg0YHxMxN+LjGNtySx5A+fj0zTSUbMbY8drsc6wiCc1xJ6VxtaJKeXB8G
jJIm1dnSUCzQW96nshSz7Ms5T3xGNXkzfWSP9e+SAs5tKoAVA+Vm4ifKaIH0NkYA
1ZD5gNuvjZyF2WKGAz7SPrcNzU7WlYg7d/zW+t71KkXWbUbgyawp5Djbeb+stixD
NdQVmYb2lnfLZcUb9yGQU4Fm/lywXnPsleYWwMDGSQrtwg87wPeHc1h+9JqcQwdk
PWTIRlr78X9t33TXLSHsunos+fstFFzTkxBApTR1Crl5TakQBlVM1Dn632firyRY
Cp6dLbaJlpld87g7oR0LJnyGVzSrRUHdgz2IDIw0V5Jww5CKQNYjrM6vI6n7lZbu
eDrBOVTCJB4JGZxwQ5WjmXMngef3OI3ZdEQnvEOU41/C3ldTQj7NifkPIA1aQZ8d
UwlojBYeTRvX1ptetk+G1v+vNZD32gJXTqMuO2Zm3RGsJUFjaRuuw744z37kCUZp
jIBL6KwEiQItPxp44yptRlwNAjojj0cyHY7ysLSoUqv7y2q6AjbRblScs3hHGGZJ
fe0FO3s7SGW7gKcZ56jCByk9KLsFq7QQUv52SLB9rp5xEQfJElLcPwk1hPfLOpWs
wTB7MtSMexQvn0VoZq9H3zNIoZvxxbRRcvIPE4n9DQm6Yfymj3UjCXoSqQ8gn5s8
B13h+ibON//tTXavSR6HJpEWZwBTnSlMiS7pTkN3U2ZYnUbGPGxO/slR3LMQgTju
V0NoffthpVLSHutAl2D4Ns0iUiW8NBe9zK8Q+axeacXMWo+UqZsA5nQ6s1vvIrMz
I2dNTZ9efKLhMiqeqpeJg9AkxP53UloZlSNvsQBQPZJCazjraMQBt5bmSD72PL/d
ZOd08OO0JNKF2PLlTTbcqhIIvBhHmE43mX4FcP5+F8kEO+S6OLRKoeRTP084SPnh
nhGm3+ezcF8WbBWpp0PvKQ6IuVz2BwdKxL+OzgpiQznxfSBZ/Oy8QzJqfefwlTEl
kiNVco2oLzG4HqU1QWwOGhvWq4PXrrX69iDfAgRnJE2+xiHQHr2VU6YgC/MPtQ+w
QNGZ9HMQekKKTxXd4YSORdNbpz97JxyKHPtcC/U3t2/xPfbD8ZG1uV7HkyL3JLK8
eHheU65mNPQ9/UQZDpbFWbvk5Gg+6nP6Oh7+9DoDMkSwZq+4rHQ8cnZsH71Qlb9U
tm3CQHn85Qzlgpj1HSvYz2NkUKWUfxqzxDxH/uN8tp4tvGr+vthJU/tMdQ6Wsy5K
/EtspbESxZLX/W7DRgpnLtrOvSqV60brZSXCS1c2KAaCe9fYXMiQTYKMBcuX8Dge
FPfrzmyFv9/iepvt13yGBQFtbaE45IzPJYFpFx/QGQMPfF+9uFOuKegQS2Z7WXGi
nnA2ckaSh8ttemSX9G3vppd1uBac9xz2I8K4H8MzMn9n0G9R11dgYSF1ZdpqEid8
CYGQ2aDx0d+0940ApnceLOt56jBdbT4oEOBASLh6amkulXKFidQt+hSt+f4I5XU6
fQMAkhr1l63XDM/Z53Uh6qERt++unoJjmwTvJBUQFg28mlixQv9COyRqrnZHJ9u+
upbufe8n7E6/SD9QezADFBQBVYcAdg+7OJRbAfo/CNb9/WkPhvx+K/F2eg02dI5x
ZwuydDOZB/lsx/sotr1VXAQLVc/Cs9T0l0B+OycpunCDxNYANjqrLg7dGWsidqTv
+ytx84ir3vEEMvWyufPmcWaErjuOfeEfVDdonrKfJiPJbIip39EyHYHqD+/fC2nA
gSO4f1PHXOaSHGvD7KiZWZLMsP5bFtF4oIPLC+aPvjbhH1heWslpWHQchcClbk33
c5kENFTiTdJD/Kh7KI2w2q++C5dNezFwBB/6Tv1jVq0OGKWegdjCqnyRWcUVi3JF
XOdjWNeJScekmr3WdEtIj41UJrSk8dLrHNFYycRj0YtPHCOY6fDdhy1jaAdwRZkd
Pg5ZWr2Ygl2cJBpXt0buF96YM5InjN9YWtw69kdVE0ETHGeK9Ji7qRSUgdVoADHf
pQAdQAKZYioQnd0dcsrfijyVcmZDQfJEsCkSKZ0T6tL1b8iy3cgVyIRMO8UXHGRk
vOcB7GuHU0Cxgp+2wZzNQQSNiRsSdDwRNMGshCY4O7UJ2tjhYLqgvXjO1oesLOMk
onnSkPTVocOO04xJt1F7Ni7nVWubim4rfdjKqvU3vxqvgOtjDo8Jw7GIeOaT+YW8
QY0PA21abuYsbXohrPURcYDu44WKzpVcQMa4z4MlS6PhdfEQniWFotjVqsYdyMST
4TVahTWZT81rJ5ikDYhdNUlyxWaaxCYAKZXgPUCx8wr3wgsnPzclqBJr1hzyzCaq
gZb/qqdSZMul+KtRPciOuJKMGf50y5K0W910bPMCFHMeZEFQJE8aEgB8SacMwLjj
IHIh8Exvo2q4jnr2PkvC0QXLdi7oYUUyTKRcePpi0a51JziOSM7+d+JdLi77zJOr
dnDJQ9uL1hRFN74Uh3hbQSYfArs4xEFpeZYSPNVSkCE/0d9WNymMgK0GS0qlvZFt
G2NyYXEb4cWNopbiCFB33umvDSR18ox8lQzLn2pUfiGnWFkvMiVOMK+bT5UgAgAl
7GpoOY+OxZI1xPtN6CuyEIRPNDEQHjXTd71IgtxEzt/27m539L+6YdEaDpfgfM4d
Dg/P3sItBE4IQ4kx6l60cdUMuYMqLukyReKQQgxF+xfLbTiv/3BWogkABxc1lupF
soq1Hfg70634WyaBgKGn1W2JYCilMHx57ouf9Gw3AfSSbvK9SXPon6uBJoxEYRjE
lvVIiRDI5w7+XMxDAk59Z/m9Twok+GhbQ9+9VrH/SuIi3V6qfUxvnc3a7z3U5mwe
yDRbf2kZ3LlNJtoQTLTOCJiqdQXZ/AtHzQeQmFhoEZ5fr2HwGs6cCEd4xiypPtn2
sQC2tnpe0xHZXxpSGT+j4bP210oHWsG3r+xCYN7JAbawwSoSkm4J+86RvhtfXS7n
JvjuwqZZ2UUb0utsUWrwVVCm+Ni9Pu6CP45TV1LajYrNvWz3h8zdr16X35S42yG3
+Iwxk/WR3u1aX+gh8tHTLpmE4M/BEjAkIF3iekiGsompNPdnxab6fLzR20+pm+3b
K8SnKEewfQS+E2bwRNit5+6v3leIWXyfm/bU9e8XeYsvBYXEGmNWIy3NP6tlN8I5
NggjWA0+oVBcnkJ+sMeVBhP1xbE+nW1DPJ9nHFZ5UetqDCYd5XvoMNIUkqdPlle7
9ZsF22pGBvxajPDsygyp1v/dOUkxB6lcQjV8YpAwOKyS/c+frndw0lzdl5YSHlcx
bAAjsvJZPVJEpZlqiUgdryIREaGMRj+7bw2pnb3CIkiiAJTJCtbL76PjZGjnlAK+
PKLqctum4oUlqY88Trq30U1kH6L+0y6qEeB/roG93diRYVSgaa4lp1l23cv/F33E
bUwylITlnaOHU1FpAgQ6fCsKRFZ88FfFc3u/a2tA04LCdZAk9wHdhhGKBsd5SjSo
7ErzcX5U+74v22jBR2cZ6r/nqmJZRGBX6CN/G096i5luBx+uE72ZZtJTCS4cKiVY
JSAScexiJymW+SiCzrazznT26WdwmoyYgxeqxzc9v9DnMmJ+eYZY9Pwqz96NY2LK
RBHcbI709exXPteM2pFucbabsaHVvQ2TOackMVqjwwoEnm04lZ20VM4XVX/iiLnd
DT+QTca0s0XYU6iVzGJNmh0Sfg0x5a4F9aQyP9ngiY2WPPckmVHj+CadLIB2rfWW
tohuwukRyzT9tNCR7WacvNKg60w35s6rQxZHk719/O7G5WmJmI8A4XpX69is9gA2
HRprlFrWdrSP691uIOcORlaHBkwtLqs/q/M3IG20pale0752zDBWAmfATDAuhz1i
ddmWqdDSYA/TZXJIZX6aJi+quxDhqnv0qqD5/E6l/6DhEzqCo+vjA5v9gNxoHwoJ
22l4UFxOB8q1fCX8WiyiOwxoFYjRrkFXpCc4lpYGY2BpxQpJ9rmrPsMqtGSGuj3Y
6LbuGd/XKaZatq8FTvBd4a6IP494MpdQt1tQicMSv2+8AE36nNij9M7w7g0Q6dwq
cgoh8UFI7UlP0JItohg/6dbP+h6rwDF6n/3a8V75Cs1nsYgw9WSNJnYcRKM7TQcl
WTD0MjwZvoxF6JUI8rb4TvarFxwPbIPMUJqpsdf0mQC+2jSNBzpuj7BC0uRMUgQD
jchWTqjzTZ0N2i7JmJwrgU6GhHXdIEDJJqYprma+LLsaW8lbeR1mqBnl8Ra+PwcM
UfaunVzWBkfbUnpiBBShcpmtX7jYaaS0G9e/5lECzSMAce4j+oxfz33Q5/Rc1fF0
dgS1TLhEOCkA6uiBjo6hySLiWAipZcgCselx+cpySBAX4Ecg9rmtUBnlaz56xIVl
7pkv+FO2vApKxdeZ4NrQHnOxPDiRyNYqd36INIRr1Ht2pPOrNX/v0JZoO39or1W2
ckcTGtBtrfwMNq/597+GETF253sdbgt33ZwRTKeBHIRv4sEw5GLtefx+iwNzkwF5
Pp5t/zowGFMJrZ9rNWRDxPTs2yUcLF7wMSBGPlmHN4u7HrRZ+VeL83XV3Fa30G7Y
YxLdSBJ7Cll6sqmM48hDReE7NDXD5SbbJj4w+aV736oyF+UqU2/HAbLJUA/MNLh4
6/iM9UT7m+e/+d3kgLsDGfkPIYQ/Xl4tb2uLJhPP0U6lMKoYWWh4+zMnePT8AzFD
p0cVE2Ho6WWTK92q4K9a1ktbw5Cpru7h/NMnmwKqUswPe/cQua9GE7q6o/fGH4/0
NGPzfxmUzMrN26WqnZdG+QAiAZpjFOlPRbn5TFd0/ahnx/DUxUbZDyzCmEXidhxT
d8pZmKlvTeMW0Ke2+w4rzmHY9CWAHxZFKXRnDRzMQ2d6T9yBzdVQQNDJRSQQ5KH2
9MNLV8A6ConfOgzeAdJAd+OEjaPZ9GMyydIWmuaY1uhC4kyLCPZAWEktbYyskkom
UVJsJGjpe8BChRkya6BseTYzX71g7r1Yb7REHwVKINGJLmT0QeSfiMbZc/nK75v2
/8Ewdz9zz7b0g/kOy0noAfF+nB8ekeAIYSJiOmu7bGipiIC+C80hw3FW3J+A5Q/2
JtmMi8WJqi32VrNJ3YFU0as27ytdM+7xUOJ+N5+v+V7V142T1IWMeEEq2bxrYOxV
FoYUyslm8Lh+6PQtMXWwt0H3Ktle/l6o03RiwrW7DyPmUXzrPpUjeDfKxqQio4gs
Zzw0DsavQpzwNm7wo/AkXqJHEtlAS4KoF60u0SRCqkPNrvvSA3LvHBGMuBoPlvij
mMF6dD+mq0q+OaMs5eumvgYVkqWCix/Vqh+cRwpmge/efp+RU7QX/jGG4Af9ZIxJ
8KbmnEUvvUboUiptT9t+Z1NGtLADCRzIK6J3jzqjy1a8BWaiKVLELe42BVBwjWn+
Pzw8VGS7aVIHqJwTDeMPRJtqLzkoRHgyqolPApLWHf8ACGMLIp2c/5+PiNy6OU60
wSXJtqMPs7PtUZTi667GOva6i5fKsVONbLhV8CMF/qgxvNErfMAmEve/L6d6vAX/
jd9vKLApysf6kl7USTQJ6eG5QNfFtl8lR4JgneiEVUC+aIGfzrZ8GTpINNMYDVBE
cTU1Cqe3zDc7Ntt0B3GiMeUonPRA9kHTnaySc7o2yQvstmVTCg0iwJdD4l8BdNSn
sIN+cDsvI3zrvdJwzpwaeIgNF/hJ7mQCLc6TJSZd15QPfkUm+faX6X8YVAK9Dgm/
FbSirwL/LlC/cSa10FCud33PN/sTwYOMc0ZfheQySvYLv+NzlA40JmbWsloJS1dU
fP5oddkHAUHAxZjo/Eyx20PcRhgaybXJL7T3HQ/NuHnolAAnzrzskNb8jiSijPnq
/ccAlMlzdmqNLmwlj6PEaZOQJo+qFgTc0acV5chqg69OkAeUjEM6Lnk2EegZTP0s
oC5VuL4fNS8Qo0Wnul0fn/AWOlpyX8oWsypb66Xxqq1Q0GPXnJRpilpjqUHLKX7L
uyr37FeHjLCtqJ3HO6Mpdxr+yTfMEPUZ4kgHEY89vm3th2Gqcre05wgz5woI2GZP
mQdAi/tKh9EXNWfnkE4zMHBhuSKTST/iyBYgVvXQN+zctN6v/lwtjiu3OXJ8DrFU
0KibDeKeY1e2mC3p4ue1iXp9RyqBFsErY0KD+FBS51ERyK+XHnlul8cTnSQy+38k
cJ8SjZ2VFn75epFQh0Vlgx8y//VSqJA0KJTTcRJ8Zb8J3NngXDG8hlT6AV/6BtGy
SJar+x0dUUx96z13cfHLiIRfDA0BdJeb3oYu+Jn0Xy/DG8CJRe6SZaj1SfmxIPt3
Rv8ogxzIdTnzotoo3NKFGMMYht94Ib9XXsgCyuXSSsZI/jAKYoSeHZ+cUWJ3XkRE
QuZtAWUB8wd5cs5jdWCCIs+lGZB71lsTcxRZQaQL8T/EWo5Bs7ZU3ltgFL/TvxG/
0+bK35RSC56b4FVjDkbAAhnbb+Eun3KNhuKVsckcBFcPsu4COUpIBAw+Z6uLXxnl
z86dMmGG+S9O8OmMsDiJFiz8RiReEfN5JfbvpkAkSQdN8Z4OjsWTroAOUqs3kpfu
tQcEsgPQxJ0krhFUmwzcbGJuraBhOIDMr7Bs+F9L7PPBpk/UyaaWhXh3hWWdpwYg
L7dJVVJ6W8sKm7Ju5jjvYXvc6sK4L2hLA+23TAhQcRyYCtcLeApiPMRc5NUMVxkw
28ZAo0f02XC8Mbgply8Ha8BhIx5s9Tua7+dWT4kOXLtDXGtSjsw7BqH/cFfFE2ii
JWcZjh+/Fr/HACoGFM6iMJh9smrScFICCcENz7pPbGeETYtGTu6O43eOAUHn05lF
tslpu40PXMTM69KaqtH3JnomzBKoiAAK+vknNMlRpTkIQPcZ52oBYVN3V8S3YQq1
HpKpBcjrzbg8Y029okAhE3tU9Fg2l0pYA747NM58odta86NK28m6gDC5WQa1DW29
xRm0vwXFkb4h1A2ST9BI3DwmGVwsJ8sBoRZmZYPo488ZTsy3NGEEKtl23Me5avcl
UuYSJP8N+vlBDeq7dMddeESSDFKMj8aqPGKoTLTG9PF38hHuRtbJP1ZBcI0pP2XX
XHibPT5p8GojPGO0FEPj6elBdPxzAlwC7DwbkNkvWqJyfBlUCyXuVbyrJa0Pov5C
YrJfR1VCQS7aaqWSVS1oFG2X0kT5MMCaBv+BmtvMwH0oLXs6kcLH2swINnWk2ozr
oindRAXnvB4lw1elAcOjZZSGweEHBvPoQuOLOnhIYfzfTSuogqr7TObEb6QrHhDC
Rz4x7tcy6lPVfpesose50wmZRQhd+K9xZtb+89hHcJuhLBT7GV14dNeHZCP+fKFZ
X2dPpIASaIJPLKYia8/7himQYUxpmW9JrN5+d0jwYbboqJ61E173C91naIk4SYjj
9yUo8zYRUrBiMRsToxMkwXDY8aJYo5PUwbJY+cjFqrVIOmZg2RI4RSg2l0C36ty3
YBx4zp2X4/NMiA8y/eOH9icnnryTWFL76Rs6tohd2A+e0P6shTyiNjKTWC8k1pKv
4E1iG4yNq90OZ022v0CVp2fPACWsUmgakRRbxVrRUMGl8Ui27TjTwkuuK0cSIzlz
qj4jlVVQyTNbGAYg9EphQWwBSxdOVPqifI5eP8l2JPLclR3LHfy+5yZMCD/rOVDR
X9OjLjrzHw1RJ7cz30VKiJwcuupsRS1NrIfOW/J9z91eW9XvIA+bzj07QUkJF/xf
rHg58sO9koGWSh5qe+RWTeUnHyY4MDy06HrLZ3+uuLybhuKnwjodMCKlxGoEzRQJ
s85feaEScS8QEo8YyPd8HDI8DnF8CE4H/qhv4QYn/0ZIELK5aRPvRb30UafYNjBS
/Ty+LscY42ZHBgDWjRtc5chkiOikQQo6abHvBWupAQ2l4i586BlstiJXY8mdtAzl
Y8/GB3EoTcjc66j8w9flNWGcxOCoaDYcDVlhY12nqCHH4F50SITVZmugRVqBygdd
7iweFueAXpDL1BcoEVAH3ahOiNalC1PCi9VKrxS665BaHG509unbNr0O+y2bLvWu
9k+o1OteyKzcn3Oa+nTMFwWdEWvPhz/Qr/bXkRE/qne8vsBjW+TtplmT7bGAZiuC
WN6Rar/UteTqfyTZiz7DziXb3HAlvNcbboe0Y2+rdZudaZVhrmAR0MWnNtA05Yn2
maWp9DrIFh+4mkR0Fb+JbKYdtNW0FB83HXQle28J3Li0xhIkwBzrNi64YGxmUP1z
QSruDkwq3HHehWI/sCJfgSVTP9A93l5Ko1uUF8IiB4+LN95Hb5zxgLzjmdWLToaE
PK/c4Uq08qp60/5/qIcQMYfT6SQGzDZ1HDtMWbLdUlyJV/Ae7j0nVzDBNNDCDHOs
qx/Coz9UCPXnP62dc81l0Mvhogtnv/4sf/JXHyAd+DU5J/cPPDocftwbnJSfv1ZD
JrwVkXYN/5l2gKY2pHu+2xX3kX5ZUi84UhN24xq7kKftUYft0VHKHGJhmAgagF/E
U7LTA0cSqzUCw1Dhd/qclxwYVlP1/AeGQOtT9tucH9debNk1mmQ21YOoMDCV6MVo
2WsApa67t4uE9FS1qUUn7UIcl7VZ0cWs8IXhvwg1x3sJEKk+1wIl0qPdXTzbyHT7
nJtCu76TI+XWKRPqc2Y8nzyRn1zLx/VR3tbO+zBh5cijbsshTfn+ttzXTDC5RCMA
IipbLm/0hqQseJzGm2lxUpb1E6sHUulKS6/4vpZ7dukADY2QMEtZCFfSLul/nub2
yFz0wSv/Rt56MnIGz2Hp7Ww6bMl1ju5BWwqm5aC4FUYb8eRbvaKUXGDSW4ZkI4ds
Xn+XKkosSliYkUSs9eW1jcaWJLMlVZQfexLWrrFqpb8bsXi6pJvTFgpJLVav6gic
2nzPx35QZ9UrmvKxlhtkZOJEG6W9NGn7bhnP1+XE1Xp73N6xhCVgePhTnTWgjO9l
0o89CrLDTiCzMAoahLxzy3lTtUEklw8kOaiThWVxB6/xfvXW5sM+R1IWURVKUjfl
l5zKRzLy9EZ/pLe6alW9FO4jcEiU+8BoE50ytl9aA8l3LQnbMsNgUendrSecKYDp
lIsrxHIuNBPcEdlIBVOjfZg5gul2RHhbHaxge3akzNV3QMtfKeQRjwNrVzbo1DPE
aM3csqIO7Idui/fCMl0Wc6SvFCsRgHHoATxEc10aq2+0DtHJcp/A45yzOjhVXYHZ
TXHdc13I+JZg40NZoxuBT0YpoKgS5CQ3XxF+OP5NgjFIpdP8m/uKd/dWPZA97A2J
ukbu/DFK/mJlJplac2YDCmGFuq8KQbznDjbKwdTOClmbTb7WEk4FkMcVX/0Kx58J
Py0o9k39ZqyX/hzXeT0+q3Wa5+1oJa95WMKnLuQWlZAL6dctFvkccPVdqjJIsqjc
PMu+EP84DOGDeL48b4SNrEiJg+M0wBP7d0gTqkdLfaKdf/nSa8miLTZIJ6Ds5VXS
XhW7raSRoZIg0WcEumXxJ/BmwjWtyJBzwM8xEbe8tTwvdzQ2dgacuNy8F4Yh6UPe
hIeyheDeue6uD8PYo/kGCYPXOD53eM/3Zf3m9jYRcqJMvjU5JYiyseKOQF4Og8bh
yP9YKEgdgyMnYPZ2UfkJEwxtrUjUbCWVLCu2YKPZ31Gud6nrRwOUEjaneGFd2P/O
7x70gu9EQ6y0AwaDyBpRj5fzZ0EdQiBrfth0vsOOrOSXyY8M5XX8rn7xUx0Tf9aA
3Snmp7Q8Zy4bOMl1fWppny7oGitZZgbjY6fFULg4ln1lpHC5aUZNsN4Y9JPIy4Oc
4gGrpmEpPQ7RjVGeF5P6xi+XPRcaIQuNECaCPpE7snJaj6s4dE4bXA3EFzqwG+Bx
I0VBj85sPVtq6d2sjLWCQbbm1A44Bjhf+wgRkeqkzvPxCViBzIghoCvlprxMFmC5
wPbiO0uYVSAOjKqLUuhRL6uHuczPjafh7s9D7/0EB+FqR1pE0Rgz2ukE0aieKhZz
+5HUgMWLB7yZ0xBRlG6A8SdKeufyGe4h39ylxroBn1YmgtM2RHS/KjyC8cK5V1Ku
fnkL7vRcIR5O6WPuyeFl0hML2AA4Tt6IvWJ2uv3HSGicqL6HGy9gGhOJjvTO7dJE
kx8TKRkMA6ly2zIMS4jE0TuqVyDYyj1qu/J17m8puoD0/ZceV/SnvxacGPRZJDHr
QfBfVXvdvNzZgp8Ddiqm79JBCx08VxSXaSP46Ei6ScvsuJfEz1mB6WezGYX1jFF6
Ymf2GcEbUhZJyDV22rr5hU7iurqO1Czg2N0iahEz0+aqWiNaPjYc/vb3EPg/MONX
V5OWo/ykU5kPMf2lbeqJYrRahEObZN5+dGf9EhLSX/52l79E12VO7mTh2uAw3iG8
oyH06VKwTvGcKtCPRJyTStt7vZ4alpBRgYhocjQI5zZe+hPaTcCWFfH9LlzPVpnT
v3GJ516SSaOihbRjEjqaY7O8oz005LeR4cVv0dgpbfUeW529+IcZQKDOSoOGXu4/
0gZv4jYrbrUhGvYGKd8H6XVShkC0Nh3XPI9w2hcRf8DpjMAXdX0lzUddT/qvkqqm
6snsJ+o4o1j+JAyIgq34I6SlgqcRGVLYeXwlw0mDpp8/+lmm7DBnypPPzw1dhdC5
JuCmS5dJkfpFr5zhQ79YvcbZPQfuBiW6CuUWpwUSHqMUVuumVs6FV1AbfrxiuAtT
eGoX1ldzE1K3PguKdp66gSPKEbcMXM+i5lu7mztcIj2Gr3P7/5Aad4orJqpRwTMR
lB5kVCpeen/qJ+gulMdVZLAqw7thlF7VxqbYAQYL8vsMD6r3jHawON2X7oRdYdFa
dTVffggPpa1Q3StPbwAiEdgD1Fww5bndIayEgdwbbX1seV7mdKnSXYS1YQKmgNYs
0IYi5pudXJXbqOxxbYI2s1dNyfcS0UsOynLEx/K93oGpzNSytoiaNv3oE1/1PURy
P77h3Xrc84xOyNUjEYp2Faome9zQQu33ILBVOQr60aT3C62kCp3z23A65PWXMuTi
Qqtbb2chjN38/dZw2XbsAxvcOA41cuV0LK+uacK7KJtgk9+nJB7KHju9Rw4ZaTTI
k/oj5JvRXU4lfpM7wulSNwKKje9e+5iHRnfEADKmkaC+Vh+ikn03JrieyT9FhcH9
On+lrB/FjtZE2uAj9q3/Xtr8hx0VmN+cRVOzR+MmIldZ+PZdHNtP+8yL1qnotOpd
R/JUaivYaxvPdVxm4gxRamEv48JpROhan/PMWnztK1pwDJ6GoyAhbWuQlujvV6Se
DBDbgF6mqW0XYyPcJ38ksfvC9Gk4OQVHE45JXNRwseTwg2Sr9FhTw2prxAgRERrV
5iz3RSWcdWsDbBy91um3Xh11RZ8Ak07ElcN/uDz/gCinQrcRhhNCfW7JDTsPuyhU
cDLwnBTT8rtuorbx/jkSVQ0pzZZa1HoKcms2ZnMuVoa0v9m0cPBNJNoGXJN14Tad
i4qHwvc6c2rqdXk2WEm/iZ3ywA0/mpREyed39Vsux7Cs7KSubcqNfucePdifkTut
UAvxeU6gbky6CCZNwWwxkZQ/PJDYNkx1J3AhW3roju+ns6FemS1Z0B5uEZMo5h5T
Ih/rA9OrEgvahr9Y7lt3MtRFmQfz8Apf+Wj2RwQqMjprSvO+HSerRfxSpvDiyyeM
PHHDBYhhfe8mwpvUHi2B5FqD76b660qL8NMvOkhafe/Xi9nmX/Sqgh4RGgl7TYr+
ajylGO8/DI2t6QPYw5airiU6u9YpILEYNLqBrjFBhcZbXFamzgJsJ4TlBH7QM2uF
s3hbFM968EtIrRFnNuPutuX1Y2iOpQHpdUDsLg8sn06XFhZbqiDWuzOp1YyYhh5Y
h7ZKgZ7C6ZqsM7q+7rtR/Kvu+LPZX+QasI00jp/R9j9ise9RYUTHKrScBJHnKAT1
uj9lNsN5ezoSuD0WnH7Jg61jTrYetosXJ3zBZ4KtuGzE8aoHaL3RCwYgnwQoa9iL
CTuMj7QBL2iVa7fEPuXdCKRpLlJnRzaneiu/6yIIsUWuMXcNbYm5a+WKRZuOOS0p
PvdZh5+Yz1p9kBXeNj/MJNnc6E0InDIkJajXRbhnxONg+aHSBNXRE013eYKOXlYC
RZYqNFnR8eH8T9sm2E3YoAkHkRsXAKlFhU7AXHQ8IS3i0SCHx7trSgPrQtdRQ0M0
rkVSeG4608+e1XlOqT20FXdG+r/QIDujjCO6NaY2HzrodI7rV7fQIUGoj6OJliON
pGDO8/YJsjQO3QTRUyUme1Xuy/hPHyGUurVDFU4SM1cIxlJekhgPsMS2TgLbMcc4
cGpqeLGEPiKM+X+Zbbff8kBsys+lwUwM6vL8PQZc9I8szj68HZwb34HpNBATtukS
iNTt8AICKoNLwsaMOgN3uKJJCnSut5gG9YnAO0P4J/CTjDo/fhZw4O1YABtfEqXD
1O3rNURhDKBsWnyZgh2R6/XIqYT4YaBzYWUhFMe4jwwoP82eP2lF9KrhTb4OwKMm
mmm6t0DMntOuBU2hLWnI3E0yU0O+x0B+jeCH6G0An8TKfmHNzGnwTLeXwcJFTZ0u
QFfwY8yE2u/gERInJJgHaQB2tiar5E8txEqWq1aBzjl2IbO+AOpf5PYZFp3coC7y
lGZiwSNtgxZWzKpoZP8TrJLNdH6KDR3En7CNLuSLNu0Cl6XGFLraNWIJxCnGNDeB
2naBnV3/aSYAtp/mNbM8zHrXh+oN/9l6MBk5adm4yyN7/zP6eAPSXR9UqeW3seLA
WgZWbq8ODdV4+8C6suhQvRRif1eBmMGGnhF85ydXlO36RBOPUlZGbeG4LlPa1vo3
tgEM0SjWyDPBNq6AJHc6m3HyWuhNByL8tIXS6o6jGx3C269ORPQQ6SUhewnMYUAR
fQd1J17lLWrX0fowmcJNobHNnBpn8xDOzTGNYFYUUTb4FJHvrbJTONGfTAyonfiw
ZgOEjRnO6PpB0RHa8pABo9jUH5SFNtMR/7kADlLO5XBK+SoPvBknnsbMEf2siO+H
IFRNuV+9/Kgm5/XFFENF4qNOI4n5U0Jz0rBI0jd7oRaLWEJOEPQcsqPS79dF+wZ0
HN+z0tJtANyAtATh56+f8jwAsyWImAlgjsSp6OiFysiTfB1FJps79FoMqZn8htCw
JZtV+bEA4LPZnxrIIa089thf2AFhShqEbqnAdyrmyG6XJS05yWOgc18HBZdvytSS
ZAE3+KkAUlgqH2rKJBek43lvnwpd129hmd4Cbb7JR/qi9vBu7WQ+/5Xaqsdd7ys/
mWOTmVOTaQAXwB/PSdYGAtcKQX6xiOcFEaGDkRuKCEcbSxfWEPAP9GvarS3j/5eB
w0yqEa2rl8w+B4Tq/u6WsCqUzmb+76URyECX9B/KhCPofvrMdDFx0mBmgMy8eTl5
34xP9g/zP216PiWgmGn+PnwVhSc4VOP7uhATp9OTZiWF6Cuca6qSd5QMttS8rPZl
YWMD9zjW5qwIIZbxV8FORigqVtQD0UvGDQZtmuwOWtBnGvLWvvG/PZIBr63esFjD
g2cImM+IA5B8vSGdCtq2qacYM6nJKm+U5XrE7edgbZHfv93fQAi2WOSsB0pY03bT
8J4QT9Ks/LrCOS1dOh5HpKUeUKCQrthb1q4tsP3ki8SopyLu10EsTRNKof9ASWPX
Z69RRigBHPZOQkL1gfVN5GmUQq8KfIRZL+p9JH5jIS247dDFF0qgHV1rHNEzKje3
feGnDc7fLOcWSYyCHJEexqqaqyGZ+t3l8SUJ4x3SZvvo/UZJHU2LpCTN6TqlBJ4O
257Vtpgl8OS1YGZNWqwl08v61bzlqXSBQT6s6Ch7VkXE6d7T+zbxooFswB64QSxk
EktzpWW8IAV6fvLDaArHyIRNjHnT5F+za7bor3Np3blC+022KtI/p1RsZmhY0M3B
g96hcBew8WMIZ1UnyydsSWPw4tPYFrEysbpW+nwvE3kc5IQbHV99mBg2QdvtGJjC
eEmqokb4BgfD/jBznnwa66Aa+w+EEe7upmnEQU+IUr950uFsKXE97YORMG7YliP7
z5vW+yLM19++m87fOj/ABlIskcS0ekTLlfnuxVtA9XegIgbJnsnJdDizPJHBEQ0S
6zBHl0VY0xjHiG3w30JZTOO3wtgvchkaTTdE2yIxI0Y1yXadqmSk6+vyq+64YWqY
uJ1FkVkOWrLL1xmt6c/oP5r9F95X/3N5ySUJ2T0JX0ryl3D1oRA5PPeoSutksw9n
u52Z2Ff5+pSfV/Z/2R4YaQm+KpFX4caqKnjymLwV0UNSwc3tkIZNbGoOhHRHnFIh
Wr/HY+X5p7oMT1/ZJ2JKfuVNjokUIZwK/jZFQBsu8yPcp38Ra+yVQL7gPcwMP/Q7
3eHF2pCDIxBU2FAxTMZznUYNa2xz1lPjmuLl9WsrfMruwWQJK4H8t9rfXKlacqhi
tQiL0FskHhZtBns8VM6ZBNa4VSW0fg3uS7hZ4Od0icG+nY2PdfEO5k9Vl9pmvNRT
J7A6X1P4FSr2cImfdOpDvFIdmF8clyLf5rrxh+wj48dBkfC7ppgVK1W1L+crDdxR
CNF8yibi0LUXGzFbLAxKwhZBhkXgfP/j9/vefzq9dVY29GdVpkxkjV6kUxZBvVV5
4Bq8ia3zd0fAywzIIizQfFJJWgDey2c184SRNh5HzVBGOBl+n5OOXr1SEl0faq1h
H1m0tq68iMP0X/XHSr3ALcx2m+2ftWAPRNJ9sCEhTHQUnPbdxWBXfh8xkMWqaocD
3MkcGuzQ2PDGiTNyQ9SXFjqL8ETxdfcZlW7H7imJNkbZhnBggw68/0bS/LnQugxz
bXE53rgUWjNZ6Ceuxj00EO/l5FzzVUQ+QGaD31sgJC8pF2/wY8MfNnGOBQqKfXvY
LZXG+GFdggbQGByHlxVUbikxKDaI+R9HO2suan9+MwOu16o6MDhK13TExATcCcjP
06PZ4dgf6KQpruHRncH93ul5hu8FlJn9bHbZF4ifzbqPS3vNEteWF+KCemI+dLt3
6uXPL6LXOcnNsBrPhg0DtIfVbd5QUF/NM0SBWfnMvWCIH378AB1dM0X/YI+ihDE7
vXF9ZLiAhgBFkQeXQjV99irj4/om4X0ii9su41ZYjP+aQms7EkRbipihkELrOcIl
3MqQo38dhQGn0V61+/yIjINF5Tg952VAmqoPG3FqHz9rdtDk087gOPWe+dJDFa/s
00n4ES++ji3kF2UzU+Is93+g7jHZFXxgWobDX8aQ4AmSedRSI13Q8yWL82reuYuP
lnMG9urtWabD3CAAjuF/wqidzoF7440JwKCg1CXOC90kt0sFIloqhYyIq1Fwd7L3
AOY6UK0Cpheu6xMg0SxwDOgeF3r4EjNbdCyhSUa6o80ulV3WZnfTm731P8OBdxHJ
TSUiy0fvqawdiP8w/Q1d9FShz3UnOTV7X///1pn4eGC4jUzaaOm2Qcc8SDXI7OZ3
+f8N0DG7upWDkffbTxd9dRvg6lM1FGZ7ayzejwIMVsG4OcJyXBCXnEvHiWL9vIda
5CV3jDG4FUpgMpwcJ2LghmxRFHETHlLjJ0hQ0ddYCUkpu4S7sR00DkRbYRUijq1M
6m9B6wnuOW3HDjrpOtuVmTMCh5tvX4KTo82PBFbf/+3TdfIFTyQ/dmU/1uxTYZAS
Bv7hss48YDIjoRxzFSFdWLQvcNfMA4bH8z4w1H1pNjWXKCw/JztI/oHuNMU1dveV
5tayb/glBomvHfseCIf+KXmM+TtD4X+YXkdiuvXxKcT6mG7u3aFiWujbsQFEzZan
MfB+TsVHu/aO9J0HvswrdvSXPR3Up7PCASpgbjrV/0qNJW81ipxz3hehZ00EOMCS
Mft5TGqhiJ1plwaXinaCULOEjxp2A4qOQf+Ml3DIc1udKjUKraVDtd5d0cNGVTTl
AldY0uFvAFaVLbuDrsINMhheRTf/W6sOBaFwIDsKsFSMzDVkCpHBTOHfdxRo94c3
BEAyX6NQ1wWSrp2FONvuUAUXCFHd6/JiLfv/UTnezoMFNrUsrv5F/iI/hmO3ke7Y
3ztoRWRUcCL8CmnxVz/97gWjwK6nxqYm4+/ricz4w6seO2Twf5LFQlXlA7Q6Z9ah
YazwJkUlPDMoikd8+N7/T0y6Qj9CulNT4cvcW2w6qO0ZMkiusbuuSmEEyPwn6EDb
OSIxO4jQcNxLOhlbtCv/2siylzxVp3dilb3oceFBzrqLtJQ4K+NSaXdlO3LCX4YS
ClW8lY+HqIFxlTc38nbLo7khYxUTEcW8g33irN4eZzn8QC57xh9FMj5M/nuZnhPU
DK/L9j5UBD01Fg/gIrS+cP3Z8A8kfZR5PyPkLHMtESmMWAKc9omR4a/arbZfkQze
0yMVP5s9dirkeWQEJzhYhKmaxq5iz1Kv43bG//5NyI2prZZcet8FR39dnxOXLxp2
HIAagfhF/8Uh7gli0Duw0ee8h95wo+3yYthSgg0GOE7aHC4TwWQLpnBpGynTw/Z6
mEGcD4BVCa5OB0kRfOKyd+Cv4ElVrkCi5isp/u3EXNUPCVTN6N1gEcwtZl+SMyEl
laxmlQ8JGNgFO0hCO4FpHNGkMCO7SlVEZ9/tper363/pW2P3HR+QyaBRFKWfqcxK
9sKZ6vHaxilK6D5Gyep2aYEvfjbKex5S70o5UVvQHyeU9Y3IuMlZ2Ti9zxHL6yBW
KxEie/4xfr8mySlJ2wCtiak4OIYPY2swgbUesZC4oLHriMUtb0K8B9+DXF0li4H3
69TgV85NyyicCuY62qfzxo42QohBBlVMM1Hrl5odwvHdLfcMXVi8LOwfs62Dc2Si
jYhqDm9xdy5+mzRJzr9B42vlsVRzSnsszX5sDSi2+TDdqhC5gTRWLRK9Yc/Isq40
LZJSUcgQOBxXyL20nL73JPnKpjcQ9+wdHov/FctpFcVch3Fn3sMWsOeKzokJ6QX1
jxY0NjBmmYhWSb4f6v/h1QwfK7O2JYf1J/VQBnPL3DIC0a1zLHlS2C0BOPn0sN8o
GwtROwf/Gery012tSOoY3stL9OaVkc6Ou8Tsl7SradQYJYRnx3cXyN5y4GX+zgNz
koUlaYCePbCaw8cgDxGisffdFuNjwaVQxEPo6Npt/NNfNP57phU+uzhDUCaW7jDg
rpf124ie7GohMO5G4Yf6YVjWgc59mQhr06YnpnMUwYP2lg327zG0y1Wv1kWzDAPC
t/k/EyN3pSVN+VBOPnXQ1bpJkA2fvGj2LpbO77oVm0RasKT8SriHrHkEDJITv3GS
KwHNptaBZ7JI/Z6BE1M8HCQmhEKljO4BEFhe3Mn50xpQ03DZy+Syr8R48EuLp/Tr
cTjGbi1UVhTNYU16vnTpAgAPG6kcnZ9LJsiZUZGvdeyEz+eiGm4FSIBAS5BxSE4f
lsmD3P4kZ8Fdh1n1zNLhexxtmfpo/7jSURY9reabLL9lOhNTLU6MsVN/3nOouPrN
iafYTNZCOnflRwtWE+jHvAOqjOAGCS8MnCdUrRJjEjbegTNwFNBXsFz2RlKlFpTt
ukEcJOIhPAuWyXOt02YdQLhvyry2QMfXLpsaXCXtNQf/3v5wg4pJgeff5HKo7KBx
SQHBG2ntXEWyPIUoWayP/8UVPj87qOfiML360NF8mx10Ut/on8l/MTk273CX+KxB
g2EyQ6meyGB1ULeTLPk1pUbgRheFiCJe3nDiRj4QTzp69qjuKV5Ra7CV5CXMZ5Ab
caYOCFNJnBBLT+Pp1KFrBfSbyVp1Ul9B3BFtV9ZbGFVU1bpuGRqqR1OAGVZLlqjO
eQ0dK/iC4rVZNLuFHUZGZtz+S08iwhORQLdmhLmUGvARBdRyNM/4IIEC4ON5Qhk6
7GOwlxwjG5nYP+LennFdyGz5zrJDheOndWljdFUwFubrX7eZH5xbKXZTIIsO40Ij
yG46XsTUvrVey/zWVSW9dRZ9UauD+x76EJ0yhI5YN7bQbqL8nyb1BdNjZfyFJ9i9
uOtTrRIngYvlKtMyO0to1I0eNoZW9tejJpWA8nIdS2S7dUer8J5lMfmqO8noFDmE
1/OYI0hmeXjji3T0N0b+G05+vTmd0UYczgEks4NbP8RTA9fN92WFPOlf/k7NTdFA
ivhTYygL3HVIsA9BzbenqpmX6lMbZpJuePC2DCgLUOxZC3KXOG20nXOmZ3Rftt2o
dKLSXwS+kQXBXjaDkUA2UPmXLwihEhkXtxofZRPovaI2ggFeNaRtTfc8VP/wNz9I
roT1dkqdT2HxPDxp0c47EBBEIBlGOdYFX+0/DLePcyoqW6wqQGeFlnQ60JIVtgBy
i2pV977bREvWU5dcGmYXMx18bYULzwGVGGU7xUYmNfAndnnD33N/b/opK/IjxtFk
79qbNq9m2boiPEemlWAWrQaL7FMlgBJ81golxmm2prQoC+2gBfw9Uo5t+aPKWjA6
bFVLv47ZkYx98NDrWpQDg7s8/cwHRMPV04RsyfBdlgbM/xSduaIWzv2Upik9aWyj
KhHNI2Ybct5EaiOrT6aOwr3vWDbIbDU1GiZ3FLnoC+OqijtQ/YYaPkpLeY3IlM8r
AnuZVWfeaaeE6KNihIvh+cHiMWOBbpKboJdtvfNgacoZdgdjwargaJ/c2D/k/xGX
PdGLfpkmkj8AzMclyDswjC+QV1aWT/W8OOY7BDHjJWOT5QKxkhoyPdFQwdteFnW8
TITdd+PCn0ECwjM0RwjVJSOY6J2TeZdH0+DYDgG4mkcTmXmFGHUMIBW0mwy8HJkq
P73eC8CZkHVImfxhpeQgKhVdu/CVYewI5371ttG5NejoWpitQ9oMpbgZOfHrylFE
BftU4VH1p1cI1x8Rw2yjLvkT5wLJkfAqRTQ6lOvIcCxozsNe/eboyzUlm8jF2nOo
DFlwMDekyUy8rguKkQJVy+w8Y/lM9rIPF7f1fm83eY26yUAn3nZBuAbETVIpn1Dj
Z/sgooSUxyyZdWnIWwA5n1o/4YMR9ObMZ+tnRVAglsPc+u1qUhs0OsrVl0isEooh
I1UzA19kM/91FyrYcxU2FQmrDIaFMfAsf5TIQACT5luRS4+6jI+FEXPS++fSidrc
Sg4tlndsjFjIVZvtYmzhsuXaBYP2YEq1titOl89exqaA32CsbBDSGQOikYRwUZh4
1t4dQWTlwmmguGHA4VKgeOHnR9ldqy4jm6eHN3ypfoaotJr0tDyxk6N0HL4Zg2Fh
RW1sx850LWNmd65fUkO3Ok2+GzPhIVIBO2WFcALGp9d7vhP7aWz0dRWUAofX83my
mu6Xlji9/rm6qnJjieb8mG9Yxw/c+oSJa5N9Yw0V0/TlU6N5SGGgfBy+KfltoX+j
kdtJhyUWnaWgX/ib8Woq7d6ciJUA8bu1Arrx/B86cCcIx0Hd8XITYc+mQgT8T793
b8rK5C5BSNgn4TZvaA47rxjO/AGJZWcf9YNv6PGTFsHZohZ4NRpC/pMiOWdJCpbn
RhLshjLbzEd/efqEDTmwix5Vq0nopETRxOs+3Sq6dFfyhUcA6oKxyZ4Fxatj5lyW
/ObFcpTR1CcCA+pTWvlCty+yVWU4KtcXmU2JJ1DDX/Uqrng5bxl83Nj8Eesuojq8
DeAe6efj1n0tGqZ8rzpTtnPtDmCKt17pf2zXMR/LYpnh9Qu1jizQI2f4pEJpnCFu
PyaUU9BX8kU/ETQG4k1x5KahYjClh9z6Ppggf7pu5unvDMbTQ6QQ/h3TMyVoNC6t
5Geb36y/B9rNDgLUtCkmnqQrAY0LUKjF6zybqmH170lB1bqry5SmsPAASqO9bA3I
vSS8Dgus4lOfwMRAPGrIWoHUZyIorv0Vyji/CM7aFJ03VyWK+jaKojrcaPMCKhtu
QSzz0iaO7Y9zYB+8HKAKjwT1tHo92snNc9uCU6TiXIZC1lnP4qT0GZ2KVH+wWSfM
O09n2Y9MtGk5P0uT5c/ewKdmnSdLu3gyUj6OgCzGdSAD62SOrE/liSEKACu787JE
XqQqPeOy0knpT8OGvFODgs2KMs1Lck/6P8zgFSXN2m+iQdf4IL1VXVVDrpRxsb8q
oSeD2i4VbRbrzEqn84trFHqMUfmXDj0CCZF1sSEzuFY95r4adm+dYautEWRMVDBa
hN7KXW4f4WvmBTyOY8TXIn8sTMD0SCofFcafDlJqqq39LsyhXWwRPkHvN1wjCSgu
3B1xzGOIed280QR3gCnJk3+K7H8ANz6hVShWo/zpix55OUUonOiiYSMYe1ojKfFJ
HtSWeW83rI/vGDlkCc4qCMYaCa+k6jBoKOHmlFDjgzqdfwvDnTVwef9YLLMOIumV
grwOdlJ/9yHXb+8UBw87Umeo4fkjjZ9aYGW1eennKaP3JMixZqDKATEkDl5TBgh8
d1k8qOMvVytnI//FCZSYdVQIapv2YiYYH+XNsE6A74XS8boLlN5Q9zR1L3Odj8Sv
G5A4iDgD0AE5NvgXBv5TtXL3XpnCPVxfroWgS3gAbEjpl7wKCT+HFx6cz7pRA7M3
0zESC7BlIeqUBtTQX6jaQQ4ogDgyizjgsAnjKrRcwqN1/YyzcIZm4GT/z8c0pQMY
rvnZnCf/3ATetpF8VFbGDHQvij5+NC3ffRL+npylzkNm5dAQ9AeRXO3wxdP0IOcL
kzG1DmNorYdUBheYsZ0rdfnQeUVTQT94CRryG4u7b3Jj+NaMP0SPVoi80Ri84x1C
57hC1cEVoBPG9G7noODdxr2Fks8Pxr4KJS2E/qqgO9V1QXu+q+XZeeU1HMu6KJDP
IIV966Msr7NGH/uXVAs3sLLqr2dGbJVMR48aeqWFzrED7SMy58hxVmhxrjeWL94w
6NvTWmKjhNvXQxYjL7du7BFBnDvYKy1vuWusFBVaZieM9YaiM+a5sfQ7uuujcuWW
Tv0veab8K6GtlzESxPIRsHpRdWlUvb04A6KcpK4Ta1Ut4LmF72FREfWIvYfn+2uY
wOZNlSxkf0Fhb0GfhPjYbjNhpMGHa934rQZnuGyw80neiXaa3VywuzAZJQ2pxyvY
CO9I6e2iXgFksJbRUeCtwSha0XR8pdb0K43gEae38wfNv5FzyDEYF0Q6jTomaFGT
rTqO5beP/CSEU6Hg/WPHkviSrARq0ZrcgoiGwNn1gBawXK6JBlL25Fn/KbwWp5b4
hQWbwCA0+mExuIEtdoYhwSbxV8vnRDxlvlphxnqIyP5bNF2SzDCowuowdmj1Fh9l
LTRe7xWZNAAPrxuoZpuXWYGTAEeU/NSbEdOnfdkI0fpk3edOAW38dmvci19HAJhx
6kfR/o9k/5SqfwztHRTb8OoR1xZoeEl0TKmpGHRrA2aCZ0O/lqhofCHOGS3odEZs
ZWpyghLUWRU0by1gP/kTpVhbVHOIC6kwiJn9gX+N24jtf8MundnMiztR+ybTBc3d
AHW+UXkLt2xQtl4shEiq3Pg2JW3n9sqbQBdjU9w8+bd8Q97IdbEQIaK4k9DRFtpc
C/ufEKIJnH1El0A9aOOIif9F3TvqQS3CGXB9h2CAsyCHl81iQjd0saGfXMfAn2u8
qF3MUiTBHeCM6+CXxTqXQpfd3zo89gx5rF2jDTF/BMfDoRbjRduvRyuE47iHRCip
HcfHbQ7hv3N5bwkO0pmzKJgIeddOQK5yi+WdfxE4hOroPWVxFjQno/AM6APkhGcr
zd4ePTQ86poRel+Yyslln0M4Tmsa46aLaJstVe6GfNfedWdZPCrCa6JcRpr/dFJH
cu4RkSu/eBHAmIGpepBilWk4GCwtMbzlFyjWIq01E7+tRfuD8WssyJ3bgo7DRbHh
Zd0ovUuI5SJ5g+yPBE9yKkP1c1G2bT1CUQkvWd2ST3qSCJHoRuwNCeji6Cr5YqwE
UycS68jGfyGdYApeUl7gRnNkMh/A5ho1CMLsQvLPWNbjM2M9xAzFotbYydfYO6At
6ZXxtxfEfEcipUo67DbbArl1HXd0nwtsoXXvJqHlAOzXdK4QIHIKCTI4z8mTQise
OXNf67xPnC4fzIf29Pifi7CYbsGUdM0Sx/qTdcfD+GFjVNxFPDutomE/lamM3cx6
2eDZj4mX0VnzjhYRQUgi4ZSQpo0g7AzJ0U0X9J9VYVkctEvdykSHRLknxo88UpYO
7uWpN2VGPjfAa61Ivn+Xf97GM4qcQ4j8NLcCnsfuLmTtn4z5q8eg0/5HcqnkNmnO
ikBG3fmc3twn5CgBRJiLxD2EogCrvVXJ/6hIT0lIGVyQ9WG31eLBPR2iNkUOW6/j
/ly0KeieyysGsgX07x0dXxVnZ753BFphm6L2i9fWgQ8wPjdwpOBtnnPSxjM+m+ku
04WByUfHHJM3KdfC3x8E6LIbS4jWst4mV9UTD8K8OI3cmJrzfE0vuA3MuceHm8t5
31ZjyUfDMj0DiEgQiavmA2R95q1K/mG7CV2g3AguUaGfVk4k//gtTf/tOpyaxjJT
86sRmIUxKZXtps49+Hv4FJLm/Q1L1ZXSU7l7wd1tv/I3PeGQPMCsexUhRxuQTp4H
WEkq/oW/aikLupyye7EuoDTzFBLb5GKYHoLPB7w33dlaSs/GgGIYEUUCKm3dUcG1
8kGQWtv659gSsrchVjesvP4lNihgwaCccFOYg22mkfz8zsDDJfv758DvNAb8tp79
BxeBO1aHgh4IRSkPriIcPzS6uslg/7byrRb8MuAjh79fL+DB2s82WcV+ETiSdBoG
maqDwcKVCNWcKhyR9RHkuXPPx6UbLGdDHtaMhEjiiTFfU2Hla2y1aodaVA2jf3KW
/tMb83bZnaQK9zICH4UP9eX+bTkl09qzINdoMzx3NrJfWzfdAHnoxXblPcaPZPW9
YKOqyJ/O6poU/5nJgCzSPD7Ku4iFDsGfwUBtlKAk59ES5kYkXGfOEWupgoQ1m8Bq
UTVjysBje8OM/aFf06/kk7Gt9qgtOGPdatvFzIFWGaxtvxxvzHyWnNuAwqicD94w
KOMm0pKdl0aPigrx59/aAzE+N0w49ea0aVmnQFDOD+FFebZAafzBMXwBih35FKxD
0/T1ACO7pSJU9oSR/aKMg/4W+DJNDHxp+rvNIYgy55WFw+mcJLz1qw6BwKy4BFNh
kSAjwx5Lr0YywgY8uJS43XmNFPqsZW5emx0/EY/khnThMNtgoZt7CIFFT+PbJhPX
v1xE6c6paCMEvA5+DvlSrkEMU+EzHNUwCU4IUegq87ZrjMl7GiCHUHzV9+oqdL/R
EK4mcZMIZSJwvmjDOuSB3e9Vl5cRwSB+zRCRg/QQfUxmkTEQblPAmZ+88nqhs01u
POicptMOcZnl5ik0rCdu+BobIApIIsqNqDr6qR6WhfIA0DHdccGk4iAxXEaLqc3e
ZCWKrF/1U5h0UwyCo2gZZH0TsEt6fMi8Pmvsw2N8nGxRvFKDzBP5JGWut9TI2nQH
2FX/KiczSgzDIQCyi8Raq+M2QYOTzPI7CJohDcrNNsxZbcd+WUxZbC61EhoMvom6
89/DKortrBLdUOpLYpX4rG4quXfF6R4Pa0h42NSO1RscwwHRlHO0BpOm/NcXUuqU
MZPB5eTYJdDJrjyr/WpH7uroaHOjt1hJU7Xr1ssAuNOiZslwSn/m+7aEVeCMOJDY
Yyu47bMOZztwEJGjZ17ml+3VulZ4EnKc+oK6FGC6//3JY49aBooJJ4r8SaoplEyS
kyj4fGo4ElHgSvLjJVJR0Mtkw6z8d91jqH/dCcFZWKBzGFNsUrJ+elkRNhYED6uN
ib8lN3RGTqPgmGeVRDctlykmWkpzP0JoENtu1mg/3SbALGTm2cBhzJF/DUKrnZQj
MkEcxDVqeSNmaX6vnGMxke+mypd9+uLKvUPqBViEM/cApwdA1Fq6R9udlyZVLIt+
tEc19oP/Ia4V9cyZcBpYbpiEDJhRajhyDgpamrPpFaY63AwsW1bRa8wK51UzlDKc
eZctTrLu5HYkyNj5PQDO1VvDTV9RK6CTFGZ7Of+BlHTecR8AQtyh5VnNTx0czoxo
RWm3ta85bopsOY+rocNM0nsw7xD1Up6cYDVIm4NfTdL4NPYBCUgOHaiVra58K/R2
XKHOGAhHsg6lxFTQYOH8gRJFlc5PmtjnzKSEZMSwL6MHTlurjdpH6aX9Lf8wXpQe
XPzIHqQgLbTtMCKGNQEFPsYcbfx3YRtQ7FtriJ3kGFJ01JwsQfPsdjQzgy+CXKVf
OMYqB1SbRDt5ZGm8+wsTsFUui9rVcx+T6Qi2yX7qnE1lG4GUc4LjSQfKddU61TtF
fU//YPiATcNmRx+pPeVKEWE+0a5LVsuyKOHbO8dMjSDCzjXB+/XYArYYE67ww+Vw
J9Pv9Kt5zgK7yI96Ch5R8yzUnQGMgE4GioAfuJwW2NYLipAyjzXH+Nt1pILT1kIZ
Q5nM61e0dNFQcw/Jtmyc/zxszVfyatexF5iI/CO4+sfhFcyiZMGQssChxIkvKGUg
TDrCLxun/G0fPCilNHwM8uZfYdcvH4DSgFoSZ9DMPrmc0vw/5t/Y1J4iFm9opSSW
c2f7i06GOQAeCeAmqPWVyMN/fzms3kWDVJj6a/JPUXFeRxaffhjLh5boEDxX2czs
HXDVhkGIKOK6aDGk764SlfqL383btvnJz6IIzxBLjJTpXRBeHswG5cn++oSMAmJH
yXgfqvFh7V1AQe/twa8Yr/gU5LBxbKCT19dRSdbkiZwiWslLBR12QP5HoYR+wsr1
Z1TFs0TJZk2tm65GM8Vsuf+CFcyBGVFFOI5lBUhQHrGtjGdVRY4HDqWRbaeqCz/u
DiZfACByJV0lSyKhFKK3JTN1tAiBXVo8TUUjLViU6iGnpe7ufQUEejJ9onQGOunD
gocQWoUrNDOcz3oEgyvHHUFMXJ6E69ApkRwLNuQKNWaokRKbwSzZTVmPuevyL8lt
CQ2dhlYFGQ4Y63xmGLiePvPBHUxl3Dfud3lZRV+a4K89EKZUlq4XhyyGeLNQwj82
C/63y+/I2yScAotUQubzLLBwFzfCxI9funJJjwz7v6qpIwqRz7QY2jrajYWsxl1T
SZFJ7dj5ioBQyVHWShm+ac4RbsnhR6rFIwByZFPuRZ9C2x/RMS/w02ZZBxGxciPg
C9oYVvFw9saEtG9K4rykGrQLYYEOYYHCtNj2Y1UO222oGHoGThuQiq/PMOc94jnX
2llt19AuHguSF6EM6LG22vMLG5EF7bgaBzUC4soBlwmBXOlVOGTUK2i3MMmN6Pbt
LEXzXOwtBRjC2SGEAna58nLFIbFBeXSQJSYq38bO5SRu21+5jf43HbTthp79Eiol
ueP3s7tH4pErDN1Lfm0j9FC6CHvFS3OVlwQ0CZe/HkWLNFr9oRWvtqw3xc4nxCdh
wYg0yO96XSCcPq0EoQJlt/VXzheV9ck801194m2izvZzqH/DlwMMgZeg/7QyvR2T
iUN/F1uCs21i8ZOGFbmVL1YmaZkoZOSVRhWcPv7bxt0cjHGjitPnExgJAcChub05
bl6yaqZXlanawtk+YdCnXJd7xNvJ1w2pgfTb1tNxkpLEYphrq4K9STIw+RkN/u74
rwByqrrqOYdbhvrrYPfVJE8Umnxl2RKuBrmDG2yKb686xody8u6zIqo9pHvv1mRJ
ABPptQ8BF5ZC20ANc9/9PEQE0dKNdnIJfWedTQtIWwMquafUWVIqzMkYkc5ryigv
rX1rVJSRPmL1oxGEkjy6D6bXV1FgOtHCDVUYsE+XLWbPWY8FSp8+C9J8Ct8sIuZF
4G0kv698pPhToE3ZJxAKVA1VH040kX3KolApResuSgibeE6iTaBuxREHSio+lPEd
IRgmvtK93WugWny0Ev5dJ0iEfELazhOinZ++k4c+GBZXNNITexQkYWIKUIWtQwQI
0NVPx12H7Z5S9GNgpr1Q6GgC7NY+1v7UVWqM4hXUNXRRjsiUoMeJmDpGjxWAXL7w
mSyJ+pP2ZGK449IcwSKL93pBdWo++mWX7bmgOCPCmCKV0CHoL03lyUqkbfGI9UZh
KLxBmORiKh9+L/HpQYBpaOu16s+Ler0dtVLSziwyrKKdc7HW3yvemOqnkGRSKmlv
he7jAAH7V4JbQJkxgOI3LlNVFzy4rxXiCA9uzykEBKg01bhbaxGcWvt0+FTzfSgB
V3hiKBqYqq7yLViKTKv5UvU2LRh1FWqkqrM3aGnY8B7w/g8yJlWioWh0wheh2S8i
Og72ZF3DcCLxREEQ7JhwI+/hNqj9p6EnthCVrWeXYTeY+4fdxg1MUCCgYq/9xF6M
oSPqGsXG/7e0apRtTdXKy2BLKa/pGM87qlFphMHJezvOVXMl8lGTqQNRjtM3e5PY
MwaAr2aJEwyNwY7S2FvYhM3qtqRE+OsVsIQQGeCZ36MHB2pGSmXbasX9RqD2hQCi
l4rkHoI422gWNcV0N5uLFD5WJAPz2Zt+TtMm3LfamszsMwIuH7RBLavv7Pu8wfA8
a0GsTZv+EiaFkLS3jAaaBtqzOS6VanPQkONrEmoUJe0qXp4NHDbd4EYeYp2pC/ts
2KAAgBGRrOiVyjU3vdJ0/WhIZWxaTJPtIR232UC+HguOc5Xt6C4uZw30VpBp9Spr
Y3501Md2nrjHt6+CvNKA2PeYt346zVO3qPnbQMUdSCzo/0zNflg48Nvje8Plsjiv
DhbrCzCLYaHymGCAXqhxCFL/EY8x14twKx6l4FwbXFD+CB66Ka0od8z1c7c6rgZ3
haN1h1SzAdsdeQKrsRkhOPDstc9bwVbMqJ1X5a6TCtEoWDFDkqhubf6eEHFfb/Vu
ocsBrbBkZIdkSiMZbhXAAyppUPVQQo7Ma8tWAvkTSn4YS5iBn1g4GHNDm8/VL9l8
oKxd6C82YjKhk90l33coxwIty4qJ5nLvnNbH68hknsNlbs4z7gfaFv2NNz6nQC13
E35QeHxTysX0W8TwV25MH/OH+VrpGKuiUNRGUwt0vsC96LSiQdPnLvkjjbahy1f9
0xzlbWKe3TQbo9xV0cQxPH+L9v/bUMOo++eanC6RP/uz3eRJ8/xvft5W+iaHd1ye
Dc+9gzh1PQN4MSo67Q1s1JbwjbG2DmWzA2aIKS17j1PHU0csje7tAX0LQw4Xr03S
v+6DfWEAsYbii5+olcpFb8nv1sUTDWKPCGj+sbHKI6DOpcLSuEjdoTCdVXpL3B4W
EkGJ4JBIWJBvvsDIJZni4mqtgB51k5qZ2SExkIoYmNj4cMIFC8B1Q6eenbt0GrZE
oIXo64Kh5n18VHQt+lrjeyE44/OwetY/i3VhE7Cuq0GJLiZ5fkqTwsbxMZsip91v
ZcCi7xUVSq+D82WDYTjTkkmf6pb2tTcxbm6s8+MbTPV/5+owkruEA5ntJSxKhSLC
NIQ64VhQKlfxa4E/LljJn7o/k/1JdbMTZOvcs5dNmPe3P3F778Cb87yLdI2PP7qU
3+L7bzMuaEST+WYfNPuIKbedu3nulQj7JFW7M5hw8eEiDFh1vGbYWKuWNYGxVgnw
I0ProgGR9EweX/zCXY+9MjGyOyu/u17Fq9P3A2jm44TxrjNWTZT0kL9CApmGe/JC
LXETNzoZ4ivc/HecS25SYNq/83MGQ7zbUtWP6EbINmWJ+hyTblKiZrV34crIB03I
Q6MeM+kVeb1uIpl53ja3XnTRWHuAUXjhYlOt1w8fFGQMB8L4jWwlFn8VOaPnQiIN
fVLPunNr/Z0qZqL2GTwy64Leh0IBfHld1bkwS8KqCrta22j1jLt+I+qjSQUde73i
COxrcx6WLfzLSdBUyhOKzl+caBNiZ69c/LinV+oTDhgHvCS/8WN3azOV5p9JQtdm
Ona/jltuuMMU7q+5sXjgGWbwxbs4Vqu80TqoLxb9UJ1ceZrzqBPHCpYWknglTh3B
BJbh8RTZDF4NMEu8d52Gklbh+qUUMnHoS5QcEXA8jpwRx85qbUAGLixr2sE4Ilsa
X5oHunl4z74pf5mA8+72I7V/Oq/CCzC25HImwEnG75HyJcRRcGkxayvCvzrzK/S9
Nk0RnGMpaqv9zJDBo+QGNk/bCmfKlW/BY7FbDZXOVYSgthePHPviO4oucXHVTcbQ
En1DfQGUOMGUmKTw/fAtaLs59glBgq86DPqwr2bwsoZvNkml6MhrFq/UJWo4tOOT
Co+DMVShtter+cgQdMJVKslIG41UPGp7EjrPhTbuHgS+6RebsOuutpgXRLN36xTX
VC9LeR07HjM6GA/pFwZy908QOnDX/IkKDD++hWKjDmotJ+4f9VNJHGOuaRDWysY7
IgRKjlt70xw/o1RuoubAH66SrK5FLnpFyZnmbvvDbYpz2A10S7v26H995X2EJ4hb
rGD9MpqN3D7u1ocjJJHmGlLNC2lXiXoYdjfZyA3QUYDk7bE1Ew2d44I2gc1swBtK
loYtI3KLTWgkxbwRsVyu1aAdFRkOmJ11oLfy9KyblabB4tpQ10af35u2ijwUsmOQ
+NlUeTIfzkGtLq2lU+pjC/VB9WCCBbEiuKySYivuUq9eclH+PH1A/bV4W6zrozpV
NUEqbbeeds0TvZ/VbZI9CKJZdcOCBSUoRN1qg1lQGlaO1l+tYbOO73pvgL+p3Mcg
+Vzh+p7UcaLSD+a+wEkArjbZLb+gvM04bPHi902kRPKsaRefxOp12eyK8sNVuzLl
94NJM3JVZ6F8GVntBi3fkvkRw2FhT3DCrMjSC+dXCeKVUSARwwcti5k/kPh5J2Ni
oSM5ynoZsYtpoVdIxcv1RHKKfbXli0GrGr0rrXtaK496oApim0S6mhy297ED9s3v
lXZ09Dx/dUyQmQuD+38BBJlC/5mvbOBodi+g6nBZsXhQjxaSAzUMJL3ELcjgWoZQ
GKZHA5pQUya8UngO3mismrGJgEmSfK2eKGZv4JcC3+vX1JbvdDFSrhEoJKtTTiiv
xZbitDY5TsIf6xwF8Nov2AAxhp8Zhy8xL4m2idyaUFDqW7yH1DO18qfxGD1TC7iZ
YqGiMqErlx9s1yfqsvuLUgD8u3mgzBie83YD0g16h1mKUgwQ6+TsoBIqAiihoRVt
KM+7t4VsBfv6n9wPV9ZUf+HGD6ZS1VFhsSa7YQYpDzYpiwBaGRANqlFLuADuz5Q6
2UELMWyBwT+mM4V2yugpBffsKcPmnaqAm3uxosbpJmRuo6mz8Jyh9HLRzONdtCJw
f1631vYeGilBCTA5Kr5QptWk5TlgrHBXkLEy9hHVUszhplry6AgLfbDmp18P4/M8
4RlNWqyFREEh9osSbU5g8n3rV+I4LaRCVkG+Yy20aQk3u5FsmkHCoQKmse+iUo5o
wUK/txPJ4Jpj4VjFj8t+K/BtnH753J24EVigdLW10tPNkQuMtuxOb0xA95F8o/wO
VyceVjbmZNrHR7/ycd+DhTAh7AN4/KUMg6IJmza3tywtTRXOHx6Dw8JhDEs6db6D
L9oAxZ2IJYgcIBRLnbQUVPTwTzW/2dsgwldEtYiR8mebLMy4TOPuQJWUV9QVeVX5
4wdCofFia9YmykgvPBiDZczGHlNfvqvnKzwaQdFw9nSZJjDiKejp4+LM/Nosypag
BgA/fhTBYDcfIkzwv91+gBZMwHvdxmqtSRqQ/Mnxo6DdiKhKRakwOgofFlzhjici
X1Q/heU6To23cnUs6JcYjYVirX/3UGE/iJklKMqMeGY9lkxQ/dNOuvJ6LPZ4E4TN
ZMBSnt1HP66Oh+2faxS0c1LI2WkH0ULjYXEzbv2ZaN5HftYAksQQLcRCjmVbl0CZ
4tMmGDVygTSaeKBYhHc7TOlIlx9td4W9VRxhUH6EuenrVL4R2R21IJAncbPK17qd
Bbl3DZqYQBxkKEQvmrnNWYG/F9fJVNOUwhyTcAEaGRLyAkOqCkJAVRY29q22kSE8
U/ZRrJS8y7epW18yPMjVKwtXqti99bF9CPh2gw/sWylCr/CUHfy5hfXf/tjCnOB0
6zNCxE1MZ6SyWEU13bNpP8ocSDFbMyc7lA3c+3OnOaXJrJAT3EtCcFwg1O9qSsqB
VLxZEMKxaVW1t1GsHh7Xs4SirznMe/ndTEW7JfjWFH2X5mYgIDL8q4+IA7BFs250
KdDREJjXx7mIP8JKsTIxBj0ZHgBXoR1hQycsiLBslp6Wxzyc8JA+T6QoLo3mWS9N
eVfMc9k7bBFnOhVx0wQojh+8S1eC7PwIKWvWu7aazXs6VYHtgJxwiHuqmeife4B/
N/doF302jRQoOXxgPIEUkwABuZOjUg92F3azVYzN0sBFs9EPr7a5tU61dp7x3is/
6S8a5lmwMDJdVaqLFMn+VPai+5yk78MKg3HDvs5GGJ5GBF9AfVAd9VoeuP30VK8D
tDJdmddk2mJ15d51hByg3eRsY7KRPJ03nZKViJ1ttsTYY3GzBpFJS5KGKVM5v6qT
EebZVyGMt5p6+p1LdyvFN3+jw2P+Is5PrhltFt1xelu0ZWjd8E3NMcWNCc3uJnqc
nD+EmSPzBuSH1+XmX81UfnqzkCgdOLU63o/FTyTVwWbbEZm4PjnVEiE1A0HR3Erc
8974grpgygPPoN2Gin3zk4sxkagi3NuH/SgveJnWq5TvSyShlpYwQeGQ21agxYF2
PcvmQDPrH4K9/gxfEpY/Nx0JpAA3BzTPFkPPQUPviW6CRH/lNzszFbKR7MxiIecr
fpTLGz7tcR/i09AtcvHOppOLvZkZMqy1dC59Wz8PEgVAC3fAmdTN1SnCbcIKNNld
393gSLsLfYaEVhiyh8q8s4C+yzN9shv9hjiysTmyloPkS3lHtkvC07liYwki1fn8
ORUv4RXRtJ5RMv/YJdX/FPxrELooiuggSQTEYnbeN0DJcn8u05S3thiE9lGxcvek
WROZOD+iMyfF0T9uNM2Dva65GXtfTrT7jog2NMh3ykphmDOK3bUcZI6j+nazNwFV
9HcNh9CtJe37uFn8wUQxU3WKH9+AZ+ZbPUlgwbfI9ijgarTM/LF1VnT/ODKY9GqY
dt/7uoc24EZZMuqFMORXw3rwZkgd36xfy7jFlUmJJl8nAvdHwrh4LG9MQWXXXzlV
+wbHaFUih/nHkcA3PS8ze5GgWjwCc+0/IDhFf38f+n4Bn/YENSJXw3Pn5VKeIPnW
cuD6fFA0LDP01ClmLBnvx4e4u+NFwAuftf2Sp1sUsQGrd9miW6G+VOS1AFdpsypJ
`pragma protect end_protected
