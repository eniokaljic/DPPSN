// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SLXD2P2AtmilOfuaF+Alx5EIjXoXy+pULxl9+GV1FWgCFvnq0UrEEfBDXo5J9Anm
OpLigxjG1jcdOZT5QwMZ4fLDmMOUEAC659IVLMOHmBZTnDvanebDWMydikTvAUgF
4NW03Xim2yi/LE/oU8b5a8GPwIG1d31NuD03Jk4g1YI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12352)
+Oi3SFEZaGYCbFHT6r/mlIy9sibJTdQrQf5eFPbObEOG8v2YTJyxpwwDhkEGMtk0
RF6ds0q0X8Vc9wj4cwNSxfFGnEe/fb7hyc+65A6grHGj/Jmndw6W1UFN7BbK+4zC
hUSL5AaB90cpVOsDzFn88s+Y+WOtIhyfzTSTmYwiWV7O04OVdbr8AfQ+PRAV0R57
Myyt7c9xNUuXy8mgmOrQTX+GYCirHvJxzoz0LJH+KXvIGEEg/7aJuhAGJwjEGMoM
hzPvMAZ/Sa7ZOAqCnGv37HKEf0aVCyr7wFwzFnu8sFB8SsPwu3AItckp+Lk+n4V1
ylhDyHiMr3lUGar19eLIdHGORvv6eImhv3M3Yj7eiajY4K0oEJ9nUBIO+E1FH2p5
8W3oKUoEAr7nfC4GONq3D+yphe47BGfsMTN3m3wZf8ege2VDLnjYcXFYX1KjG6yl
cGckKkEGFQSs2mTyfF/9XJxzoUq78ZIiQIjeR/NxCMpIl3HWvCn8hEEB2FKdsaUy
YxTxaHD9s1CZIBrorRHnbeQqGcgLqlFPCpy74SnvW27eqay+/G0oRqSARCvTo8iB
41wNajWTiTLMhDKYA0Jy/FWpHp5dLcCRj9YoVItJSY7AdNiz3dDgR7483x6uQ419
85BqcLe1RC8JGEifVgQ5dfIV9kTDxzmmlB4ID1TNZVTMbo75Nx2g23gUrj6frQHk
IuNFo6hQrSgqeoSC+iESlGmuM/2UatBLsGbIcX02QYsZJkF3c0dIaIkA2ZRx35XX
+cPKlijdGnKXGWBF7iUyhSoaYiP+uSjwiqMoO3VqqwD32WNUFETBvKwW5eFguCL4
JjDlHGib5n0LyBtoQ1xljTU9DhLUBfX8523H6xn0tbbA2xCaYGcRZSbT6Uj0+WL9
UopNXYev3BmJAZXHfFhoj8tG2A4kpfZarbL+hL7jrGB7nLmyaGVPYh2epHmetEl3
NpwxycNFJjLi18zlfQfENeT5e2p8iHAlBU4o61NPLpvvqqqd6DagS5S/ZB16+Oqk
w6SXbnJH0uKK/H8pV1Jy7tEuqG+I71wCVGXIUONvx8VExis0/puwEtAduFnfn7Gb
f599O+mUHzKmKqVBWY1NdkCfMk41q/ZCenl586rq1fiZrSwnAX9sV3tsFE/aG45w
2QhkL/nbSBBzsjffoEQgB+7e2qQIAaQm6ze8ZOPQx9kSiKQyEIrlguda3ayNgEIP
mTlLp2sWcWtxx6keulhK6WJLcDfdgCOcEXnvDNz5M7f0U5htIViSsxEs21fc7ppm
UuhR7cWi3wxy8KgOMCfS30UOn8C2oApr0NxEivx7C+hbIHg/7z1EzyDSts+swDz6
apaxFi7PAjDoQXT0qdpYGRXO8RL0QB3Tg4ZDW6WRqFcUV5QWlUH4/ufXitHPViAv
8SLPsQJGwqkBtz4Wex7zQQdjR2tlZ63bW/Cfbrx/Ex+U7xnJIFhlE1zQNffAKW10
xKNBYnWvg+4ONmu1IrM5o5ZpkwFZXVcoizxDB3DHVy9sTcsPSm/nF/uyew3hGMaJ
sy7brUeR4beQ7gzfh39Q83KhxH9NkyAgcEy/00BqzrxlUVZkJoHlI/Iu78r4gOfB
CRt/fG+juxrsOwXBZDdLcnextNsH8Q/K3o6JfhTCMW+XldK+3qiw9EVTdQPgJELY
pN6MR0ADj6lyhXuIHRsrHdZDEnjzOSRL1zZih+lFmBXcaEIedcArdydWF7kao46P
uXNUURPxyfe58xRKdPizeYedd0zwVQ1SGWU3gyEVlhH1uJoe03DTvQU+o6zSH2CM
p01ow2DJgUCFapYHtpyROv8FoC2wyId+f8lQtnovylk54Pv5bJfBVPvebX3+syFL
0n+GOLTyKPTWuTNFjeymcI1F0Mfyol8gC1rmY5kRYk4lKhjNQCoNSmWt9SNZiV8u
4MwlCg7YFfhLSgiU4gttoQ4p7mRsMetBl0AO1rYsBi/lTcw4gM/zQaMlLVRgbCOu
PvN9c9RwL4tsW2Vc+MDipq1QHehoLsR00KSCzCN9Byz/mlh++if0LFmurBmrlGMT
NC0UmCuBnnDchGMd6rCgUN7N2zymCwLj+mt7gIDVgfiNNc4po/O+noKsznQbvyTU
/28yTKpM+9O8S58oi5oS0JnEy//fHmkoT3b+RTxuEsFXmaVFZwk0gSVOLyQtyetH
vNJpxeOsVX+PK0Yn51ossr8CQfsUtXMlqzkBqK7vHVfF0UErxSIHX3N7/zHZbpbY
i1I2V+E3X5fY8e30RgF0TNAeYM8+HCkABjEVFtGym1v6EpouFwY3Xl37oOnJiqhE
97uH0SfeLubnA67xHLmvGjyQ6qICygRkQTncjErRRaXXnR8jylynLb7NrX6i41IJ
pUuYdZ2YT5ZLvdD4aazZmafVzVI5q8n53D4grJzT61YKi0ZLjE2SMjRIStJvBRNJ
WtLTqpNQJzfy5EovvTUqDYreCe/kdtLBTY7piowQmGm4P0Ejy5oC/wkk/kbeP3kh
exkhifemHSV4ll7MAV4Uo6VRMvVCVCXjMZY6wZutmRjfNpSWF5xTHgcG4Oe8J6Qp
jF0Hf8XDW20ilRf3xYEUb7enX8BmDI88dIVN2JF7wcMrqy52YOBSD94ePV8SFhKR
LEsZ8ojJ9CIbG7hHWcFVd9FEZ4zWP2JCpTtx5pPWsGixilggTAlK55cLb49C5/ui
qSBHry7OMxMWaHxREBgqLCSrWviD0HgR1mdpN/DmEQ17krsK+LpCCg9YQix5LE8v
DitYX3WCe7ABU0bvprShJGH8Qy8zBleLyv19EllKfq4y6eQtAXAixJV7zFf9XynD
uW4hFUrE0Hw390Dl6e2oC+rkZlAsyTlnXkh3J6kmog7S3yRzv1ZcmxMt2cn5w8ut
3W5xOUYv0ABUBM7AHzbnaA3vnvqD60yVEtyaxB50A4FfGhoACCQvYq8zWiMPCwBc
6TSlvdhDrEEIRfoFnzz48gmSrSXDbB+mt5ZJDuqe5JZEwsaQjPWYImB9Gyd9PdeY
46CNSaKW4xijT8PSiJ1ix0EyTmrwdGxbdLKzHskqwyLmPy4W583aGk+VzQ9pOTyY
obfc6K5w48Q2wiruLA1VuSQ98N89BpmGDN5y2A0xpK8PXdNnHCfu8c8P05OIF+qN
MXoisNO84DRfWUZ+SbAPvFCQEt3F8g6cF+NablsB61RJ7aS5BwQiWFpcCr7Dlzgo
0kyoqT/3z7xcJoQ8M+StueEDhelhUseN82Vchs9IBrpdMLBrq55mmo1pnwcVMyMD
gS9XxZejX/L/aQJjlORSzwKymIzggE8TK/CvaqcaBgt5Umn38Mu5Vl7xjbiICGY7
bXlg4EfpO8ZsRV2FWzMLIsE+eru1TQaY1jS5OEYcU4MltTSYKijTWqDslwZeTEEx
jTaU5APvAPP6ywz7J1d9aDrKE9UOtG9DcOzdC/sEK6wkpp3Z6WV13puUTtVSLwQF
XFh9Qi9lTNKJ1UOhjkc+VvzOvYfem9oTEjhaIO1/MgoRi6J8adLSJRWBdvEKo9/W
sjr9B0k28paetfvTpv9+GOzzIzTElO1xGG5EC44XaqdefNmJo0BIJ1CDmIBIIhsu
/Sz1WQBFoG0A5Xpa0rbDLDoUUiRgnfOdh/pf/8s37pyI9tC2H68z8s82X+MMIdpX
NCLrMv9HDdGKbEWGfqnSsp94FmZeCSLyovMVo4zU2e++dqpSUlIgZOJViAqBPeUn
UMup3g+Q8jdfr5nHDSpMKdS3fxiRiWV981p7xn9yQan+OSkQu1Aw4tKcwKF6aK6u
O7+9CanA9oqOm0JiXCt0A3Lx2uEfhj34VLDOZ1gTqTIFSsqGLHC7qTQKxAM7uTti
9RD6nLzQ51cMHJl8fG06ztrrzD1hDfdbCqJGtZb8UVWl2VzYTg+V/CJAsqbUkd1l
FFeesh41uRm23/drikmf9xrTWw40To1WiJFvZjQmTEIRTNt3uvFfSD49PQo7J3VU
ZcUTXj/KoqxZnLkhVBeDiTJ0noVegdqkdqr75oG7lNyCf9oIWrjKTrFWmwBiBGhE
jSoFNe18412DSXlXy2lm0nh1FsSY6wYnZQgec7hcNOiwKHEnn5Woi+ux9BHyV7ny
s2DBbnNTDwHTgW6fxXAkcZDCHMTCMcN9LWnfpnRdTxa+86pFw8WAsJWkT7PXTwEi
KCfrR9BsRYjubFSeuG9bUXMXhEzDILn61E6ZdqwvTB8aXACCETSkDDqP1m3XCvJ/
gekOtz2l1IPkAg69SxE58UB6/LSedBjIu9vSEgelvRueAE87gKLEBFHQhPYSw59d
5BN0Ib2VfH9J8snuwHmeltNfKsssAX3jE1lUao25cLnrOlOW+4TQoCw1Gdc6ddC4
QfDgpzrmNBBcmyURMt+bv4G/K0o0tjjxs0jFlWgPdFhU6Dh2SflRkJECBrkf50k/
cOt+UEQt6YkF9rIA/Q7AkcIcznyrI3S2DYFH381AAfmX0zYS/uYPmKRdtdtP9ewl
jBUxlc4Jr/uNdC9JfuhtscqkiekI5ym6oj0nLVtv3GGrIw+fykWr7o0kWNHIBGQE
ua3EH/ubtjZab1p31OSe1iV2VsqT4oSh+ZUidRPakppDWui1hQrOh1dLsgW24vum
tZcEDlxbNptHzr8Kekz7kuy7ncFXggVNFcGbM6XuD5SDt9wpYrZB2MOPJSzQ/qIL
bjE7dKekYuzRLsKnkQJD0H9yp4fY0F2gMcS64Vqy47JSo+4/n5s0NcwPF9/jXM5i
WhTpGQp7cEPgdVtEwmngrUpkqwlgb4NmYUFPgMRaJq1fq567onaw2REZJGn1hSAX
wvEcHzuTnKQW2cdv6Jma8YZWx8Itc7W+Ux/nKflRXjJJFDqjYnsm1kbMjWzlKPNy
C29zXSRwJ4m+2bijQvHwly0fLjLq9Cqww+otLl7TnOY6QRun3snW8hlDTxozM3gQ
5NVq1PSoJd4U9oeOWcauJ2f6rKEPcogjL+iMYI1RVSpqaxqAtsBNYtq2vKtP15aC
386B0wLD9DKJ3by5YKstpafoKBihSKRSMwE+CyL3PxEtczb5pS0gxaIG+CMxbxEx
7SN/bsw5OPxzgQdtnHi1s6T2s0aM+Ejc4OltZqqoEcp10BrxOb9wQZXgF3u16uah
lInWsB0Y4YsM/GAg/BFxqxcRsr9IDQzj2eI9zHKpj5YYYp2OR5jqlvSlVysRwUjR
Bp+pwri1S3gE0Qrr7UJUQ3BTPT2oTJNhcYQJC1XJUQYWab5c+Osju7jysmSMS/fe
btQsL09vtke4fALy1hc12wBQV7MIQdaB8GxJovva5pDf5bpBW3Gk7Uh2xjiVi3n+
PZr4uAdFOFkzRNC22lbPiLKc3W2YsNmRpaz87SWBkrUQ1AX/FJekNeTceEZkYDzM
VqtOOxAN2KIP8nbhaN7F8N3mUm5wl5fZnOdSQkPCk9lkajTGlWLqWw5Z5JBjEnY1
bnxfADKMAyVF3ikCsU4ZtWMSPkUqMNU5GGqFradEw5WOdc3kvvnbPHDmLjB1v5o5
sqljc96tt/JkW0+PfIkYB/MInpU6NBoNIk1A0x9L4eNJOiewvh9MHMVmmcMhtA3V
ArkKi6zlG7B8aGtZ6sCMhEPHevWebhQ4+9bd/iJ1Wb8FL5ByRAStFR8FxF6/WOfu
+q88aj0nVje3HY3u7r0dUa8IWIx/fkealMhdf11z6HL4NvUHpuJGtiC+msYoU6xN
2V6VZIu667CfS1G5Zxy0DFoW9OgKDUgQHt/axOwVk8QRMQd+63201JPIahRhUhvy
nQrrQ91rFt0+uH2hm/sHgJqW34dprhh3iCq0Buh/zY+eLCljTH7BDOpQSqUVUvcK
r6RTMhMB9tNLw5S0SsMRoLDqzA9JiJ5uCSHfwReki1y4aRWxFBiS5JIN/OFuQChY
/2Ra8SaVf25hM3foVLLR71h8QP5G/n24tTOlc+w+KEkarqoZov9MHoqbJrJrcCR5
9sVQyoqeS8+egsDs7etf7q9Zx01gJfd8zU2ZSNplIc4ulcd9m5RnEYnVOr3TmOSX
cKHYo0ScB55k+QrVeJflBtnePEHzKhOU38RHoJGAlkuGJ9+EBM5f4ESlR4SDDHYi
a7nUPChvgPA1vdkJxWLyNGGdzQiRBaM+Vmhn0wLgL2Fl/n4QBDPOhVpfMq4Lil3P
V2FBm7N+eKzZ05ltD7fwr1HIvc2LFiSRm4uZz/Lo+1UojNwGjnOuY1DBuIbH5LJa
NBvTxW3YJ5yMeMhMV3HjHQMA4SdC2C2TRxCmWcZn+Z0Blpvotcjxr7nv++bubM5g
FMN/+GsGsOXwzk25rE+tFOSh2L9Z7siCDjGhiWWsRCYbrrE4KBXX7Ff3V3T4/TdK
CXdMjwjd1YLe7vDZ+SjuZK8dvNbl7NKlwvBNdkEb1jPG+9l0RSHZcIhpdMq+fOb4
5pVrIwD5FtFc6UEzPUttZtyVFJICwXNz3VAgOliHedA7yV0JMm3CI3Vy3XVQuZ86
1YPUFgVu28qN20POUeeOeYmZ1Jkbgekd+bFN5ZUdSkEw2c+AFYFhM7EF3ROPLASk
0/p99RpQD4i9fJ0uzYE1lZIgR4lJ+pmXs0PGzt0QeWnohyxyqjKfbOLUjqgwjwyd
I0DBjW1Bwi/Y6GQo19y7lYqm+sq/CJTo1pPyckAqIX10SDaNhyKxVYh7ujZixLyj
jU0TO7iOdeQgKc1rGobYJjMsTPACmHNIZYMs3bKf69jYFSEWnmNrd3vhY83iSVeT
sL8XAJgdYG20XSkh0P7uBffACrI5hktSo0vWL26io5s3XQaxZEfg5r3PIT9LcxnL
8RRDb7VdhrRGxeB0XH+opRcjV30yCJM88IYBAsLPqkiauIAnHjHIpI2u5JORp+JF
nwzjaBocsNS6E//maLxeKN1cQ7icdjvmGyi5wajCPrHFxXc3W1UgXOpTM6+d8/Ow
wsTH5kX0kLCD3WQnszDCKb4ZWBjdKoLaQU7C2pK76A25Z9Wot1En5GMtMceRQCny
HTIs4JT2TXmAb7BN3UrXtn/CCWGZaNBMvbNcOUtqjabsq3D5fcgY4tJMRnzvPQQ3
M9wy4+wkVLPm24LHdrE2nMlIgkCYahZJCJ65PIXhZ/YaNK72vFNNqEGsdNO0Lk78
7u0/vXhBxsRC4Ac1dUuLueoxjqgI92wIW4kNm1enV7Y3QJpz9YwBeCTJPorOfrQk
uw27dUpYQiUl8M9ZpmzQDcAd8EFgqgAhef+GOwm8CZlDWDb3585E3VLbtfcgF6uo
1LevCMUDuq6HJxcWoYAjMz95D8oDfrqbRxw98LqyvJvXDmOhnMri+0+Yopih20s8
TvxLkNRNjKQrWBM0jyKASagAYVdHQrgRpQC0FUmSwWVLg+EKQIgd0ENdcnU6iuMo
PyMhfdlD1JeOavLRvjhkcR6c+9+d5ObxTJJ0SM7Ps/z+2K3Jl0k/OQSCvACkPneD
ym2MxduCbSmRKYgbI76ZqDfND+DDF4Tr7EioQ2GTrY+B0P7mLcL8M/3NntKnsTE0
xNy6L236r2khqiidfAHQjSk3lFRv1aXjJKuPu9vgGf6jKGSj55ICo/MRISBF4aE3
KQM5FU7RH6/FRufiEf8mOKo4/H6h2csWGgbjO9TOcewkd5H1MxYBsRVHqh3ZMGvR
ctQuHRfTYldW/xMivGWwugA7Un+nHqaLXiQT5lDBKnncs5oSa99RS4pwvmmgPLuG
cQfVt3siW+yiJ4ZnTeiG9cL7hGP8NmiwzDBGMCws6WbO9tVjcCCc/QwsyV5ocL+t
j0asGN/uov9ErLzSSerUWD/4PfUQjUYMqE+cFVfSDW/eUaH5IeBSWoWRfpuaJ9WT
4+jfTGG93alnvWKa8pD0YuRO/sJNcLcYBxRIF8y7ezonYYWb3gMz0hr8oFnWTnjI
ViNaWsQA7smlosWTsPYiJ/oADGr49prlF/3Z1EbQqTBZFd0yo4er7A9DfckadwgZ
+H/ulqM5qpsyBVGetqzzF7Ey34QILUrkxAzwPSwcPZIfnUIJ3vFsRtmXwkSmI2lo
y9HXenvegx/ytSRZbhtVdVyDj/n4x4tBu99sGmsj0nhui2vnv3xm0E7H+zFGjmln
u7b+k5nNapIsExQrmufC/GdYaOUKF8VFcvhQlFPTHQb5T8W6RPlbE19j4XzY2uAV
gWO2Ozl+qkh5nXJyxyeGDY0zc2DYOVr6wN71aWhGQ2PCziQFTWNsWY8SehpzamtP
1jES1EDsmJVgio/6uyUWofWA0N93kof9wh0vrfVWUv9eo9LxPVpVQOBW1OAMCg8g
kBUyQ15WhVv5vGngeFFA1SnGJXzoVUHe7Q4vv5MC4eCRQfI5VjsE21Xk3aiR1iSi
Is/qdYQTJL19H/P9MiNCPi20Dib6S1SpR1UiPyXLL2yP0sF6HG4VUj0x7EG8ljv6
jWCJPabYye8mCdi71cDmNtpQYmIb4414Uai71HHZZHklXEX4fkdAAl2OyPGia4Q4
DYaxtBkCLO9QFKgelS2rpaAmQ6VcVpZwRgkakYXCupfXEfHwS9CHQ7afQVDYRC2v
tLRgdRZyAd2pIzIKePkLY91gK7hdtpy1b6YsiTa8w7uAOczS1PFnwBn4yasn6jIU
Gy/VGzzp3IiswFg+t+RkETB1mT52TScuqwGMJuirpEJM1AGDvbUv/tdAqziH+jgx
SIT+6pH3083hZQIQj4IEH4gr+5GYYUp9WuuVIFpS9TSGRozyQXNPM30zb/HXala5
PgNKtd6P9+uCJF0nAJcZJPCYh9b01iFIFnvwW6v/IMfmdwEqUclXcuRHwaP5zTWG
wUR7I4RRnDnypSCUAlGhv5pflr6aCndtsIm6wyky2zzL3+iJ20r+teVi5eRo+XOB
hSgUMfdToquF0TpztXbxVv+PCYoyvzDgZ3jxDP7pHB3xEqermXcqXmCUDisjEjx6
aIVGcy0/Cm1T5uKCW05tIZLCvUhHeyOnLDgub7Di50gqeUW8fmenAOLpq33DpwZD
FELsaojmqq4LgvTr3DifVqBP7P52LLZYw7Tz343/R19sj9Ypy4y0XPBs2odpFgV1
aA6q/B4C9tFVbwQWii6+9aJ0x/0ZHb/Rj2+7K2fZk9x9lrZpGsdeceouxq4va3ma
6WMqGf4XyQy8Uc3FLUwzclIpYFV9EYp8e64oz92Yd4eYRc6820fGBuEviq4b7Vks
ttgLmNlauL9Wc8m4p40k0+hrL3hQvEu8uNC4YBH3EJ3DH+uBVyIGOAh3Y9riFsaY
128HLXepqsPwF1n7g4on9lbulPN8A57QEO3ObncwE149oDi1hXA8f7/Ps36dXfrS
6Eq+5QpDUU9dGfHPzoGLZmE+zj8X1YAjVaUcDKvkMepRYu2DtWIK9Znrzrt6xEQ6
gms3fNlMYbAs3xD7evX53m6wz8ga1ttzW8zhIhbk3vtpsN3VnhJlfl0/YIkK2vmn
0pdHvcdtAyG8X9dM/DBhO9QeEfIdi7BVbI7Pr+CBBuMNP2s+RCgFt7zP9kdtSY5q
JUzbdL0a0gkuhIkk3TZQYCTtQ/BzXIgxcKc1lnZI8TgJl8Z+pIiOA+u8hjQS2yCL
baeWxYAmLJJ2VPHQ06wN1UYsDT+LoaNI2UpPult6f4rbbnnLlbD0DUptxbjpW1g1
9EksLBNeGiRD4bZAwJfXhpuKvFmT2ih9MRvnlWEjKXfICzk2jz9g6BT6JReLT8wQ
2PWBLGwdwDHUbVIhZ+PDfyQErNOvFIgQe41cU7RsOk76/IgarLQjDzVl8oUMeGiu
27sIgz6KI2w0Hljtx22oCL5dDPBu06EtT3aCi0/6GI9PpFsMrCTw2zmtKkAK6Gp6
ojFX8oh5NgJpLxBHfxYMkp78zOtaoZQyfh9SP6GCyVsPkzlrJPWQ1LcgXtBgYWtu
2lwtbH+STfr/9u6yNN75wZ3xQmtAIcUPCjjg9yyImivd4btx9JjjyzwhokCjnLDC
wa3vcPd1coI5opQTdWErn/n4TfCPf5SXJULPhmKr9ynM4FO9ZJwDgtpSlZeu9GAh
Bw/RvCWWHhmPn4Fh+ct+0vA7p3V7L6lTmFvi+wKg1hHZjlNIIgN7n3rgDNm7AD5J
tLn66s4hT0D5ItFkP0wJHFXNWWTH9ntVcVh/y730lnQktcL3YzOlNZdffw/3CFIQ
DBilLc9Kj8mr2KZX/O8qEKGkqtDkHvg4Fwq7NLDEUQ/U5BkAyhRLh3x+6mJaFSnQ
hnftPkPGVu2tYke7841inQCJrsb8u5tToyeF2Sp92t3fSa7vbPNDLpr0l6qcNuxF
tCpMterRYyI8tIHp7HU5JbEQPbUfwFUCXbt5bvEKDKAfJgoqwnifbk3YJLbX6Czd
XTBhXg9hFEpbch2ZhV23v2LMW5lv473jdGrfpFSvzLj8rZqNa0AkoirnTzn/DhHb
wgogKue9lRf5yJpBl5bN3a5VS40EiDQgUk5vVfju3qPvDDUoaYaYL1Mb20ho/Gdb
+J1W7Rk+7PUaVMgra/2ClpQKMGp8BEID1UIg7C1lWDMEwusFwpfnPYlODWrnDJd0
CmMo9yZjAoAkk6nTKrgS7aOIHbaG1yjmmBFMDmekAnWuJncb4lenEkvXVkbUEv57
bkXJvdTmCm/4ncDZo1LR8OZijSXBkVv+HI3gz0iEsEC0PvE7bbivCYaosNE4BmY8
Ywe8Shjbs5ZvjMCssSieWyoVa9OCu+Q8FKqG0v/8VFj43MU1hwc0qEtXDozLJDj/
fIpTKnvXq+yMzSPZSara4nZXhqFh8AxOuBHwKBn0b/TsDfvNyBwSZYx2IOXCdBVq
wD6zXIkxVyNSU1ZrDtSdjkHTOGgPyUfYg57iOBYtB+OELWv70wKUjIhnvHMkTrS2
rnboeeBrL8embnPsiUd68cbD94ZygvfGX212iYxgRiPrpq298BqhSpbO8mZTG4Sn
6LiJiZCSZI9ldzWuRDmrhE1H9svsWrc03oyOpDVhRgH5qMcTfLrC2Z5bwiSSniOc
6yzY/deooU11HxfW54w0B647kBeMZffPEPv2zXCFydZBoT508QNffjiQlJJxRTch
vXmkiKPObhkLr+p03BuL+RzEgF+qq+m6C1ndCAF/LHrykDwdkU7PGL7zjWFyMr7L
aX/DeSrI7XUC1IO27mUUWwmkHo8GYNkQQhYF3vGAIHi5MverJi5HCkvk7NsrDmGy
4H+AGLxYvcHh5caL7vl7Twjfmbp423XGVLyioV1/IH24HFE7g643Rgx9aVYrfL5Y
iA+v8CxpIQ2BFeIwTWWrcTJ3NCxM5JGKnHHthTflu7NUZt1saOFpLxJxzYg+SYoV
zub8i224WGqbzYJezDVQ0UXF9JfM2lCDWztAgcPMP/Q8B56wVKO8gpR+GZMbLjQR
oudn4e4hn69VgQtdX0q+zJCcqGfAJLwQTf+7GwucRom7rHyWmt7Z/heo4kRW+fqp
yZfMcpd7CHsgKj1ddVI1YqoNA2C7eot4RgmGXRgVSKbxm1LVCeuT8wgqmIf7/irQ
7wG4FgIS5N0Y+e5LLNll2ydBBXpDJAHiDElCAJzGjY2tO5z56joMPcz2eYruwoO5
j6xaShkF/Rd1Z/VM7uqhOh+45buQ9nbhvQqzjtuDm/azRzchdfRwLsct8c1z692r
aawoBItzPVR82x5FV+LBi9FKlMKonLLS11dJ2vhzWuVO+fmAihvQFYsAL8dKYcJK
FKSUAvBi6m4BI5E4Ok44H82nJg+6in8suMcgAOQKkl3UNJuJ0FCZ8yLN/q5ctgKM
4t05SCR4lymMXrOwKfLH8fF6UvlXJl0zWsk+8rbF+Ku3H1bE1oJVcbEdu1TIShcs
GUBZ0hV0P7NOnICLBtkMnptMcTCat7UCW6Q8jo0K133DPLuODn+S9kXlX1wckVPH
tDMAG9Mxip3ZmnvPHdA3gL0f07f7Gi/dTwpU4JKO7wgom8q3t5OQUqkwpYRUU7gd
BPsX3ILkWY5aKMTErKguxo4TlhbtLn7bY53InE/2Ju11tuEKNaOxSBbW4rli5QZO
Czhj8U43Mf9hSwa0a9H0OAmtHlmy7A7LkBrJsYX1LYP5urta9FKu+xWisRWotVs0
OZBfzQEJAIKJnlVj0mrkEmqCa0VZji19sOFg1hwqGyn97BflmSSfPerveaX+wwuy
4GRvqJyYJCiIbFztLrDtuVowiGyFAFMgTK2cP4TRxAbXGfSU0Ea63RHyJl8DygTJ
YQKkm7g6X+9lhUo1EbzU/eOW6QaTEfwnXMU9AlD3JahF8DSJ4jzMl1Q4PpSo9jaP
2aq1yZMK8+59H02tjjWXyBmYgzZOAUm1yIQLnl2MtAQ6LLqqxdPEE+qZkmo50Nn3
3fNzA68rtomCoDxLcq9dxPlmOjy8gyyHuuylel6u3r5AVvYQ6oaSb2QWmsGzoEd8
t8pLQzIlN+i7r1sl4CMdA1qms3rI/CMHdscK4hU50x+/Fg11uiv6HoFzG3EHJ2kW
infob2zapVo07sMA/q5T1PBxGUtYcyehnPlGZccEfl87i8lHroP39ibr5K4WtSGX
sFD5cc32/J/ahJZDljLioE2m1Lpi8OEYdkBkwuqDYCKurEZW7hndjbdjro6x8y53
jtcUvk3TFeit8UsiJKtJ3LYMjtFq8p8OomGkVctid87V45u0HvxAe0Qt355U1LJB
ET8CCdB6OxHxcYOvPQFnkt0KHXwVxn4rDFyXf5DY/3lMhdR2SgNabzk8aGz2v+/c
51ahnfrttzL5byIJcyu6oZEab7KKNLuTJOa76WAHJ/G8M/qoNrZ5U6WmH37NfcAL
dLIHmr6Y9ZpiO8YuK/jJeyAHiM+E8gDX2I5A87jwPwNLXtWAbvbP8wRhAFlNE9zR
QVA0ybYpAeNNw00tkGRv4OWNNFcEVlWta3KnTaI4rqb5w98xlPH+6ym8VRqGzjh7
zbvs+SwYxjgNKJwF/Aqed167TjdDUU2HJC+lxTwOrJMb1BQUyvvBYRkE4BT9hwCf
uPQjWOttSQ4nWYxWXbWDQXPOXzVX51COdScFaUCBLB/8SfFHLFPrCKskxGa8otaZ
TZld0wrN+fw/2hNCABQRRHqG86P2Uq8+vjaxYdPGGL2JYgRDc1tatPQfBv3vgRo1
jB4u7bBMxpwuHmeU0Z9Z438ivMgCMEqknJbYCjyqR7b0RARyJ8iUqYeGr3Pn6SR+
i3Mpos6EYS90aVLtyWVeorkl4LKdvREcwylcpaVSe5433INacudp1QeDXIMBoEtu
VKtl6x/Wenj259bAkvq670F3tv3AfNnLo0/VNlOc5slEZZmzp/a9Xo9xSCRA6wgc
iUQV7vmIwKmmgWAwXdQI4nx//rzNHMl1cTU2fHdAtE/QPNUMBcbU/ek3P1W9OB5r
aseUynYmR7tGt+1sPvS/VuAZrE2+2u3kACiTgsnGxIHkYlTWJO2vekrAP0sfwG8x
shgsKmyE32RjBSjuJj0CNiqpE+mCjSJ7qk3hgmzfokjNM/i01FOCW7vkpS1sPfxv
fGjvRDy57JLgrYXSLUACJ0yKycy2Z6B1/OV29gtLNOpx31xYZ6QqnFhcIk2LeD7N
WzO1lFtji7l2Y0P1kN7vDc1MU5JTLfmvvzWSq0PpfFADWN+9hFbSoho+BtVuQXiy
Ac2L3beOgYpfGcKPYAWIhMpXn513nM1WLd6sjJhuu/FZiHpF6VqTQrQtSktpVjhT
JVAFrAxU/vb13zyglyoT+6c4r+H1LCkNS5nEQV6jZjyfxQDA/uc+5OGNLyC/uhLQ
8c4jyN4ggR7KAXYdi5fXw/YIRk2miUYZ+E+QoT9pVkTIWOSw1PKoUWcLD5+oQ5fK
gr2g/O06rwzu9sFeJW14cqgeCYCMu0KmuTCskiz7aFPaZDcpjgQjKWlxkAgr/YYD
n/fwtgBZBnRznCzGJcku+U+l6iMVtsNsK29Uwa4I++N2P737IHs266FJK02Xg2Zz
1op8uGeGbBrhi8pNjL4gYP0EsSB5rdZjB4YAQWy88detTbH+T0AqailFemkwAj0x
RDfaJqM7zUmvJS1htCyjaZq/IH4aH3xYhJht6FbGfQ1nXeXbRvsc6YII7LsVwqcr
UfS/lZPJ1OdYSZUY4TCPb+bakms5BYOT6lPklGg84oIPOx5PPk3ahrliClRZUzio
9nMf32WUXfiY8bd17pCqrQ2L6Y/kyrOHS5Z1bSfvLm71AyaRY6epLDGQzI6bqsSG
4tNOMhuqnLkyfVTW8uzNLrIr6pWc0IwYcX2UxxE0V+DMWktGySfA+qD487AgWBEU
ok5inJQ/hwFMAPMlzPRBl6rMDfVKdPbZzDzsI/wzpJCIIX3U10WlxtQj+ETkWb8+
N0POzUlDa7iyAF0n5/uX8pnHBgZMLJUYYp73Q2zC8hfrxYUEAiHX8eOrsoLxeQ2q
rTaLwpc4QqfESU90prc9BlzJTCaXuoQ7ecSPjSrw7fLuHRFhWRFTK7196p5jGxqG
UCt1NnMbrxqGo3MvyJHwSiGwpnKePzrAFqmrjsfwz5azdLRw/ar0Bv7Mmyf+6dOp
ijPJr31KYIl8niAavzJuUo+yRttNhMafPS/GCpPlutnvD4s1tSSfhKfZ/CRMjnV3
pC0Ska1a1Li9PPKGmNaMc6dTgX6ju3nVOBFJHfR2U+JfifVVT7vyrC+yJv75CDR9
xvDYe1GgFxXAtxo5p4O2iyB15r37522ZbQI2L56Hf8bWn7LqIG9jRxhGaVsA4zxj
kvekspTH3/ZDERm3Jruj7daDEnemxaO+7vxgZkVuc19CMV6ra6j4jzVPfcTUtR2d
dir5gTT76FBQTv/G6Sj/+yPtd/44Y9wklj1U5dgThGCuCj4G3Wg9bsw6t2FQgTYw
FDdO74StthQ3DGHeV8KMTfWB/meen8RcYuj34LR4G0rR62cRFpwQsgxzCoKqMiNx
7QnwQippliOdsezIhkCJ4eASJ01BvRfXf68JwsWKWXdQjE9rTahARtcfG+9MEWac
qqp355oWde9UuTlAPUaem/I8hxk+HaMayo/jSYlu/vdOsUrqvI4m/kiK2Yty243R
G7JivZ1l0JgZyNEYsiJHAqRqnQI91LASvePlfTjwBYQax1rdVf92MvxNKi3ZSU/j
3t8KxRtxadq8PiJ8uoNIh8KXL5v1yGh8H3TkfidH+jFin8Mw8U5j0esNKeSGuCWA
K+ACNxyiT356tgyJ6BKIWCZuCRlZEiud/6nvCqIX/pZVNnlNrfz9TMoYJbAoxlyT
AXfRhLLPv4MObK2rB5b2EEUONx/sDELnBJC5/00Q7b1F3SLZ7hSQ0DDezS9jD7ca
voz5V/Ju7qqBQQeg4aQaloz5A10UepGnM5L5BLw6TrjhhKK1wUhbiISU9mQv7ije
vfGs7VyX0WjaBWoAUbVFqkMeqMYPYoYt09h2Ww37nLWK4QKo3kOWo9dTczqyIY9t
DeoFMOOgClinxsxAqr3y9boVcwpMMpRkK4JRD/0BfyetzJ9Rzjj3WBfv99OLI9pT
pkGJJt+6PSMWNzQyIc//L0zlgThqTvHa6MkAAYEozF/02t3aTVvMsJbaShkYuMYE
IEYKP4Mpzem6PXCyPb9C09JgeTwj0+TX2inXGVXLzcSS77vFUq2AL31u3YicuP7D
YfZoZM3M18mqUs1bHJ1oir+mPh22Hir1lr+YBVry0Dj32YHw2x+haSunCpH1NYDx
6t5/fCz1wSpd681/lClFV0Vpf5O4MP050NUnts4X/KWkVfKr+/tIoDJxLa0wLcvO
9pgBIEzjXPG4kj//gh0EDwd6kBZPAV4g8YFkrA9PgpHf68DETstYNMI1lzueyXK0
gC51koTm5q18ReMte4Fh588WszBH1023AcQsr2zw+gnhXUvnwCK2Imi3SK/ErKs0
4CMVDU7sy9MdrY1NT9heLl+E3/tjNHK4JgkwAwwgkZbkdryQU5vWJNiFc2h84LkP
ufyAAAIcXnoZuBTzemBHJcktDH5PbCgpcSYj3u71RRspToRZz7Tg5+FheY1kVn8L
Edds9kyCDdNCjpiUO8T/TDQRUukHZ49J6Si1Jcw449Ihv6PcUSuT//XKChh7fjej
W623g9EH7UgUl3HZ2/eGqxmUhdZ2K28CzSQMN67+5I9T/7Rs/4Jd3i4SjW0ifZmI
tpKMbwM1aXBC2au9Gbg/VSVgPUDaJ2K3XI0VjBMqhvRP8WA21APZMtG+M1ciqaQl
COjfroKvZFxDXvWXp3tRrjdNqwATckYZdeSgUYqbGOXwjq1Ta6NpAG8dY9AMfo0M
lOpgjBLQi3HyWj2sTUDh/J+3mgHmPzjoioGQQbaSZWyHLGg3u9v67eP7ZRWG8sfN
a2P578kaB27bDVMfDrsknB73Gz7kA0v9jOz5sc0KhU6XkRNKo+1PeaLoLQgH6kSc
OYR/gP7L0ldGljpFWHzPkgMJ+JI4AKdV7xwt5ZPVsthAEmmiMVNygyZtuBtyU/CI
Jv23a2PO/aII5LABY384Bsy6o3FOgRrmp1NDUMsx6XxSK3ISe7piWcflQT+bWGGp
EEKTUDAZ5H63ehosiZJqug==
`pragma protect end_protected
