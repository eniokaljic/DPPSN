// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LD0HN/+TgwYwvKQ8JvE3URmnpqXf8bcovmCF7fuJOtdnOPJCY/pj73bGz6UX/vpy
7atr3IcYe5U1k1I/0bAo5UbVJj9vyro1g81eBMkq4APxUaNzZrhgj2Gc8NCmH7Q2
zeWbmjr7zIGgarTEU1oZ0ek+3LK18RpECcFHicBh/G8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 195920)
TKrvBD5L/HcL0i318lXiSDC3MVYX1To/1AjsOUAOylODZxTbopJ8DVm12f/bywkl
/E+pTJAB9vFyRz20VCRdNQ8bdlwFrxUzwbm4iLAkhHG3G6jG8ReMt84yGABitYNZ
wYo0vN18Czb8v6wLG798a6E4k/uFS96JTjImZ48NQuqMAl0BtrWp8xfY6KRtoZsT
GYX8rm2pzPJTKOPHct7KHdwGxyh3J166IXsPqN50qfqrPuBOKZqNKL2zSqEvwNaT
Im4oU24Vpzu+FX+BvfD7s4rMXqxyeullgncQawwuJrHw0TegljlX/QgECZj3FRxY
ktC7Doa/rHBc7Jtb3xutDVZQoInwjwf6JGhlFNEhm+AtXo9smt+3bdZiYvr4m2XC
JE5kPtgbP9KQ702x6j1Cz3XaL9E8UB91ylTSlMcJvyEc2tKGsmod3aaSkueWlv7M
aiyVT2De2VkUUEsjiS9TXjZvtIJco1hSKXrP93xaWyZ791kPUbbmhx9gKIkb0Kl8
KYwzfliuVbcxBag18wAgtnffzealOSfnski0kHU1MpIvHCog4oVuci5Sm7kCeF2r
+wimI6DV2QpSQFIXQB64GFimvllZrAy/0JZ9EDKBE/qa9iOsofiISor8EDdWZM4x
Mkht/ZIGFq2VvGtpkp0vjrvMFizsHO4RivMO5VVlbjNxLYuPfuA5ny0uHkO3iwNJ
ZbgXtnL6PtVBlPdxxdviUe5nY+TbNkmpp59+Rr1nOQgWTg8lHZ9BFBEPD0ncS9Ie
UCiSs+JzO0juuqb4wWQIEuk6S8T2Mn5CvM2ZXtrAflRoOLY7fqC0F52hrFXPQN3p
NVa+TvR0rkJfM5ZpLVhV5HDfiM14bdD0uI7SEkDI9dnHZmfRefTYKxMkB5QAN+C9
oFa9eNRjZYiGoNaVrTFj0XuXjNDSvIBMTBDQKm0L+Btlls4JYIy4Ex3O99kNC7bg
TW/lPsDAQdSd48BCexql4jX6u/LWtH7I3LDggrdFpIoK2iMgIYkF9DGva0VOr+6e
4DaNaRcWD06gW9OrlxXv9QzhgCrbT07u7wGwfNBqkypP08vJ6rRxrKBuig6vWhwx
9FVaeQzbXsJTLz46Nnt1CKg++DaZNw5kbb7vks382iYMIjDUv8RwY+TcgJg4TDwG
fucXjV4ukGNuRgMRCT3Q9heMsqMhLaKT5Sn/kCSaHAAX5zLqTcnsNWVYwPeVdWxh
NL4m591XMpAn7yJdCpnsZU0jtvWmemFokLkdvalP0AyX1C5zUsYty01rcyPAVRzb
kM1Z9Hdhb61CYERWSY9G9s4X4h2CZlb4CGPK1pEnESFhL552h2AWfZ/QiZ2w8WLV
i77vGFn24dOUTc+NM7y0uh57DsQD44ioOv5SGX3t1s3BspL/wRTcYD4MPiUaO7zP
WVmM61Qcu7uJg+mssuBPiruCJy07deO//JRjTin9isuRu5JNe429Vq1Tr7jjnc+2
Fg8CjJW799+uwArFCOoXcHnFhGW13WADqX9lI/wLOC19/JW6EuW8DdDq2v89TP/H
Yr8ub3fz8dji+/GwCMzfS1tWB4Drd0stoJ4PsnOVe1+6goNjVD8j5UcXBa1vU1eU
ojW+aKYqytlRINTO+b4S1iFIIw15bGk10d3C0aTsaA1tmsXYc25v3R90XtP4eBtV
B4sOdGWJ9I0QkDFxJ1l1h8727WTPgzaFR15XMNm7AwfdDTYPQmT3fli5XRUQDsuN
OdEDPEhXWT8kkj3zQA/RPXMmKp8udLNgEZ1GI/YuIjUwPCgREgIB08LJZrUQv/oh
7T3NYl1egKxWlYs1OFrJmF+EKkacQxe3INO4KMOMBQXuN6WE+ONGM0p2YwddaUpO
9Ca80N1hW+lzL52L5nguerEkxbjamKHwjNMpkZZ6NhtaHAwAln6Nrguntf5ba4zE
QlVXBfi3tPpJf1NIQH+Qi9VH+PHsfi4AI0FlQLl1wim/BNTvjMxgD7hkIFblXjWt
QeUrt5Dp6yjQ7f7w5EUFhzoqIS1P9fFInAbkoV0pZffTivAq2NaC6Jti+HWbbqQQ
p1d6gMEQmlBCHL+6jIkfmqFOY5+0xlAcywlubqLMp0oPl6YRFJFiROUPC5peG4M7
JVpIwbCD99/sroJTFq7mPb2q3Z2rYXrbcTRABwzsn15n/50PigfavbkHnx3eAI+m
9RbDM90mQrVLhedt0JKfTHF2pWWaf8EPMMFfMgMXn3TqJtPbQ9QoiDjZxbUvSs8P
rE39pPku8/xhXLB8eQqX3YCSlguiKmvqzF94GvTtZx5SWG23bziVrxDBAlTZMtVM
kzaxtxxUfYuItFS8WoxJaNLR/PeHLUw2HxQlhXi3XEGywRa7+878Ff0cfsi9gLVn
/qTaDGRNy5xYMURrrb0u7edUSKU6/FDh9zTpsTdfqPiIgvudBy0jlWE0Dr4rSE0V
Q9g3MvV7WrqsX2VkTpkGg2Xexk2Npe6OAkq7btLXTjNmsMeKICiid8AuvgsbEh55
UA3fHvAr0Ha593E74KJDwWNsU19woTfvMGeyt5bjES2UeqhfkmDCfN/+MAS6rAxt
459oGqh5Zse6El6zpy9Jh10WdYI//Xb8TY8HA8/ToevwERPp4Wevt7OeBR+RVLqF
G5qaRDU1OAXIDciU7r96tkMn2jJQLUc2vWl2rBevW+0dxTJfZC+TQEP00Ew/sUG8
NfaYx07eM6hPXn7ycI/irQxLxUoRcGOTT/H5PI/hfGG8+/dJzW/3oxGhbQx1n6Yr
mdAMyeg26Ug3CXfEis0/7alkynQKJ+9vq3eIYDHhiPVaks2gNXjFrhJracen/bZP
TX1hK6G504f6p85Eg77iDo+25jBiZML2KxAfygip9Di5WWHjLgefwOMgrixZ1Wsh
/HrKECFhyhmEHHBL8OpDsWYu+0l2RAIZIjErJsd4F+daAW+blnKTv3K4EYavq203
2w8q4fa7hb3gvWLS1Al+wPNUU6Y0HahdYGGwKGbsHjGp42jq3RMof6f8UZVMyReL
mrOth3CP+Uf0NDID+EgSdLkhJXKUMAB2sLxcGwqqOGqKYWbaeVE0aWCkdCGw6NY+
uwN8MKWu+p+CEBK+SM0XUuDs5VM/lKEsvoMqlyUci71IYqd2945b6Hbl6s2nONX6
R2ZmB0xxa3YZmNdSKHWfzXy0KRYRLsuZJNWLXdjx+0obvdfBM1Pj/M6zQ1fkoJgs
YgoKtnH2T13PSJGlfavQkKu5gDgIQ0TS5ZErPysLRSdyZSErPGJ2CKib0x9sRl+g
MiYozpUEBgB8kgEM5SttLz1yTnHERRKjhwao0lIl9Eytlof6wvzzAW0Y8Sdk4Wp5
U/2y18edb/voVeCSlUOd4SHAVm7LEbDsxKDf2ONF/ffG410DcPmVyjRHpz/9eEgH
d13R3PmKYjH+t0cPJcOWvepdl3lqaOQuz0qsJ1Mc9m/Ciku/IhbOx46vj3eKjfpN
SSiUcAs2XsnsTeJDbjFe5x8TztUKuQcY9xUWDl11Tj0DVKrPL3IlOQyrIGt0pnl4
FKGsU7n1h5XFeCq+ZXmgIhD07pgBCL/OhnABTOo1NDFq3zXXCN2j/MO8dkEod+UK
dN9UePYi3Ta967sVg3BzF5M7OaGTqFoQmyUFCvzIGkei7F/sev1ph0S1lvKK5wln
NUYEd7s4b6lxmxpmHBCIR/2SMCP287mCfDzRhyj8m8IUZICG76pq4sMh1qpB+nQ4
/hZS/zZflsZCiNixy/L4yseZqFI94k0RTH/i5dZAVGynLWSnJvaDfNGe2Y58UORl
3IeOAw3FrAQe8ipARxGAbENs3oLyNIUk9wYY/EmmPL0YIBo2/V/nkAOVgkwxicrC
d6JwhcWSMkRIcx6BZvbsw9CF+zJfmKYJZNZovebPTvGk51eDsABBC2y7shnHyiR2
LpqyQsdUiIAAT3lhYPhknrkeDqe7uNeW/nGrsI797l98neW7ELAGw5BBNeukH78r
k9ishtmKlCU4aOZJpMavkgSP/2vsiYOmCBboREut4QOQ+fCeTr9LEeX7fqvOUZ8C
xyhr3gTRGBisjkrNu2xNaoHAMq77bY3PgHkeOtQPLqx6lpi+mf22o3h4TLlzLp3H
GfyuIY2m19ZqdrEWKCb8jiCpaJX2NDOvioG04wUr+Up6xmaXYzxeDcKCvjN9c1iB
5BzRDxK3lV6AuahUPxXSWyeoxe0NEftLFDXk/Eb94ykHSNKKjQ01evWtZBGMSczd
KFJe3tB6GSlc4E4OobMePd6Lx7EXHNoMS9JaIj+564/a/90rwPv5YGNoAMSnyFLI
PBIVKQEFxJ/Doth3InLJHGSYOCUIVAYC1HKRs6UB7l4pWjC6lnjDwOUdYREb7DVg
pJKNVIJ14uIKgQF5eEVadFIjKPLCIf4QcV7hQtZtZMWYJTHYMB0aaKQF/WgxhKOj
OSMSEgja6ns34n7/Lc0kLQT20exV9KPScQ69PUschgALoxnq12ffk1NUFPHeyZIf
OzvxF2leJxRMKnZupDVmVvvoDJI07mlqRl6dTLy/LJxLXf99DFP5WcAHdN0tu3/Z
lUTNZ7+85m8JYjjHAIPMXDEWYRsuzLCkjhcSU+Mm2WUzMPJ0l4GvMv/rZQAUyKla
2v0gDv2g63Fvwf01W2YEHR1jD0jcJHp99dOt7lL+TC0U/VCSbqRnjeGvr2zVX8Vm
/7yXTUY5UD1lbFHi3sbzrS5bWgynwCfW/yMj7LNuKc2myWwnu2gy6J3pGwEEsF75
bAEzsqgCGGafMIOnM/KP/WYjC41Dm3qAV6XM+nDvxWHdEEQbhkSCF5x7PUp6tuaz
1YYTjqbtr9Gi9QAVrLgqoq5wdQYZYvRCf6WRtDe1W82KQdguxvED6McmGLbsHgqv
3VciZxnDTNeU1wbZs4vs1X7H215o2RN1zu8rOMWcWnblJNjaFnGM+1Hu808qQ+GU
X8yMlC4wG33L6sVBaBVI23iIBWCu6kxJ1hFly1S7XfUD8CpXDs1MsLlVK/A+Xryl
5jBnlrNP2fYy/4tVUwFxpfGhwqFy+IHq1X63R+OmyZEW3fp2B25bXQmLInsMcTm2
8Xw9UvzpDRtPeOfvH0F5ZOIYlIFw3ck2XE892KqmXP6ILs9TehkUVNfsbvweK/Y+
2sOqkg5O5V2cAzkKVdKZlak04I8Oui7KZZUqENTMjcy5iPBuka2YWKJ/a6yNxikh
DqoQSvX2e3tvyXNE6BSL9v5lWDqDvWTZkpFJ6nGaTinhEy6L5hFa1oPbyTSzqr1j
ET1vq0/QfLK4DgBXJaEM1NVEF+BcfYyjiyjh6U4Jnpw8w3WgoT8/+DUIA9tiCnqK
rJgfCB3WzcBwuF7sf1D3sgexqPS0YyjDx3eqE441+ReaOqfsSn5IVCMUMLixzSXk
YGYCY6iQUbJwWuiqYlkOF9TOCpnnAGTB9KD1bSuJWJKg20fhelYBzVFRE6/lLsFk
esxMHq/vVBM4wSuLPvjzJE1JWqU7ssYBcxqbPtKJahc37AoIzG2XtJJIOY5azPsG
tfc6jYudBfDje7fDY5XmHNkRK2VqDuDE4J3P38xbAlJ1OFUL9H0ebI1fzM5XefzD
6nnAvIE+FBC8CXYRkZXShS7J+lmyUKGAj22jZAjo9As00ff9hoRt+/04onDnRHh/
B1yQE5ENV8P76ATOVbLWN23ug7J6IpCZVV3fyD7ENei3AW/TPsiYKoU5ynEGz+x+
jXl8Cz9gPhLQKce8RBswHetMAd7MNyV0fzhw9XzZjqZPG7v6GyMF2gqkN04Fpjsz
AnAOVh+3o1l6QIIxEBg0NNdGZSjirmRfCr7vEASiz18LqD2/BFFvY0BSurGIIz+I
B19fawAXl+MERQUibGEnX8RkooE3v9f+3xHaHpz3JE78ffitP/Egeul4Lom/ZdSa
Bz/eD1xJIxozh+FsU11Z4z8uJkASlMaj+Dpk0r3GHYH+PirpjB/fvuC+PjDUsEsu
5OGMVBFU8+3OYtD3Bjrfzkx1eLGhfp3V/YX9jv8dcTewbUb0+WqplZ5QhD93w+bU
ywgrEHZe7Htv92OGXJUUlISjU2OnSRuOVy1xiIGr/dn3hcAskyD/5Vb46JZ7E0Gr
3NKmzb1lpl7IOeShVkk3Gp85rnD7C/lqu2pLM2Hig2v61KZh1Lof9busQl80RlNz
MQ8se1zGp9n/rw0ZZ37DiGBQ+FF+9rJpbb5Nki6gF903YYNaUva8HTwL2xBxohCI
YtRDffCao2/tEIgFSJgMohkOvhaV6S+E/XrQseQ6sYvCiB3ysoMgaeqy8Phlh4Xi
A6iHyAPC3cXVSCWunBBfJ5CTlF3S4uRVDlufZFD44RQnyV/PkHWYA6CXXv45yLaT
k35HSamE5Z2/cgMOUnDkHuHRjMab43BxPNROuepghyxJFsVERx1m77sLrZ0ENEFZ
dCnXz7fREDwPxjYzf38Di0Q+xw2pijwUwcF7BKwIfEq36NROfzA3b7I3QP+kXYfG
J3/xrC9s64GKb5P2Us06knjxPrElYD7Oa/jZMUVoT2L67qI0N/zkGE+fx/4MfVWb
b6urleebKxNdAoUxdHfHTeyUjVEaS1i+UMViLnTyaO0BxImvwQ8ZcUhKK1nILgiC
ffhrA4BUx4HGDQ/Y2oT6eX/w4SPEmSq4TIvLn1UvBJCHRVvXjM1DWNzsMLpkxVtw
F3otkMLshkuMcRBsSExB1m2J9MDijR7PIgCiyw0x/AZRYkGz4McGr9bCVVu+HZbt
MzLr7YkriJMRXboaXqPZgRTl7FPxJgX6yaXV3ZvKmnuLtYXcqVnMOpJN2bCSgb6R
bj/3muGPQa4Yfk3loReGLqlGX085uwBwDLamyCHevFMgcy08o6XRp88ozrwWlRfK
JazVW5NSPQNU5/vbxIpUcpABu3FfGnsRr/Xxds0PraocXx1TO7SEUNoCSprBvUhY
krCAXaSozbo/JAg3Z8dVBIyCuXZudnxw9ig07vOWsQ7ImuJFrU8IOwFm4yorU+jM
tKfhUIvzPHjaH+tYlE4DVOrVTPN3CgGhf7VGoAuhQWH94NyHJ6P6Ao3UORdCstad
6hIXJIe/Xkw92PEsOD2EDPrW3SQfXUQUt7V523vnLJibD5plInxOlexJwDK6r+/C
G3MaA6fxG6CQ238kQS5ZIKnD1Fg5tkLP8Pw4Ix1mKCJP+e7dgbHqKQ7EYqWhVxcy
1T7BbbpKJCMbvrlbGupsU+bCTo3N4tcFRw6vo8dY1d8D8cLzwSsEhhFdEoBhYi8H
wOfLU1p7I1aJvpbb5Rk8UUtKfEEk/B9EOieKHA15KrldbV65IJWlmo+WUMH7RzB5
q3v69EkhdSAJdfOVUQagg7GfX6fu+VcT8bI5idnEQL6ZU0WzBzk359MW/+bAySwa
LVrLMuEvXQbYglKyjTQdeZCDv6DxIs44xeolBHu4Q4dTpzhS9xNLC1btdPTMlvhe
Q0z1VjKNAemZQn83NxIhcvCcI9hiyE4Z23rhSh0VFb5kvD8M1Ux//zzkXABbpua0
azStas5p86kHhlIAGCNnBkn3bVNRLeF2DcTpz5soaoKANkTMN5s6Me9JXSJ3Noav
HS+T/mLU78+9AHZwYYF6/ZYAiTM5CRmxNE+PBJjKDNNDNXSurTCekH/WnsK2rNJV
wtPoT3AKaxp7TP8Mkxk6JFWi2U7SP/vQz/xcmL0HbM2gMwM4Y5CpBpc8FUQYp88O
fQUCeSiwv+r+lGiM572ymM0/f38hZRD3lT82peiazvlbJ1HjcuFONQ07JE1JTZ2i
wsdShB7v5KELGmKzgafP08U+c5d36/dvo0gRfhhX/4Kbr1XuYo9k9/8icfyfREqj
ToxUxtUfbIcQUY8Lcn5+aHHBqqmRrhUaT+Rwbt9qZxAemkM70mHQgT24JGU4kk1L
tMyuWug9FykT5N9Gv4bfUyzsd9eUV0tWVLzQ4VQx/zX46btN6GGWF+8mAQTDgELN
RN/ITL7Yoxy9r6shnZTZ1JGSP5AKefA9J0g6gec7fF5ikxP22edWH1VVeeWX3eBw
se1FqMGxpSBUinZBYewJSaWPvNVlBeOxwV7SSKgDG3fXnur7Y18zKVZBbW8CwcGf
J5E1uRAv5JHbRrceWC/zapVMI2otMmfYAzsQ+9P7CVvDt5J+6UK+0+AJ6KljMd27
79BrRx7BJsUvRSTB3CZiLJ7fOkkEXjgrxNDRN005h2fYh0nlqqDcFNEo/0OPlPjd
FIKi/Id8zt9hKUFa+4fDOZeQRMdrvj5DJPshny2x2xq3BJdVXmp6ZJe2dPuoGMy5
8+MUPIdwY+wrGZAzbT4HzMvzKdOhyIxKNxY7d606C4p27GAFu58LMJxg9zVeCIt/
tR49Xp2h/Gk+P7IPDtF8G1295DAMZXtNVHKwx1LXFnL2Ds8ScbVDt5fghXKH5K+G
JRAdm6qYVBaRBruTrryGag5aQf6vpim786HuP6wDFPzvIh5/Za1A0wtLxMY3P53m
WDNiQPAUZIB9z27qudJ3U0kh+ZlyoREmi8mmN8IXoIXt8gdYmNudkAcudtHtzVPN
OhPMC9568UhVaFKuaSdCd6La/RLWMnJ7bN15Kqf0my0kbIksO2YmD/ROSsew5R8n
U+aFjPXe0KY5kZJNrYrMjBmJgwXvLCMfWRiWLCGvrZzUpw93JWZnulmeYG9NmJUT
Xs3K1m5vN2ALzkIpCfImE0Lob67aJ/hkKnED+RnVV72QMYFaX767PKadMnDHajn9
v1ZwKtSBoHRDw/urq+9pQ9VxANYEoVefmOLJgTiEr9n2lsZMP+B3pphKSBM1cAR1
949RSsZCetM4EbWlWp0AkJqyPymm40aFpAXgvR8RJkhqB/2/g0xj3hnzD+tLIAvc
+HW2XUCD+ViW+GdCxFqx79/RjcRKzfRctrcAMX02r/OwfY7ayJXeilhZCC0q1GVV
gKntaxHdBYBtuEQKR+Q8/iul1BS7NJ7ixDeGrXIZ5ALN/Q/17WsFuMUI5iqY/GlN
hUtFrHYeJlz3bPL5pZVtBmVQy4zMMUTn+fWGn/1gQdNmc68OaADe7nniDbUUmYek
oGIo65f5H6tFpprv5NSHHU7eMR6Q6QRoXpO+0f+XT69miSbRp2dATNQy3Ua2JTs4
aPyZ4MtHLgv9havuNxC9eT61xVckhZe6Y1eSF37eIltkXVACiKkgpeEPbx1JLQCU
2ngftZo+cFJPv1Ncujrx7MtISqy99+KnjsEuUl5bOy7x4NoATja5cpD7xgeDJq3H
DvJNdc7UBG+/p4w/Ata43wz+mWiRRy+3bhkoI3q2Xj+uoV7V1b4WJPsmzPeWkI9v
U8QjJKoI7HLtQtOyUJNCnZtW6MXqb0gHWVmO75x6hkbN0R15Xded0VJKbdahM/qu
JQaxp34r478gIKYwSJgZVpcbx3sU709Om0TOsmXf3TUBH6Hk3k8s7FySiNR3HACM
JBpKrcl5KDEUqVfj/8MIF6D3VwviC7rCemA2IExvky+cqIWDZg5oVPL+Lh++mhr7
2D/wYFwAYNmcyQjonHqL0ZEfATlP9crPJpXQHgx2K5DGfFOI9zt3YekXzqvbqp1y
kuQi4KKb/B5mfTtiJR1tiuWOAiXR3H/I0PQcSX6pgMzat5z/5D1wMR79glni9HRt
dsPg6vOJ+d34pKQIVqXE8MVP4qHn1WNKxvuLtanF6Chy1+64nTk1/HR4K94JNaRV
4wh/6DjabolpwlAIShPC1FmfGeJKVAnFynTlGGEZQtTEF6jBUk6k/VBv2sDAZqRp
Wa1/VVa0pKnREiqmCL/xTbpt+k1ivm+SZmMGjuZB1+EvkMnALvyOlV6mMgH3UYCp
10MCGnTc0Jt69zkmFQDwzORDn/JercCGCL/QtIyNQcFmfBddLsKICiRHVlr0O2m7
vD+4SnRoAyQOLry+AolTNrzidzvSLlr1ScJdFSh2lwUKuh53O3NlX5z2k1HDR3tY
xNtU1kIxpYPfAZj+AhOZPd9FtmKqsa0N8L85vwpzp20Kv1+8EiUH3UowbMXbXLfJ
h7V1k7XOd5gIFVa7qZ0+TTVxgVBcEVOQhR/jDfDXegB2IBRks5n+tSR3okrHRfMx
mhPPedgKlUO1GB/Kv7px4y3xO9Ar64YWdOOwARc6ZwU8MndlFO+h699hLE5UXsfb
HJFwz3X0q2ztroDLaK4AB4MPqAgQOeGPdxAwzEHBnq4TrXnQra1O8YaTYgRLK3XK
4STzLx+brQOj0v0PTEAzPP5KX3MtTbn7gKM7AtjDYp90gaqeK7jK+TCXgBHfMkVg
R79craSHKq1qVGfA7Te34lG+dByvjSFpii4obqkpAjt7vMxCDM8pt2CeHdD1vUxs
zPWTlTMgLDCoTDiWNhqUzgXSomQukvZ9YOhGgkP5jpA9Bx5x1NGPt3RX2Ea5vecG
3Tli7I9cwS9NXRNit+JS2ctfrIK7fkzSqE7NB/FKXcjOSlqrevaTDIfHoLAzDH9q
KFLMN/gMrECEi17LLdtYA8ItRwtarZouWpPgTF2OE6cf2toBXjif4HqDNV0wkqye
enZXSDNAisSytaqhWwFj7LpqrTk3U88cgvka7KRizvl76lFGWrbr/YUhsxxJybNp
Gy69FSdl/XzzwJE7QViLcpDV2tWXxS54wf3xrscRsrO+C5fexKzVKWDBd/KgDKOn
GsboR+yOx35Xqqdftgi+pQOa98oL3qwP6B7iR+NDabfyq99UoZXeWxXewmydDko7
8t82O2g2CU6gIqLsGVvAmKaFl4S1cVRr9SYUSsHzpE/967yZmYxI8eT5LHQG/4NN
1eelbUL9InsDsxDEIP0juMmR4EAyI3828u3qllOvY/COEVS1a5zMgEnsXuyuDIRj
nyW1zJvtALnbYq8jceixuTfIWTdyFgZ8PvMQ2hkaNX1E/9VOB795fUFw+EBb9tKw
nDd0JXvlpk/PJef5Y4CjD1edE3YWparmEH1XdD2Xw/ay8MQDU93yRpuzltlNCPlX
vEy7z3/tT8LRonEQoHnJn3/ylJiaojGBGWjBqJ6bcvSsLpK//wAInlhme7CAeyJU
x0TFaRrX48W127jcwJJlm1xzG+bY81sNecyJ8Gxyl5FU8qiPBtnISgf5Ba6D9wPy
JEOO4L33j5pHg9MnrLPc3gW/krAEi6sbO7HKI4OZwvdDeHicuhRJOX1Hq5cXcu56
SLU9DA/ku+RtsIzNeeKmtDbOtS5wU8kUEy467k0/st2DLxkIU08/354Yu2x3TmGn
OQoyc0AVEJImqmfYO81BOltwhfwIRaknmRijB8Mb8M+1Ltsvt/tO6ewtdxmNg9OH
M9jgc7cIUio5oLlYFGni/a0/bioobeAMa/QVi9NivdADll/K61A9MUGgDBLPu4Ce
zfPNLzmqJ3YScAQXiWeci7hMlW4Y2df8aZMHzgUw4DmRtbwYqgB4sQ0t0F7jC6q2
h7gQ70D0sjpJvZfoZsR2DGIbA7n7Th9cM1VG5FMAgSi7U59AMZP3jxsu14MC+N8b
SW0Vcmb8Wmd3iNjnZLaH/VFp5JcH9d/DTF0QOewIJJqaA8D/ATGhvhSYIcbTLGHz
/TKFSMYXeEcJytlw+GZF0LE2RjITZeatk3+la/xCid6NsyRkeTxEe2wIX8RfaPP0
7i1IiLwT3Dd+KDjj4vjT0XLmvHlYHHDClhaGK5ElwRComr4O75pVSFe4XXGoJGEh
oqnrIC69uBCZ2cYNBtZdZC/bYEIRyJf7s7fyom+fhwMwecXLxgLTswvCtcZAIHZ5
OiQfebJahVDkzaI9tSTovHHqGfivw8jXRxTBuZ8v/qMESrQgGn3gWVzDMuPPxGm+
k6FJACYQ1t/gTW8JgcHadQCw7DNi538lKPeQIk71HO8AIbPtUm5N9ffDx5MfMAUE
X7KcBlWd1Q1EoDFyxmJgvN2/o1lvbQmPxF/rkLu7R0ztr9uNFFNfke33SkK4EGCp
oHVQV1A7WFp4xISs3ntc9GblDYYbAnuukshP3ks4V526dH/5ingFCyJjwk3HBfon
TARrzkHMMU/+nLa3ZnzsHbBCcKzxHpkKVzqSsCbk68Ae8EdA909AxczLoLkMiOY8
tCwe5WCQyuQRNnWb2fJC0Tdm/KmBfTudyDZFPqNuUmpqdhTsYzubmPYMRG98BcE2
NExgX9QOu5tD1kefl7cW7ZZWq8lTOqpU1FUhm/Ke6ZAkoPsghwXN7iFOID+OdZsW
7piwuQEZq55+9xs2mVuIA9HHKF6XAk9sEaYxFCcOvpdpbESOfmke3RadStCPvj43
XHzgavS1GXpQsXV5BIyvi2tLopf9cfarMz2Bb8gwHwnE2zZral/jurCpnPdVIpeo
8YU5vqr5Em71ZRlWk4ZYK+CrFWB8CRoHb9zIqfzpFMKM0U5cZCBZF8I0LhJ9/zdX
pXme0P+TPBECDgPrkOXvy+qS7xWhCajKr0VBxGWSHRINurtVQkbGGoFjdb1DXKDW
y5g/1fg6JEiI413aFC6jISQ6fwhxXZLrNXjpbRDdPiujCT8Ou0NZNybyRjIluwDm
4jzKK4qyQjy4zXfQuw6tReSk2UD/smhGdN8vvCD6JJYaBc5xZsAqDDaC/ycSmAty
fFcEONIedr2ZgtoBvkDyrt8Kqov9WvT0xIjZ9Gdr6BNdSZzxeg6zMmJiOhZyCTJN
DW8pRfFAA9ln1kvN3HlrMn9u5KECs9DjXClQTPSboIkhxP7MxxpWqN9Gyn7u4pvq
j6U1Zg51mazmtYq/sq1IYwkJVmiI5jjeoJBCKI5S7U8hWtNW6uCI7n3EutHcSHd8
rW/Iuwdc9FT7TZ45g/hAumOFE8DE2n0YzZoMR7b/luAsQkN9TVtJa1Rgc/tf+cGz
kUSMJJN4Q3M3C2IkRJ0ZtrFUD7o61T0NscN8iYZlQeyuxNd6BGEMxCYqAfglkPnk
lmVgCsJCyzoWyr22sQ0VftVSI8v2uOrLSQ3C0VX/7mNok8NFNKuRGDNISFLElqsL
jl0sAIEGy7c8RLK4eJzepciJAAgDl0bnvVolcRL9Svp6O8rpv/B+FWga4+GHSaR6
3JVWtsbWVGNv+3Lnzn8DSnqaW/PjqOElV38XEYw7ZektrE/N/Q+fn+od5LQ4J3xt
wKdSWGBJ2rSVLoQUQM6UFZR2okm+p3515q/dwv2BGjWXz2FE2+YkAE1Ddt4/m7cg
JGZLwrFx76pOYSazRKEDwQZczwRo+Iotwsh61hzPRVc9ClUQj/2szC0RRfB3nsdf
HfdE5v0/y8c28S/fVmArVYPz+eaNd6MgcME1RhkvOCWQtsy44pOuEESDFHBWi+aB
39CnpHoAQfGViTq5YNH12U6r02kTgik03gCHv/Yb+waeVQfCepMPIVVxIYrBi0Eu
ujIodcx3nocQQXtchJUg95u3Vt//2Z7eskNfObShG5335l/1OMw9R5ltQnrjw/+O
99V1gWkBHN1Wzu/0oyVhmvtouO+G5mkZ1TyJI8jLs45/jY8CSTXdxkZO52zbkiHH
dTRqiXSu8RR2u7v1+LTpsYlVgtBTOvNPpUjMfaMFWIDwQkVrBoFK8mrwk5cptx8s
tMjfv/BtA3/Cpr73+xWnqDjdJdVbPwMXflfVCgs+5+tXWk/PULronSDC+hom2Upw
G8QPctsTeNDL3h76Rg8aPXwkak2SmJatv1H2DU5hp3mUDpYbelsc1E37rhpIbgXs
gb55nihK0sSAyqv/MC7chQMTEz+1RGNDL+uUgqgR12nUGlhcR34d9u1o2IamBJ7q
vlVOFN31q43saUOBAwhQ9Ydo8aCakqCxzUWL/ljt/J8xlSEycqGv0yAn+qw0vxPm
nsSeCA71ioMWAs9j7rFNmgyAc6J1yKuvvdSk3MBbBDvQMEChmD/YntYh6kaS+So1
wDOGYI5gTJ7zxnvqxhqbITeOfwqpWeyQSEqcTTa5y8+SSg8q3e9z6C/vtoIsuhEV
JaN1RiaFqdSgWsMxSD/zf4WLLGSvi+GdIfnEAL377sEbDVQpHQS6oAkX3QZW3kD+
L7kcEDfhGzEwZbXWuHAU7NhnPACBqbySTrsWKNrlNO9knvZRvCHrLwxGcq8F7HYG
c7AOgmQDPZMZJXE3BKyYAJ3gv2pkBJU9ocQsxo6DXpYcvxNgHC7iCjn75B7U3sw/
zZC56Qq9E6IB7UHFNT9uPfjuFY4ZmyroZhamimpjilf4g4CecTgO6OnvKobBzhz4
Eo7yYmEOMJwfwBafOwL9A8vR3asOnZZN4WmH4OEnUCI9u4w/uOwtk+5Lqs9NCSQ/
0+b1l1pwa1SP6HJtGAqS8C+VAoc0fm0PtKkx8ez0YPAzEjtQOzJDwStzlYVggXjB
f9SiZg6FhCBHwvShq37eqUQ1QbdTdju2LkVjPKlt6diGBt/bolRTUiuN54QxJ0uB
om13n+kJGoikEKsQm1pCQAWCLiI+Bupy2hnVqz+EX+ZNpfPHXWruW/079pSzYud9
9vtEyYa4V/+kBjCPO/XTQn5JlOLPzLwTWuCIASnk82xFDsJ/YQLguNnVBMllKx8u
f6wks75sgTD90Otno5cfH9fKMyhLH0riZIPKb9sqH5VFl7QIn1BO6UpoExDQTSvV
aB50wK4vsj2dRifSv4zDljGKUy+qT/3YDx++d89Q2ey6V+JEcexk5eM52uLGCccm
gZb68id/raTMQs5ZzouIOe6V1mSeBZ+9X3rd+/Aszv3j1ZXCgxU/Y6c8ZZ1TE2So
u4vAXeuEyMt/Mgzflve4//BXR9UXgz5WlLvFh4MZ/WICTx9R9ODl2PS48btBeOva
h8i4VNkCRjIIdMp1ew7nHjLUkD4/zQUj1C0BRM+1j8Y0HsIVN9XgpGROzyNIbPkx
bEsiUdi3DVyO3beKMJiD83qwhiNucZmyDkbg/GSTZI/vHL9glsGUS0SJ6yXJWPA0
/VvrkIRTSu3QrygeQR+WMBDBF6MKe6tUwFNE906656ZWejrUUAAdaCR/C/y0MWkq
p7h3nVXoCJT4TukM+U42Cw8QiEA1dCOEueaDqsnWSD9JvGrEBNHdfbF6xJYu/iP3
RENUtVktXiZH9Gd/YrasVaAOXCxDuCJH8PKwgtiYfPRwbsMYCMxU9RNY337xqXP2
70zxZ3bCwc+I/ueoAwYNGWADwwtwRiJ6XSAtalzlha8gt66oTe2ZpBu4lfjHoaNu
XZTDNsjEKrHyOZlNgVUdLuMShS0XFHZZ4sxjZbWPhGZNcxgIZh/NSQLOD5gnSMGL
wwkAdLCWA8o2hFp8TkJHTcDzVo1lZFfHbocgNLG8UwcWzcYChJ0r3rFGuO8USk1u
piBZrKN9mxlI8vNc8X6Ba/uAZPs+tMkyB+OApAhQhMDn0rIJGReNZ1CMt1jNTxeh
M0kf+xjFa3FKhX9SKo2hMEr0g2lAlGVupOnz8GQKZIUTb1sYA6AL39s4C7vxLYds
tLyYotc0Yfe842LituZ/iFzUbeVKcPY9sddBUGSqAVa4B9jm+elOtmkVwdrOb2Z2
Fj1RUb2tUHaCDy4iaML2VzN64Sl5zlpNdCY4KMcZ5NVEZ1AzGFlQ/vBl7oSAvODP
YG24/0IPYRc2vOdWlYneb6NDiyd8JPzKd0JggPvFqXwAs98vauK3/cpEd4VbI/d0
dbQjFI21JyhPGZldZk4fAWM6G8Q07WpRAunVq7LpLhq5Wxpp2oxVCPnHETFxQkfW
ZzWfzU52lRS4jYs7AzDRriNPZhRXhOPW+PihvUPcRK5jZQnH837wPSI2mvkpnrmI
j6PDfWY3jTLuHS8/E9EAEJ/75Xt0mSoOZ9DSiy8xAgE/2JL3jNugssXvhhWCpBYF
40szLH80nwt7uAKpienLJEbgVpvM190lCcA5+eEA5ZTi7HGfv/Au2h27LTRRoZWd
o8F9uzAaRHbvwCrbH8s72ns70o/aYYV5Kkb1rDL2ES7fC/vh4tqEnZ6K9FvkaLxu
iz+F7iXfVklQEuh79txGIG8XdiNkKw5haKtfouMc04jtiQm7/VSCKcDb4Comw+3t
vL+iTqMgmqBwOEyrJMPpOdXqt7Nqy6pIA0bLx5vowAlSGGH8czAbDHZiKOTH9UgW
+2gTEoymeAbm8oUhFGXXADYYEf21al2GA5SI4cYntPNOYS+zO0Oi+q3aAZWfjhrq
dyAvkcEbFNDTlZSoSnKCzKw1VJeMy0ElLGrfMhYW3hCT+lauFR5sAxsNXwGw+xvq
C7HoqlCV/GmnQCikOg4IMtQwbmAkviGRWl55PWOKVnjdWQ0aQHe+4cNoj6jX0kQW
wiyL/oEcZyS5SN0S5WevDuJZj/YfcpYidW4Uijxz+l/T2O5CCso9d2ZPpvGk7UB3
5dTt7xlASuh7/1Jj6QvwvUDwQU7RXmptmMXcbN2ZYoy78qpz7AzQDPEx5KuSj1w4
O6ImZYYOHc6Ble6kvWQM3UzVghM3G9iVTev9voPHLItYA09GDouFWxChWCYb4SLg
Cw11pYz0V9Jx5WdEhaMrs34SZPtnrOw3Bf8Znp5leZakiWpTYThe1xN2KEOt9QY3
uXFbn1rR+6WkyUo4fXbNuEBNWXNxNLjIFy775Ep/BT0S8hNe0si8DkcNvEZXPi7O
m3QK1cY+SGWgSIyy6JtVzI8eNXDylfvc6GCjycomfJHrJQnZT4yEpQmn0CisL5Tw
yMc6IlAxR0DnDMzte2Xdu3RyROUlqY4c1N7XyPjxL0yeDEUoKaDx1sp3mXKGb4uO
IZH/EpBKSdQOztypekBaYS96r9wsomP2iTdjJCwMzYwaA65MW/IzEJlMGkC9fS0t
AOKibmXzHWRjA3M8txTfhht+hT7g+6q0RFYbuuysmex5Qrz1F8XWrKUgWRBfcRH1
uwySQ155Xkz00psYbxkuOLNCYrITMEDQyN7TIpG1WEd5H6nrZM77ZwB6/Vqos6sy
J2u5JVEhWipVSNsyMtJapZzNWGu6z7eLgESoAyeNcSK0BhY+KUyKh4n6q4xrhjfX
DKjThMkz+QAEOLCgXSqHCuH1bVLLnjzu00P8rnkqVdu4uG0VDWldKVPDZB6LPkK/
Joe0DcddlYTgyItpVWRCPOxlgskb4b8+3ju+mUbHvHWJoKeIx79syLbboW/pz10s
KBPHSGIZdZn7QyhXRIJRJWzYDu901gHd343bVWWwSQyCxLGPQwbk+Q44LBbL0Cjd
9h13yDe6DtuEf0d6jmO7PFRG5TBnTedFPUVwslhpDui2pBamKClWprcs+6PaIJBP
NouSnsLk0PT9TcDAoYl7WYbUQDFAMzdOrTJesx/94qKDHtz22nS75ROCW2n7qNE2
zKDLsfCdrHr/z45/FVuwDOfVjX/aUpTFAAfun8FYntSHommV76TmBkAyGdROnob8
e1hCt5ywDi1ntIA7xypvD18w69FFSnd9aCVbvxSKk6Yze04FCoSQApr3O1Heivdd
Zx9+5WG/XoVYggPIczwqdymV/WJo9t4x+F+SrVuXksz/lkZUU7T25Dna5+j9SH9q
WthPMMKUfBwoQcpjzCV7Px9Q+9pWPoqbfnZTdNZMjnckvU18WJf4UGgUKPejqZA0
CjSESN6b4IVNALD/HKHm2SWJdbWl1ISWKi9gRd7Nqz+kY84aRfnlwlWUpe/2zm1B
d8z7vRvOLxL4qeoJ2dx2Je+YF2PambX64RSeCVL3Pp7bqL1Rh7IBIVoeCFgT6Zz9
vCghP75ZuqeXDnSZG9F+5l/e1O18F+r/b+oxaoiivobCrlwGeQdYNXYcXmXOdx7r
+8yqUALNrh6qPDvIq7qf/guLrT0LvlRnHPBL//oYHFZ+87oflhUcbdiGW/G7lygQ
x4o+9Dk8RcyJzk/LJ1BHfNNwzIpGjPki2zDcLXVzSR246Py35TJ3th/5jJf3dTR4
PuQAHR/Fs6SRIe6Ib6dzoxW1YlqZpTK8y/OrORQ3preN9u69E8jDdTDikJevWs96
8TrtUGGQGL+3+zqcnBzCBLxJ4ihKZOH+1whoHiSDqagzi2kGbTipP01qK1+xpZse
0ZbvygiwFmguxPQ8Q+8KIt5c5Jcuesqbmh1laDCCkkAHMU468hfAmUl1JE9sz0C1
T8wH5lUsfooxIDTQyyzNR9WSZaflGtd7HZJQJm09gez9Up5kYj4XxyVTGHATGNvm
+G4oOzFdZKjWBhu1joPO7aU7ekm9iV855iq3v1yWwLmZVpwYpY9iB+G+c8EFIpPE
l9xsWguOlPWRGp1OpyS1DYlNcZuwv+S9uiLm63yXZCGVsjDDiNAHlA8kvIFZbSn9
5W9mwrEAhxc3xiFPahN9AWL9T2g72anAkpg2lj31IHQ0pVmMNaZ2jx6CwCpWSQpP
+GvnuaPyfMGx6ZocqDNeLMVYyc7hIE9D63LcHNLPYRabiqk1QrLwvgR15mYvn0K5
hhzZ2t0WCoYsGSSxa6rDbhpCQdMO3QRjHoujAWcA6v1vbSPjTkSIeBMuAnVmU7x9
75Rolkyznv5um2R+hQzz1nbHK6/W3PahBU5vWLPyvMF8GsI5bnbpCwStepNBTMCG
25yDz6AB5BmXJOymr9w9t8c4U1UI0NBadlaeuZxPtm4ohd5drA8sFkzxniXPXJ1h
ghqo4VXWHyDvbJ1uUKf0NOdgALS7FZqy1aaLj1AVeCGVF0MQEXpkp5G0Gj5Psc9s
xREyXqMg1zHme2UUmJtHD5xsFBURZBdLGO0lbdGp5qXBRASi1EI2yGeA8K06qBvS
mhQYoUJXkaRJsaGKvYNLc22JrGnIJZz+mgFJQi1O6tPgZuuvKtG+ZT6veRjAnuOX
+3HLdzK+CsQwf3SsVZHegsyYXN97zHQdes8G0it3FbvY3WNkZsvyXQtQP7Z2BhIh
J26W4Y2ftIsAoZJ9htRio77R0Lpr43ihYlQFfgYZpBcRfVGMnsM//EeeBle/ky6y
w1/QDHmhnKA1kLHuSyhmbKdJKBVOLjMaA1wZ21mXtppPI3+kCH2cXyqU/W2ZiZc5
bDktdlCc6vnUJ22tjWKvR6zJmxk8zIRUIrmmsGyOkm6jrcg4gvt3C3me7jzGIDAz
QvjLK9n1a9sL8BJUUicLFQWlhFYCagS1H0CoYN2BloAFFaL5GKukWFzm+3xSLxvw
UwdiDRJ0rlXcx5ckM3fsb7GvqPlKhZIVEKlFTRw20VKY0ESH4Vk4Icuk+FFpdkek
HXBHOJolUHKzGM4dZv49oeUKNDURVTM8rm+S9EKGhZ8MD4Jcn0vJt2w6tGAiPf7g
bXSpseBlqxKvc7c1gQR2cQ/lDouu2QWUwKtGLqHv5o2x6Hxqej3Clp7cWP9a2JJ1
I9LRYRSdYj6KEWXjkaehln2JT/9QIUop48gIdVGNKblapgI2HvY+WN/lteFiXKw8
P2Ya7pnL+9SGouCLmJnyl97kjLK1gGs5QMsnroElnmnvgaMgzhE5a2AfbmYGiV2a
IDCVrIuroZ8Z+mNrLzkqh/qm/gsZ/yYBJdIEOXHXtPLuCK1QaF9aUiYj77fhNbdT
FuOeDv93NEXorYN0Gufs9QEF0UJaWSBsWEXk54iHC8GAkXTwA0tZAtZ7hvLfGKz1
EnuBlqZ9DwvU+hQ3kLeBMB34lXYIuQgHsP/px9NeTbdcg07lzkxNHtRCLW7MCu3X
fHH7OHknO8F1dev5kuP9nDBg9j2Vgu+vY30S+0RxpJd9aWuQ7mcGDd1iGOphqUbz
WFIS3yQJXw+zznIlw4UgT8vV7/K+Axyp5OaoLiVTGwgvw4FtPC3kBz6pmv1LuVmb
boKUCj/gWpyoWDu1qz4mSVv1Z/kRy4Ya/UJyYhtJsKjU3yiKO5CC0ppgcmVIpNkV
MdIiKEFoYtVRkkAuK97rfHYahp1XREsWg1X/UPpxfXce8FkOe52TAG8elwiF+dLG
D8RaJSvNjvgaExEsUJV/hq+KrpcsA4iuXcQSVvBcQ+87zuWBstJqfSAz8rd7ahQG
YMSh8UTayqCTx8hhiqI9JsYq93T4nA+Ntzds/E6nLi5eVPDiwACiLbSSPknGbhPH
DnWhcBrx3ANIOpzOnOQ+zukxwP9JXqmrZqW1blKF1pFXX4/hmy+e1Bqcixm/aWJl
2IYGqbsKPgPCwcsH67liy42wC5yyDmGPt3DNn6wzeK3+It630yNPrrzb7jRUEe/C
JputM11KpUcg6Q62ubJ3Y5cwzAO+a3SePzN8BBOoeQCcEu5N6OgSITPHN0lAzDYp
VIilPjax9Fux51w31khm8n4YQ4RqZx2hD397RsAY+fq4ZnZfX7oO7wPrsxhlknQl
Wxw4fL630qcLzpvxkj3asIM/CVk5bCiemHTTyMdhMahhOPduRLFm3vHjGUFMbgVQ
xvQ1DGZTwMQkbe4IA9RjoNq7Iq5kwCeNRU+PM0/AQ0vn8qJBRZQPc5AlpQBcVMW6
8lJv3N0BFeDgip/2cqkwdefO2x/WFK/A+mRqDK0PRYOxfZcJ37yq2TLIMsXBt4AH
RI72k38sFQLO6FMArC994mdPEUNUukwArsF6MIF9rQd6jXux4V3KhYsDF4snHUzt
HxC8NgO+nztBXmVhw027dJOt55olnQTArJtPdhig39It3psQQmdiHacHW5Vt6siO
X0HOU+a1fVbiyDaX0zbDASzDh/bv3o9R7tHTZHtrMd3crLQ/ychzhKVM/m9WO4n5
Nx9e25C0n9Lgb9ravrWqQwyD2H5Kd8ucZjAyNPHwI0iALnZy1qT2VU9mUBMirKju
58mDX/njES4D3k1hMyq1hZ/nIWTO87JAZRG/5vbRQMxt4OqEzAriYTIyQUozw5yV
Pb32YUzq01glVENnquxNjlYh4yEFLENYDCSMLUWr4gzsRMKbG4qk2lnJZXVryONL
ubqxcc+HBfrT/wxMbR6f8OtBzyJtmmCtzvaRXllZK8npZfv6nTGQWGZWrggFR8Yh
nCNE4LjBcwpr6XWzJFZ4/+9mrIgas1/cyPDMCS3bQ3PGXF2pqjpauxaz2MnzylNJ
3KMWeBB/3P5QODkY+iBcFZMPLbyMvNB9ssAfqRQpMtZdCRgO4slm7uymQXtYIP7j
2P7wgZ6GhWlhOvcSga7f+0+VeKWCKv+vOlCnGR6kJm23fwYs9vq0tpXLGOK9NwEV
hnaDSSGufMf34DHSf162m8WEl9LaI07qnDbhdr9T4ZuxQ6NVIi7UyIndvgvtIo3I
BbihnoiXW5RIZXDxSJJNb7FKOaTFgczLgQDaqR8EP0GhDM6SnDoddlNIPj/pS0cP
dRvmBcKDHDLnkqo4ieqfj54ZapmZAiiZc0jW/HWeH1LoeRp+UO/81KkYbSjUT0WE
ESt2Frt1nGx8MiT/kyg16WlMe51/JY3naUjFI8boia1wEiUEmSfkDKax6kYdx2uG
SecFOI/1ROELxBk5luer+PrwCu+o3RMHPI7N3WtKdiACCk100YpMKSBQ7tAZNh9r
bsPEHVn9wJRGFd3jCNoQDXZF57fP1CyyGdr7CX2aZePxkQOII05eJoZETe3LBY2F
QUQq8TWXMQsqhqtgC4yT32xmTCybthNidwV8BiJYglkV8+GrM3M4R2GoYUs/5tW6
bQUdnd4E8rx0bEx/0vG0tHIkVHlQ98jn3xiwolD5VoRTJvYBQzJuHt7mhcFoPhSJ
584SCe02aBVvVWVjH5sLhoMCk4EpHzswDWBxb8DCvEwGf0UbJPs0CavwolhGirHk
zHV0gkfLah93D6m1KffmeN7UKuNgMSzqMp1RCPH1/JxTkLEfCHPnk1GJ3MIuInm1
Yhh10hSi8A2Ahd1fm5fUv7kbk160bReKMjs7ZlOOzxdVY84PmrHTh6CTaiLeC0/O
pmxuj9YVjuT3mDNu2O/xbBGYMsiYL2m8R+x3a9ChGP1BUtkTx8p2pb8odZpzFoQ8
wtEfSr+qrUIQ0EynA26bQaL4PZpPEPgdCqEGaVfKMQxJNxFomDMgJ0b16BMjgbYn
AtXzTCAdzfwGln3ao5TN7r5P8KuVTgnK86/LEkd+HDiBgzoemyZ47Dzf+rqSkkYX
qxfmDxP2i7mGrRzqRnwstmjhiUvDYLGMVgpNE9PlhTLy3GE/NhQJUYS8iKKRPPpt
EZi33p2steTmH+/lHxlebSd8zvv0uK7gFGtwSM4fCZsliCwrz6DnHHiwaIbozAp2
3eAXeK9NJMVJ4Y37ruG1ObVSEfQHZ5/Vy/bTkK0YrjlYwNwyBtlHls05SNyv0P6M
Vox5ERg663G8S2j1eoWY7szJiXdntqYPkmTqMgRBPrxdUelO8580b2t8WCf4VCpQ
UOYbd7Pmghuh+fTlZrLm0EHjoAQ0Z0QEFeizFqv7KHsZ1PCZNk3X2R71v+aFIQ9B
resYyTF+MwjQ/03PJYQaw90eCYWHiyhT3ypVGId3ZUhCbH9P0CJUCAJJ1c54NEdS
MTcEcBMPecRS2n/2msHqrf3apfxWHBXSctN2Kd7zcn1rE/bOLEbY9LcoWgo6iVmw
3CjTCR3w3zrFxk8xX5ZXGgcZeyN//i3rq3fiIH+gFCaWsPniADrGTq9080IR5xY0
gu4f1CsAzsPBamZl3s9uIBOu2zqfih52t25B4hC/NMlEP5xT93Gm7zPLKa0QIaAP
IXE25bmwi/L8k0N6930b7Pm6vtws1otDCwIWZMoD7WcdeIPH8ul3wJyKv24sqQVZ
hoTHeof1Dc0H28tvFLpLXxTNCWK4hRJLLFXTyXfzvcYlfhcHCBtT2P7xBWAQZCs4
3hBkH3Z/viTSMF5E2aKxja6rfO5rvoiYt296FfU0GRbQT51DlS9+ENY5nYKLnjsF
W2B4rCt5RvrGCJahhV1S29eKvmCZ2c6alNTt0iSXiqf4VCOt5TmhXYXyP1mbHCEf
6pjch1l2tFOfoyFiZumDNtjWfJiAl1Q8C3L98JrQTEHhKpGNFfW4pDd0JbdHHjVh
+rMMu+k4tOyDikrsaeLlUshaiw2e3XD+yubr0nYjWhKQE912m9sfltT5S6Cs1cSR
y83XCdV2CqflQNN8tQ3hQR0IZLc6LvnHQYQb12klF3meAqxyWOVfK0y25cmbldx3
v56/pHqhETL4NFzhSIyGvJKShF4+3EyZP4EO5fVKRF1cjuDMwjBMjLqa+47w3uG6
Uc/GSjZs75uQnmPsikIxbitNZljiz62R749fZJgZRX1pLcyUubdW5YpeGIUggKgr
3NJZAP8T7sBhF1UMdrLLmhJBBAKoyKtYKWfzaKv8oxfon4mIOtIJhhkF/5qikNXl
zpJh2vIu6BZXEI1fZDrOG/r2TFNKPzOnh1D4L/XtNeaDLQyKcUDgAopdpqrJ6xeu
cmpB3nRP9x77MUoanF2Ip2D9GmmvEqAnu4PB4jMfetxhSju4kXeDHQZEwukTaBGV
04H9A1ecN8ZAoibYk/LEyjXX4IVGmvZlJRspK9sUxgO4CT3cd96uLO8PYx9Zv31T
f6KI76BWTcfWS3wP5+gpYVhL7KyCjS8fsI156e1PNuIwsaDQlEXdNbWmb2QNwiuL
E3MsUJu+9uRxzND23X1LPYW94+3dHZfPl2/vrBQsmWv3QtuCJxK+aL5ow7Jyb35C
U91JpONAV+dOkC5+gf9LVrTL0rzz6T0jHWWoWJ0YKCSPEQidgsldBfcphE8jm+tm
KU8k6RFkYlFj1smHbXKL+YFJ/HIJMTZqHnLT3XGBs7QJfND2SeSzpUuzZDt6bz/x
C/PRDd/CPa3fOqKJrWPLZEKqt4ZW936Asdy0gxfj2OSHmwit8IKbZtHpVJw7RtlL
4gQoupReieTE0F1o+Qz2VHhsNTuqQJ4TAhdv283QZN2535kLxbL6vTRKykW1Fuzu
CvKd1pmgdFs7K7OGn4L5FgMEBw2PlPIgJ8uOFGViXn2aUteT78BM3T/yMTbNmoCb
aMnnQzn0RfYyAySm/zeBvvoBO3CwFYfFg91Sg9XvnZVpf8OWAQVxSTDtCp8kl3yt
n6kgoMbFzieTNaBnq/5qwd2WH/PosI9YEIc8BrLGTbyN72knf4JAZwmavhADSgn3
foiCSnfg4dTq5D99vZ+m1kvusxm1YI1lgQXQ0rByLHhRoOGUaVZVJ2mwEHjn6AbQ
Al1J/qI+5AKqBqfQZ1r1EXzHlav9bVgy/6XBqnc1W4vZX5NwmALhXVm5Cai7cAjD
aQSc1gFHgrvtRXAkla4k2/RNrVtAU1v069oGhDmmwq9fSXhGvGnblIBYHMaS+oms
mgr3tFgkLazAl2PW35r4KhYmBwAlqk/oCsHGthARN2rx7bsB/9OjSkayoad5AnQN
PLjR8wuz/QXeFGHwh4jkdgkEMASOi9nsAEgtUcDLcMr9/dAhXBpJ5aBsrCSVadoZ
NZ2AEJNxfVMRN91b5AZk4SAAlBxxLaJ08MRLZEOSLthgSpyCEuJW8FIAyso2Rt09
em5dXOrF2iSuAy5iUMqmbOwkvKAsAamGiaQnYwqLXx3W7PJ75f7shcxrOLuX5vjw
LhhwwoSWYbYx9q/Tim8i3P6cIGbr3RVqNEDkdGn6jGa7eN1bFzR1H33Ps8A4oclV
zTpY84ZBr4HW6SPffcP2ovkPUkn6A8EQdMmRRYR4mzPpKMqAuwsXpKI/klojhPnE
f/0FquPRJpGJvTO3p5DGCDVXP7iScqCQ3zAkYdnsy3fG4BjgSV67YMwoYX62Xh7u
R6Jot/aB5GmfK+9E9Qq2TeNHE0gMtKasCkR+E9w3PmYmjoJeSP9BA7ZUjekGpNGJ
emvmOSNYIGoCGE9OcoFJuGG58vcDPGJVh+m2awekyb7ni766n2Nk3fjLFM/hNJOd
khtSPa2MfuUln14RnwumP6DaOesLekwGpEa3OtQQAWKQ1NPFkk69TTej+OxqGhFF
fDXIDZDeaXa2UtjaQbHAfzdu1unwK4DqELP4DOfZ0nGBamfU1OPdbjTk3lQdHgHy
NR0ysJ8eSvLedmyDd5QI3F+snyHV4L8+3bBT6cpbLfBuslvmSPhxlEEU5D3e7keL
vmyVmnybfCe+kXf1IbwH3DExnDNbGf+HKw6kpY5tk630TAPni6eINHqSbSa9UwZK
u+lmzb9pml7YiHOaKkzZsaO74M8IZ0trpick5JaPdBR5zMvy5Tv6tfHxeVlt5Hal
DNgFfbstgVZUcztK2jnAoEAUfwFP0H+pteQqDyCoW/cCz0WIl+DhYKwiHYwOUM1+
8NTUrVba0GiMFfSWzqOlHCxVIzPUKiv5upETO9ylclMn6JQ5+JDUXAcSZ2eR4ZUZ
srMpGqa8rE7c/2rWzlAthrIMgR5n0vrkXdNyz7Fola/SdSI+U9LTmrbs0Id6WeBb
BhmK/Xj87Kg0Yf3Bhx48jHv008q2PPwQ/SdcpqHmn4SsBmhfqA1z+rYOxMqJJPHu
lS7KyEw5ieYtvK6yOKDMuc7D87dssPceF88rhwfM/BfJDdS7wB1S+ezB9Dl6vszh
8x0/qsz2UBCWdIfMbdULPr07lQXCAylbANJujda0BaXSljOJ+iEyGiB2TcWpgJrl
obqmUrVZODg41+ed9XpNWX3NjfCUu3WAUWnlvwRb1q//pP2wa+U08cqk0oh5KyKX
vfjDRbU4Viop/j36GVwFezK0m16mpISsabj/xLso26HiWnOXoAtjIGnI/JZcZxCp
KqLNnEIGJJfTOLdXlM89bd4oYgEu9sYffibGe4NLkPTNqaPEV5yvGG9nYRygjpLb
L+MKiLtBWQEYKeSLzdSD55oe/wE9BYXeTU+m1IreLAyj+Yfy+SIQDoNzSZKaJRh7
LSrixYvx2mbmojGEr/vecwZ30xUfVc5pGQjXSk9e8SMxpBRTqxWenvCAASnol6nh
o6KVse3SY0puwqPE9Q+L6/ElkhazqIOrhXoqlxjpoaBnpEwivi3UIQP5WvmW5HPN
Esk75cB4bHbdtLM8zMXjeJ+WJjLPbpQboOW7qpMXh+Ehh1Kt1rOH9tR5QHe/BoCb
6N8S7rZy2PofXeuFzkz0BLWeZ4bh1ZCZRhFdKWsi4Rj23GQUQxPnIF/LtFCZMfhF
dsnO13h2oBgduXuLoYJaYzsmCX2NerJ47yNYoKTe6+3O3QVwMcJeqWIpj37mGH7s
voJ/kXRecDK6k4cUEg9Z7sb/Nkt8GlO+z1DCj/pI4SPcGbzVs4TbraUgrfQvDT3q
sZzgpLGopRq37Z6TQieQFY7LKePk8eO36REm9gv7BtaSdghWj8/cWlYcwW+KKb1U
M4EdTrYnmr7DzTaL5gWt6xCHKKJcBzx2xE1cv0lIrsUmWarshBhCf68EHudZuROV
HEnoVeJfLpbVWsbYv6hTK4xTCmGI3sGI6LW3AlJ3nmzN6nion4qiiOdMVakecY6M
VQIsobF+x5jqwF/mcAGKW5vP6LiZCgeCwrK9OiPKrTD/8XSYtHc8pT3M7gvcTu24
nIhI9PQ1vpWq6XRdNDmJb43resmo1rhI23Vfpt3tj/t9jqNgDASektXVJRGDrSP1
PoLCe7leAoA37ScbVGLXU5LG3ly9259/ajlRoWRQvdXYI6Yr6aXfKNJa622hDEdm
uhGrIqgZjqhrPcU76wsAuOE7bXdGfmdWdZZPtzV8sSo/RbJrisdHea+Wx9P8zixF
958Nd8yiIO3hpriX4fKGXH18Y08txufSfauOMCzbLlhBnfRbDoysM/eCroOj3SEg
u7piL+S0UH5jDXP1ygeNV7YrTu204iE1GzGXInVAYpUefv1SU9TzDl9vDYGlHl6c
Kra/KNYgsSN23xaD3kfD1Lzj3L+pMRjHGG3Oc+iaKEuNBFnJqdVVo4NExtM8v44o
dzON/ZK1PhWoT3z7UnTBbjbTFlGL+0J+rbUETcAJ9hr2RwKQfXX0tYjrTQ42wsPH
MNozDjZRhhW5vmi7ATtfOOSZs9jMxRYhxRla2fVhe0Ft+XdfNZXJfOFuFXqFIYbZ
lNlD5qmVn7BN8MeWsKR0JJXPDIBA9H3sj/xvSfxEum2IJXMnT2Aj7406g+DbT/7f
VsLpHAXcCoWJdwxvG6S2ESc5tvdFN4v7LbsaNwaXtJoqe3q1VHhL6AmKa2tCvHM0
+RmMyr+yG7gHMeVysF6OhaWZP/zjXla08LFVBcSq+isBnTgkZmnCpwViP9Ks314y
WrHmRf2gBSNsonrR6lJL9yRVXtWy6c3Ev1O2Ceub+41mEPG9Ee/jR26eHFHb+e/k
cKJK2jLd+jV2s30nT7Qkoq03t8QOMV2awCccfhItQ6eTx/SFDDsxLlON55295MIJ
d7k3OWuy1O362equW+dL5kkLPUh3i302G4pIK7EZVCVVN8sQ+dr8XjEFAC/fuIQt
2+k9DXkR2/WmJCO9bAILlkyjbKE8Wxp1begpJpOMLkxByjobsehORONmxQJfQ/6q
EkTr23Gfr/IoLUrCj9IiaRRSrB5Os/rKM5UH3KIT20az4or/Wzmp4F4sbo9+NbIN
ZlglE9XBow4nEm9FeM5z8j/spLU02jCNBNJhp72v32KPvrc1fwIo7LjI6FQj6R96
rlx0F/1W13Gjq8HNxOIPNnNXRgm3y1vnZ3GWzRy3WzvT0UPCiPpQUzgmwm8T0lmY
2sUZ5hAZrImMZrI9tlMVRgjXs/WkOogkl6o4NMyZA9LUr+l8ryyXOlzB88LRRWdf
wIzIagAOGN+gXI0MjdLQASzZOu/MPGVAuyeUkIrS2V96K2m+rsL1Cvc43mb1j4TF
hkvIrY9II37bc1G0tgLRsLNSJwnKNZ/HmVpZzg/6QeTs1D59jnYbqKAAtIiItOO8
9CB3A7ENAOAziAU646HH8+6SgpuENx+c66Bt6V9//P8AQlBSus04UEL+4yxkWG2+
jpkV6lxJmLwfT6+ZJk7NS6gljlbS90xDWLGuaBrU0bzy8HpG9a48Baa8l0F4YzEl
EG16ls8e3HLbyiNjuXfd5BQ5phFGyYcAe1DYTo3jEAHID6zoK5BHoXucJEPIXgjf
0QI1wCHELXh6wK1zO9ZugSMefEFTp/Y5t1ySJWrqbxMROR9tar/TE4lQG65LcqPi
TO2cChEijrqOz/CHv2m44MOpajsM+9GVjh17bo3mNCxcPuP5yKi2NmqUvhko4diw
43WzhOLavCMplgtZrSVaZflgMCAvzb/FH95tYYrERujkstxvOnjSuT/nR34YDPPe
eZOL2czaLtLyr6rFO1zm3p8+9bzsHPrsnWJb+0IAj9fgtlnL3LXZVe6hrUsCoZvT
+sBgAO9cWF0LYKLTqlWV19OuXIroGDuFLvDawRs8wupuITDNv4L0NcRmfk5vQttY
KD+ZnST2BdtSJqk2McN5XYt86k11O/WePY9pyHpYAfM7/EZ66+zluzeaa5JRF5VC
+dxeyw/kBMoBIzBiy5k6Wlahe0wy/mJhh6Ai/GkZukEaQh6hGL5WyobdfA7AACAF
Gx3Bj7myZKqdNuiw/KhP309GnyjBwDOD8ja7pQ/v7dg4uo76bsQt8niNngip+tM7
+cW7kzEe0Zb0XuUHo2F6f7oBkSXCBLd+QewPoQTOLL6cqWEUbmDZuJq1gM5oNsoD
fiEnfg+MIJnYLzZ10ivI0+uG1eqOCOSEQ7VE+u+SFIakVE79ECDsYNmbC+kbdkiy
pJBWAXoaR3VxVPgsiVrMvC0fMWNF0hLVdmdW78SZ/2tOPM4AG0DrcGuN8cFu1HD8
xqgU/itKeYvC0CvqXv6voQUp204hjdoZONRpOXDShCgzBw10J3g2WjOBviHXw7L/
/FBDj64MH3thaAU/vyR4toA1udXgLyZVJq3SGf6Uwcxf1PXgo43xGlybM3igS+bP
LO5/XdLUEH+BSeXpIz6k4wtA9ByWib00Zfc7msia4Q8N0sFE5dvZ77RPIOu9kAjo
4Ji4E2HOxAn7qZ+dO4fhNGJdre7qsBSx2xAFKYlCReL5VeZmCG/Kok/3efoGQ041
hnewhNlG5Xr6/L1OEq0KZac1P1c7rkZXtvTupvmmOg87G2wC0ICyHz2aUTo7qhzF
BlgSZucdq6DlXeqWPskTOO49AYygMULoBDEvvaBcEjWZ8hm90xgv24cVWBU/8Ht9
iS+OaEBwQZ+bbjsFtBe5YC01V592s48NAnsF7dnD56I6CUQjHNuV1gdHgmjPc8T8
gjIM5kkaoaiVM5EMjjsDUrYjz+8SXIaJOvphVX/Er+OB6W5k4hi8H/xOMuawal0o
6ROa+SSygIbex04ymYApnAqJ709ktdjQ/vAxxY4m20oTRqwHKgTNRL8C8d3Lgz+p
Aqqp94qfYN1zRybR+RENml1MpackiEHfTvcewpQ36DSvNDU715uYhn4Lr+I8gDZW
7S0Sft5tcEZGo0uyjlAvsGs7sbkv4+NW2NQFehQ5ZBDRfyKNkPhQ4abhbenvhr/X
R+hQPThAML+I04jevbinkgJWxYHOaP12y5sChrKbaKMqzHP6EOOUmueQDeRGvTcy
OaMSFe4M6QEfXwjMtGmzIKGXXIogbXJp0EKhrV5C2ksMzdx3KMc4nLW/NobG5mVR
QoLGB//mFd7BXlra9hdwa/6X8oJfVz9bZahlHv6Lk3wIexeUSNWaoW9aAAVbV9Ui
79BUrYVvieC0Ygm1xoVc7qpOXBpxZstHLaH+9u/NlTXffRAZBLcKdavMY4ysAOOd
PKqlgDMGWYBy8VuaMAFWRiEWv8jZV3o7EFZFqArDNtytvP1jHJKivL1vEADDLtYK
l5SKR0PTnXJrWoaiLOT7Jxov2HoQ15pDAfTsjfXbi2iDbpet8VxWO/xBfK7Pcho1
3khqWyJw4/L+i07gc64ZUkaFwY1dq7ANqOFgE+QSvsXQyqu8MHVYlkcodnSFUhkn
U+pp8Hu8TP2R0328E+RKFJuBJ4TAK2boMVD0wZMTg9l4oxKqTbTO+l4qBBLa7JOE
yz08ktFnzXm+KbJiLIT24WnuY/aWn8HWAiJgV55O1rasVRYzzO0SK6/hsrnS6gv3
s1vpLxX8TOqjcOHJCqI5BWpRb9j0p3w2X7hdIDzD2WKwqwyDn+I2fQeMdMhU2RZg
ioR3sZ6y46e4vDxTx5qOTOAZFml+Ckb0JRsE1iORB4294Q29Y7mANI7W3qPdc53k
D4qFcGbzPEYFFhPU0G1996MOd+XxZTPbuL/ZRcBMO1+mi40DceJIlkWzNDhwT+qY
+EOUwHZVJV1E+YBoru92zkDyjyl+QcPZ84QBt6vJl5mK1grGA7jrjmv4LiKb9muf
B8KeP2+ZLeK0m9djhSGw9MZMhQkhbBHFS195VYuKn2PLtkfHFAMykClSjFxjqa/d
kP+XiOmmisM13+bzLgtjwHWhCNoCBiHr6reMZTV7Ji8pYwKm6Ol3EdxYr5t8EcvS
wzbmZdM4ELFUs7RfItReLGkESLyNFzdmoTmwiILXFeZZdQd91BdVPdd7G0a8yOCb
zm/X3fHShysTUYOmjOLQ3OiXRwdidbuSxxKPATDMjnAqoeJTuBSbMESa9CKyFIXi
H4CP0tVaOE6gQaJk0ovtwJmC2WI6U2RRMPz5I4s8zl7YuUcdLxIixsw6KloGhIVj
MGJLg5n6ek9/QHH60haPJZXHo6piTI7TQB2+Z7lsk29SRYvPk90uLOpz72IMEzik
bID/Z55L36jNe955lRkoRFOYEOm1N5E70eiQcheQTplDvOHsh4HDpwXtx92YeH89
DmDkv2WZBSO1HUEL/njwF+3jAA5hIJE5NFtjnyDVIX3zwT0lKnkg9XYGR5qgU36a
BCCGyyC+e8TpOB+0KEuXgCLZdHgxIg61znMICfPN6/X+KlLryn7C7bWYnJv0QIXK
4c91Hvs8D1eVgfogFyQXXVqYXRl/3iql4V4XHNBtK18izV3x6lpsLj2WPHf8oUPV
Z8lQh+9AKpliCoLyBC2ANQhFBbzw0kkaiA2wzBT+Z+x/gV9X/Gi35dFAIYMzAn+d
6vvF609AXjEcofonl7KJteLJXInoM5a9c97CdPWnG1SUv5PVXld66phVE1xcKO9f
VTLz62Cz1sI3Ziu6qQKeu0VI584lDzJBnnYXb2BPztFFPANCMDNTYX9SlDPbGnpF
tcdfkS257p0e32W9b7Fp7d/s6zia2GyvGItaE+OfGfBiYr+v9GJkYj0dKLJiaV9V
n6yCogx4k7k1mOhfpOamh+N6PAQwMNQIJ/i4B55FD/Dz3IzjCVpPlPuHYAXOua+i
4O4WtVeXRGRzNJEVmW4GGhZlnxYRh5GbXltvg3ouFROKtPHXKk6r99mao6dTD5nV
0lEWuOPsoDjWoMuI0mgRz8CQMNWCceccVJ/Xud4IOwpI30/0VidTbD4H9FuC/BpF
bxTzdLFPIAMIGBVRE7KYD5Bn1THx3Kyt8UlKc3DzeA+3aHfgEXvpqNJOr9pRWIrR
PdBu7l9W+eIA6nuop+3M3d9eJnSXT4cqOBkytqnn8Mye+ilJwJpjiyaRh6/P+pkH
FMN1MkSRcouksTaYphP/TqSwqvrRhzq5GIVYK8CmgfrQKXhh9TgAsRAVznjyDmF/
ikxT2Qyl5NpashtuWOrASIoass4ovzcf+FpZp4XiP+5ryMn7PcmB6Z/fZzzwPDqO
ltUwld8H7ye9gjBmGqArSZQu7I1jf+8h/8vke6Arsm+N6+6JJzIYqGzgP0Mzk1Az
6gkdVWInOqk/oO428zM2O4QnmKLGMxl5HbINLz6uEQdUpbXxICf+sThANmlhMnly
vvlgq0/UTtZxll/6h+iaxLK1d/H+hE8HhaFK1OawL7ZNffj7OJ+YyvfE/DknfHoJ
1p3TIQ4qFZeQbScp72WH57ecZ/43wUApcCKIUba1bXZfVy+1NumuoY+eruH1trFw
05zNUaQaaiCqBxgbwM+9ashk9O0+TYfmU8ri1ZJINTDjGSypl3Ulxfnvx6mICfoz
Yk8DcCOkUN1fs6DSF5zvPXxEncNc6dUcbpnuJ92nI8H2YrbXkNFDMUoisXJoqtxW
6jPzHxcNPYPlz5TrKf3ZNzEQzzqWq5pbsSxGZt1BVXoyk6YgGHdpa2N5DerzvrH6
N2VTXnPpGJTGqaXVfnzfILbozs68CROS75FezxCYSeg6ePGlkwqoLnaoLv45qSH0
/B4pwgx0EV4eN2fvhLxY7PzLJip3VC7y2enDxn8Q/9ssIu20fulxNok6w6/ViLEE
3amEsMxLRuLjN8eg8Xt7h0nSyRpJ+oR3OuuqxrAv63p/woZAY6E+Askw4fc3kmch
DQm+euhXUHaZMdkex9PYSpDL+b/dLXMHuGZYLt+N044q6OkGuJ5CtfJrYj2rqcmH
4HcWN9PPlynv8g+QXVW0RqGtNR8lfTEqV3iVcMESCHhHx14rDLddd8YdhApdLxhq
UmLPTiDFILoKh3/CnwKE9IdBk2eTQlHHtHigmoMgA5aSDZj/MUWFmaZaPpiLUZPM
0BDbTs7oIlI6WeOPvkwOIpxQ6cuK/sRKY3oKmOM92y96JkkqyK6qD6g1Cy972Ay3
1WOfL7olzjvr/v3VN0i/IVYfsj+mMzORRf3b5hJJ16UJxU+YMFFCTpRx6JmYWOdb
kmlslt4nuwbwaeJztIBD5dyn5LvCYGMbm89lEjVA+Fz3KZAYUJVtuio4b3I+tdbc
7jZU819pcPgcpEz1wRRFpchNpST2xzZhOcRsLTw0a84p+TzBnqSlD2QsXD3Bg64m
0LdqmgU/PS7bFB3zAkyia9q+T3R4WjG4NJNVR4EqWAMyFHSZNaD+GjutcNMNqdYF
oA+FaL0DEXzd3G0NXgadsBxfRlsOjdTUd7OMcm9ro5PhLIhzRC0RCgvZOL+rVaWu
rFIK5YVmjVTeRpAAN9qmoasr3tjLIB+OdJ27QSkim9UkAZeQkHAkIulzn0p0MqSG
ipTR1pXbJoSxGFdtJfoy37IRsks6SJQbXESavHu76N8MtAb+QfzDMhCrryt0pP7c
QpPInj5G3QnGGTZNrya8zIvVjpuZCf6jGkzyg0JFzSmaIc7nfxd//JKCcL878tGp
XSWbHe1ykQ6WBrOLjhENlQYI8kNbaedt/JKo0b9svxfX7r/2ktlQmCkuvSvyyG8R
tJqpukes+zyiVOw7/uvojOdITs+fJgrn48zYswDsyBTBebmS9XxB8Fp3mXjENodg
j0TyoIRZR0GrTRBPLaymGgrZh+2BX7PIG0N58VxnkZ9insHri43pS8ONF5zigv+o
VlHCh2Tw3HDxCNauw6pk7mKuApQLgrWYNj88QzXy6pBD8AsciNVr55P8m1vr8bxn
yEOhA7XZmqKDqL6OBRs37fr8QtFullW60jIanxxVpqWPwFMLiNEAabO4e4LXtB1j
mI0wGRefteqoqFKOvtJCJa8m2lsM4zJOUAJD5LI2H20Mv3AyAApoaYTXYQcQ5ZBy
RwJ/GSwCmAFsArvfXQB0cNOQUiO3/ern6oNnuWBB9hk1bhg4cO+pKBp8rbcdp79E
pViCFWIbdTULPW1VUTqRmn+xW93gwshPLtef5hDmaUK1Ofptv7Fba8UPA+YZfPod
9VA338Wmpn10kEtAqWLlTMxy+oc+pY+00oE78wbYZDPrdogvESIT4Fhimbfj3/JU
zIIuYm3BHjQA8R185Yfkm1eBDus5GQei3WPh2uJ/vv/XWSocTYIjgDJJTlxJVnqK
oN3e9nDx28Jyca96xNFpqOjfkNKiD1u4ob8LIAyfhqaEZcY0rw2VGCI4Qde7O7zQ
+eeWvzKkzvL0Pdg/AfYfm7TgbkimgZ0s0VSMnRj0mNQMRrx/4fdwGszqksJggbaY
1AzXQ56X2l+lOzeEd/r1i8wK1+EEfmdxqMLVWzcy149otd4ASaeZurfeBmSj/kkS
PPbJxoafY6szci2xinfXXHZ6VlFjs/rRnUCBh8v4MghEx4n5rvUdyb8IChtKIGB7
pdAzoqPGOszvumS8o1YrcNFNtehMc02fiAmuJYOLvnGnBXX7pzhh1vuHeRQizCCF
LKsSW1tx0LRkN4/iAl53XqSvIpWu0Gke2UoRnyZinfneoUTgWqCxS81x5vbxQOXB
oz1Cb9Ra+8yYx86/WPsrAt6hTcYsu00Fm2RJK+lLSIcO40T+tbluV93q7UF7ScyF
UTGYMRV9hVi9rQerM+amPtbQP5PSIHjF3lk0BD3fg1Gst3CwEE+gWfIWLpQ/0AsH
Fq35uFfuBBEsscBI83jEegqNPowR5Yu+vzfeXp85cZN+6Kj1asVogcpLkEQy8i+l
1OFsTtIbIzc/ijWY1eCxu6bf3I3jVxHBcLRO1jVoW9v/yNHZP8k8HlW9G2clMe2h
T3sG6XUBIkPWi5aLqguflxD4jVbFq3+JK5gTyk2h8wXHOG/KsjKTmAnj+7QIphyd
ewUQwKn7rqJXAZluZ9d57Ds3pxJnf7gImYRKGLLXCUtC6laerVkTkdBFzk/F/3nP
naGvucqniRCQVVK72Dd77fAPQGKhy7McY55y5JtaEj0UeX84ovoafS5mRdJ4kXlq
HdHEmMzQ9cSkUeSiWywlZMtlxmQTpBpI7vBWRlBbpCFQFE/w4kxAbFMqiQDOnWxJ
Q0UAc7htq0PrNXD97dc3YB7FI3k5oT21EiYS3HErqX2nrDIfl77ChrA+Jks/F8qa
NQcoLnxbrg7Ra+vZtPIW83eHvZT2zjeP2bYGxcKr/F4kXsjJqG0UQcXB4nqicdCp
0LBLaWIgRghrMEC6l0iOQ1Yl0KGxRrGcvRsBEyail4rS4tGfxginugSLc9EcwW6W
yPbpflGlbq1AfEcol0xKYZ6qqJLdUL3dXWTFejWEbtBSLu/Lvz9c+Xb75eSz3CYs
60halWuhAtOC2oD8QlNX9E27VpSpxV7G5MSaLlqwtI4oexLnflKbE7F5AT4hOjQM
qp9OOec7mgaVtSyHppj/7bCmQF67E0w6sF/ARKMKifkDqalE7u9SDp63ybNqM4t9
aTIJXwMkGeumMfFxrbjeBfawdkCats0+LokEwMwaTnqufUOlEcXFKEkBpquh1yx1
66GfC15FXSJypORDKtTtjF/Xyuoo/8h4N7oxfwb5IhHQc8JP5D3jZDimw+jFhfEQ
L1fMFbmeelwBUtFuJEaviIVIGUmpb+OnH8U86WIv2BCV0j3Km57XUW6D/vbvbvg8
AVwMbAX/PpxukkSO0WEQ5EtdlKOeMPg+2RKCKxf8TL9OvcuJm0I6w3mX7vTjAdsu
zGh3PmBnjNPw6LCSSzvK7KTeUdw6H5z7fMB7sK7clEQaDIMhaQMM+yAzhhhZC61p
Ny4/jnPFNhFXkHANyXpGnSTYuphej+Ub1HKDP+e+QPiLRNfHpEtuTBzzwwHb2rQf
fbdoEht6RI6D6hh+W3+9ulxh5yRYhyxrU3GE3Md9JFYgjrdP12VME2zkUocwo3F5
H3uvMdaxfMcnSpmdLr+6rJssVdjsnuVau80RQU1jdvfGhZjAdyr3Y3isKCzMmY1R
/WWUW8v1cfk5yTkWxon+yq85SBVMcwYZbzX3XMDOqS3Ki+p2zQQdMO+73IIPgdBj
AAuhij2b474nswuGJR+XA6tqluiU8hX3p1xDMu1x8jH+L/TNXjNuRQWCAYlvWYw6
GsBeZX997F0MiN7YCJbhGwUBJEDEArdeYn9odzn/LHE4rgcHq1/IAtPDWwsXnEz6
qAehYJyyt+XplAwfZIZaWEy+i5vgzJhHZ81ZK9iFcsj1w0m5tcrD/PNM4eE2v+y+
pdKCBP8Yh3ohzJ4jTtNLnboGGpp2l+T1GwgusirLq5PNJ8gtNYIXKeISulVPfbaP
F5AY6R0JZTvoOcorCGRe6jhUrRGj6oRLhIJwus/fseOtlnN0h16BERb3th1gDx+z
Ze8JGi9ZNCJwCbh1aIHaNfVX9engh7AOmqSFtf/NpjanAwGt6qoXb6dk3c32oBRQ
Qi7QFq7ijD1BDSFFlp/4yzKhhtVKfWhxRZG/cJQaBJ1daFWCsLhjT9Wy+izn0k/J
vSl3ANokDpsA9Xw3ggnzjtmhlbnu4J0qfHVQPw8tV8meygRHsIek3FrVYM43IaDF
c1eqWEaBGAWgFNcAv0KmffhDXIxM5ePlNQUSkZcqGCLM0WLVMiB6yeCkZCs9UL45
N7Nd3oHjfEv6uYcJ8X9YNK6bIeWV+yE3OYDa3GMRZsbcW1Ocl5V6eLO5WXMBicAw
f5qEZbELhseu8GFiu1CfucSNPqy6i9dExZvRb3dxYqk0pJWcdUSWhJDE4GM1sZnJ
vtax/qFfQ4/dmXKCMV0ySeCgtDPYHWWe9omTa86SJqXhWFtnOM1zxr2xgWHGOHwx
NsHouNYBbx0uNGz8KRPD9ZwuowwxmOGMlYC6OfT1/B4InRd+sCyK+G4HNZIzUoRH
uVbzTxEi/Bg+WgFpExWsLZ1o16Rj3dl6xDNTmDPrHGg42Aydtt3PZo7D34f0E39w
kqiq3o9LTZ+IZNoFS2CWPJFLSKjlgaxjKXJekOfXncY0Uw+rAKAGMKmuOwq38E2E
0zv4cI3J2gQcb8HzhDunOuForliWxmxRqmk2B31Zf0Ow72yrY8ypCYdAlLgukkVd
jAx3fnIUN7cG6J+SBtYLLLP7KXAKfygpuLNu1lcRddjYxJboIuL3QFoQWODggLKp
M5YIlh0AOBUYYVN2WOzs1ISBFxDrkXFi4E4b6sUCzFGqv71NQ2eBANe71UUN6XMl
MAw8gWsgH+gQjQ+T3F7XrMCb8Dgnw0B3gXjpxcdfad0UKBb9UwvNCOZhd8W61iNC
rZAYXztLoI2qIzOlITs917LrIJT9b8T4pgswgL3Nk5YSaetb4fwtq0pcpAdEUvUo
VhaSvAdsqdAl9rdIt0A0vW3yWQoWzSBKfSPYG7JbJYMovF5sXTrTA48qOPa/Ha6R
nOwfsFk8s7OjJRLFm9bY2c8GuXj1MuqNMPbhe2G0oixdeMYdsnY8dB5A1LTG/KkQ
Ho0U8EhAWjM1vJlpnkAuo7TXdLFHcsQHsMJxrguLwn+DraHmcZcmoib311zuwK3b
ZzOjkdE2sZTURutx2bPwIihiWtKg+viejxTpRqPI9gKwIPG37276pc5eGephV9qQ
tXJYn+vFgr4dmV/U3VRTO/haldjWPCinxxttAi8moJ2uSeS/1irdb17nmPILwKR/
aML+NqmVKHTUF1aKugU+lhSkA72pbm4tSDGqJ0a6zVoeDgdLLwkSZh3DRfbNQfnM
c7JZeOvF1QVfXtnmuGcNKj5zQ2bQF6vTG6VkrkpAyYRmNHFCDTNGOvBcn3JfQ23B
06Ad3O52a+dv6d/IOQxLsa/uy8//QnLwO+yClxn8/9J/8k4Yg36ErO+T5bmwACb3
vUXs4zAh+NmdoF5FbIS/GkWD1Jgcljo+fUTeAIg2ijIMTwZHWWWM9Km4pRb7+eBP
0yNiPF2iwv6mbk5Vm8RM9QKHAk1bYyoHKm6Ta+C/RLE45qS6jlp3dyYzEwfjEujb
u0CLi2fLwb7sbUyAaBhYjVkWfGYAo9HR2g7Ir3uUrXDUBkfU3V//cdqv/T6wqqsb
5RSEW4KKjj8MBiRWM7y7y7pX0lrpP39CXtiW0s8sWFljoWfy7Qz3KisetdJqi6rc
rr4W7GH+wemhPxfqtRHwG4OtBaFuwsh6C/21nKAsMxo3O+tnxDhcDXNOFozAGQFR
Z3XbRmxLRjZfwV81/N8rfHMLeYB/LGbFkjREPVTH8POujL2jLj/nyQ2y8fsvZkUD
o048MVScytouerZvlts/F2LdVqgSnPeEUb+OxJZlFtHa/kE0kZSKfaFxcUqlRvru
Zo1PSY4iaMUmlVm4KPLJyegQEBFOaPhRqz0zjbp3MyhgUbsF0z8bl2oBZC/iE2lw
XKkCUw7jp4s4M4xcoL8vMxLRe+Lx4JFO/VvihbNk2WYxgc8uxHBUjFuA7vlqOOsG
+vxQGM3/+IUSq0e3nnAZeuwk83e6lDX4QzPrUbQcPlKPce44S9PmqySdnwS8vhqi
QIgpJSFA5UwJrTTrFst+6fFOuJD16Vdl9IwnAJeg9KqqTnfAEQQHIW8U/k3CmWj9
ZO0OS9Vuha0qUNtdP+9vY8NK0tDICcNJkm/igDc7CebdnP59JuoqXKbFADrre4ZL
4caGFaqpQhjxlvDi/dXnYD8FZXKh9KWFT+iU3qe9DuV5qCxifZhZ30qxolGl7Eke
HchCRXI2BzRWa8IM1zsvrFjwhfffkV5ZHOxY9+aGdC1LcsS9xYElT/CmJ0vcp71E
T9VofXYTq7kBsTw5tTo7g1QM/TYZ5938ohqat2fKjI2ttO6vAYIjWVhNNcewfre/
bJKtaaR91s7xySGwUyyHwon3D90sf4lxPgwMTQP9OjfzdSLpC5dO+e/G6BkYtiBm
sXh1NOb7MFb6iNTPOkgCzPy2zTtKO886kv9ucGVTanedyJZOIFvG90oR/YA898/Q
rQ6ogC0+XJIV6PpcukEBA68a1QpXfVjwqlO7UFR0yxbrDxEElLGKBYhzwPn/vCG2
WBex8Qj2CZgRZgSrx+WUTkGxqefMiSUM6qsrp+aLvj1QPvcqiPuamiQ7yPGQFN+G
cP6os9IX3fGLkK08HQGPZ9jdcEkuLwXirzwkOINXjHHTDD4B94BKxnPUA/Vb6OWd
PPxXHLPxD6bjNqicNZ5Y+REct/sS0DeVaBEMGKapBXDx4A24nd6Wg1OM9K62kd9E
2KHKBuOySuA9Zt/GNS9JCq9dctMz7k6yuGxqct7yiK42XD8hFpYmfSYEXRfeKPz2
YKyVXVMQ0TKwcQ862dPfdgC79ju2I417VXGKUY1R89lt0M4pJSf9x7K+sDNCk8GN
Pbh9Pa2+Z/9bxbkpIuRlhyH6LOgIvrkTBttkz1MdWy5hs5FDg1zUplPfZTp+HIMz
QBbjxQSm87sipwWJtGCS0FU3xLanufMkEQq8ZOjm/vtbYSU94KRUQ6QtnZbqTAUy
Qsa+BWRD4drm/qieoWHRrwBTX2GzexlT0FhZMJIav7hfIuYSiidn9dl5o2gauPnq
CTznK8j9zH+lBNTjcXgmkX9c8qLUv3Hwkyz6fy0l88NkYu8YBdDpbdByASkOCFV4
5g4me8DoA/v3jil+tRdpW5HJfm9iBC2PxAh84dneMY7uCONHuIIGvSZD/mL/3w70
a5YCiuQcvvU5jpbI7uq8jpdQ+Gf4ZsdliRpahCxYFARL/UWaqI7oiB1hJ9nlwCPV
o+geoER8JyD/HRwnktLAN8/nqsG1e2cV2jE7vj57KHH7fDH0ihHoT29rcwvn+47J
ALIxxNweWBak04xXwKbzKWcxy72GGZpBHqWCAf+PX1eojrz+/Cz4bmRGZYGfa5fA
vLY/p8kllODVg81BBI768y0b4jST7pyxO9SLNQ8tg6GrpJMl/jDySxREoSUP3e34
togV+CFJdRpC/heRNRElpBP4ei3581IlVo8DFgczC2iJp0lKvvtuwtL4JQ2Tpg0w
QrlOuzYQKQCLHh1JGgoSRlvWkkMALOqE+PnN3HphVNpKHquvWyHm482PqlJDfsqI
8IJbZ1tnaY/TCSvot1kp0odYB8/3uVM0BXkMH3sDiQ4RPpGfLZdSvtU5QI0Z0GuD
pdqw/nG6DCPESmGv0yeC1LKe8/MtVl9EKOVuhSsuhlq3sah8F7BpGSaxmkRmfanb
qgXjmYhLHv70jTZkIGnR6R3CdkEo8B5+irqhPxGcvGiWKElPfEehKoYmoGduyw6/
S0g3QlHUj4MeXaqtPTegYzOpBj1untmtRFKgP8r9UDPKjYAC3+f9Q8nLnOiDx2eT
iEf9fnvet5vzER843adazKuSYXD/dz6Hvun7+JAJ33DjMH6wmB9gR67eH+1TTJ37
D6UU98fkL0uRotErt/gL8cSfU0Gauy+RQc8jSHk9LvTWBcbq8vuPXdko1rMmwa4C
CUwPw18urHCRSqhsHkR8PNjlcdz8I91+rGJVldjZxmwV/Fd18xq61pJdjCd+GbNr
tlqyPSRoVPynm96VRQHifvaQIJGb+TIVo9g4UkNi+U9Gshwwy0gO/EMvubn5ZOAR
qYhyc0chE9DgUT2w4qEK7VqMgzaTY9rpPovJoFkBBtAUDZjzoX+AVhJRNE5+Kcj8
6r4+6jqNMwdtzuO7hRh0KdIOQ7WiZe2BsGMI/KHTOoiWH3qK0lbET+tB9Uq2C1KN
SRd8tdlrW3krmwU7yN83zcnIwmc5LPInAaYtEMfdhUv2rGPCTx/0aQypfc28ij0t
O/yIdt3zeZQ7L2gvFZ6gZrO3tNO0+QPxKdMUMTVJU8bw6GBdh5CAaklibFL+4/zW
z+saT572uqNCEOGwnM02SRK+asfAhkJTk3JGiUV+fLfdQkGfpxlrfICov4oCkcLq
3XIWPqX/n7Xs18G7hn/i7uBmIGe1Rbz2K3/QG0fBszr2glbY17q1vLDHkVC47goE
X8eI2UqPK+7NdWcwjO9uApbzgZUFsA5pqNdxK1/VoAEx7RzRjSrJWIREGxDPc65Q
Elo6kmgYSbATMmGjshbjnGhzvkz7Dol2uKzs7xuc8RdACLMBE/1u8UtquNeFa767
s+rcMPoIDX/r42nQEkXwN5Qlbn0tHeunCiW0zqCa6Be5FCik59tfsNRPS5SgvMno
X2Sb9qgmOkTj5btNHUWD3xCzrRq4m5yXCrLPBqDF9wOocwfJXAvp2FS8X3L/a4Hi
0r76lZP1rhLAr/e/Pp0AiGPtMR/gJ/tPRv9Jmql6au/W6EL6UcSwdzZGFru4BfmS
u16wfTxIIk2aCRUf91iRnIFnj4bJuRmGjfYfNsZY20kaLKkt2axhRLMO+dMxgv8k
Xdq2u2OKwSIlvqsFmZtOew+Vv9sAI6hZ8AlRm48WATNy6/u5Ub0uIiiAMdxLo/eT
93e//SAAOqvHhrtueOq+aI5LAu7yNMsvEPh3CL1igmMCq4i2Kq9kYYkT6/7R8bKG
HU2f/1IV8MtfWgyqAiiyjRq3nt2uEMUubZAq5vd+xevOC99qpZ/yREyI4+pMKf63
Us/UJeKUVnimENWy9KSmp76aufVUiNdn1yMvWM2i4seaw5FFqXy90nkE1eej+vH+
n3gLzjXONcDYJYoM41vMOhRJfN/32kd1wyMPc4IzcHGcB+tslTvD40Cf8qSo9ELr
Afg9wmZXqaJA/s1gIWr7HtwSx3yZdiv0hpffQeacUX0qB/grWZgUKePmmf7k9QEl
D/fMcxRdcyCZ9up4J6hdt6av7G23+UmRSj5ePMuj6j2BZzw1XMQmlwAah5v5a+pM
cAFf+YOc0/+Vam1ApkRlrMi42yUWNkse+wDl1GBs+F627lx75Lri90AiyOwC5F8c
mu6clBa49mMJYYbJidu0xesAAqjyO6Wh2KC8F+0wYBlD4YMEkgKXYGw63rapgt2P
0MLkFqbMwTcpV+usbmuVeY+RKxIVDJ9X0UMFjmpfUAYW0/jAPBslVzj1zr6rjLbq
LP8xBa4SgY+lcFZlQx/YN9EAoEVq2H3LCwx9BxqUQ3fw+EL2YEmP3wbo79pm+6Po
2DwWykdPLAFzGv6Z+smnXlANK4b2ZY0RCl9+L5eS7EJYHfYKruR/L1WKJIGDJqbN
awgGGdvo58RhX8CK3ioSRE47P3kqm+Ty9MuFDHv1Zy2ixwxHbeloqJNwQJejZ7DD
ckNSNtTSke/pX9teRaKmVbrGlQv76z9bUn8hDnRpyr0U9tX+D1krLvTJKBy/0bP+
ptB0f4E5OlRwfCtCF1J2MebZYORHz6N847qtMPQyZmACGtdy2QwsFpNfXkkqhMnh
CawhOtAHPEceUj5I4lsZthY3GxkQPA0gWjFacmRuRZEsh1TviXFVChrcorlAl73P
t4k2JQcy35406VPYTiEqgmpAG6Yy6NjC4odsYH7hZzm9mLe9oYq+wlHxZolaqOT5
3lLutIxEIZb8WHFp+W1jMA3YE89cVg5l5pz3vEIjmLRSHZFUoL1IsDVjFlr2ibnw
IBYXzgfKsX6LAA1JveY5BtNe/7qHj0Goh3C5EjijwmpE2iG3F1VCfcNoGWf8xnNy
g0sJWB81hfVoSn3JAwOJvWPEFBMbz34D/LVWZMbsI2iOUCDO7/JkvkHjHqdZfR0X
14QWBC9XHSYPomlhYiT7T9FGJ6YDaKD6DDngVOjTHN2jA+bTU9dLdJGnsflTRdeT
ZIY6Ue/zI/8Raf1EQDBzLKwccpY8hRvtUD2vUoXC179zni6KTZQO5O6gEk5Hikoy
OgHXwjJx6Poq1jSlrsjnPv6da8Yw2uHTFdv70sTOnbk9tfX16FF4iZCFcHSBoDV8
3x0y1xVUSAtCgb6DjllXWC05bGr+Ov9G2EWfEHSrHTmgzFNrI+tBPhJwVSIAGrBL
XmqB094WfoZ9TzY67bKUE9QvRkW7/+l1jVDQT7x+hSUEtoypSo3VTeVJIajbPcQp
bOGJyPB1Siq9zjX8/ynI6EhxZX8y+Oh1AwzYrpdc2MHTawwxFElgGT+3AmevrlD5
Om5nsCw1J6pwvXkBrMnG+mmpZfPiHwLoshsB1/hgXUlPAU+lyYfFtHSjoGRRTwkq
Eg6NreNRFewe6H1Er4uS5rEtcRGjSO64mgPE/ytw2CS8ZEODMeQZWIONqsvClLlo
MqfSyGwQ6lzmEcNoIrCqW49hXXQa4nlTxcxoLq9uazjIIwqEwWb3gltnp2es0/IN
R/EXGjdcNgldcP6f7PVfYLlH2hacb4MfrvSmohNNegMaQ1qMRxCxp6dng3eBZ//E
ZzaSeRVtao7DQmfl6gH5T74PzyrTrqMaLHWoKhgFH4H0GODyoy3JZcyRaJVSdqp5
kzqUn2coJWfG2W8x8tuWInzuqzybYoP49SFlH81kQGH6ogqXob4jQcFwruo1xh2b
5WsJPLRk2C5qijoEBx4EaYGckYpWB3nHSgCrORK3mUovQzHF8X1N3rYSrvTUAoJR
/r/DrfxWJTBHn4kGHZVauVtdtiE8UC/rTLWkIWReBUQiEWEHqvNUylSZUyLC/ln5
94AJ2Z6Xe8voZV6/AeovAVLNJ4H6EJfww8wN3QKleC8zwvhEOZMG2zQxfC7lLEK8
zaZf+Yt3YlZdyuAktcu2wS8QvhDYr8FQ0m5VUoWCLYG5Nt2uMeCZdOvBZjOZri87
d8WK+d/1ss5JAiVT7KBCx/PKF3W9yQ17aavbWdgaqBK6G/oUjNRY8IDNw5u9xUMd
1wHXclnTtdBygl8CgUJHVmQULXud7ae90HMB40EP9IVF9LadwQyJ7mG/RqKN0DV2
NhR/u/dPgTX2R030tKPXzuNJLhmyGt2mzVFx/ScXPheCBrqUGNFMdI1oiT9sMxLI
YAXBcEalO9OtCHKLpKYtQ9uLgl8KZveKBVJBSN7HP+GF7qyde3d8QLq7rzBDumtZ
Wb1T+/kf04npT7mS69cZAwFo5HTeK0Gx/p3adiSAOav1bdwxGxFsfl7pC9R/L8Er
4GvvIUBc7Oz+O6wHwQiWBMcKGKRHCjp8rjoVho6bzBO7aJ+OCGuET/1dfveqWe+u
TXA8ii1vx2plYmWmHqkrVlzxrxShKvDkWQxMRjXb9QrLLTgxt3PA4wtCWjGk+eTp
DSiVy94DTc6ozf9gdF1NGp4pFNpbQcGGlRc8uLHT88fYGbnVAFK5S38eaHfepCWB
6th17rIyBLEgi1zsCpQXQXYVtobJzmo7RZPAb9L2mNaX/xFjfu36rCvxaJ57PPNp
QrFMnVdHZ/NjU2avSBK5lUCMrNBFDXHbI+KM+lsnkme2UPJ3UPi9slhffkDx5M9l
Bl0ApF8jg+Aa/ZnI8J3J5ee+z9UeCAqW37s+qXJO3py7ybPY1GDbtHWJxCLkw4SA
+/FOedi+Aha2lkOKt41VrsZafdLwZlB2qXhX9DFx6PE5Zr1dg5W2qcNxFEU28Rk5
Pka6bFZKBMDK1QjKqaRskB8TxC6EjANHG83JJQHUwljAUh+DbSKjzSfs8bqzKwGu
6URtTBimGe5AALuMFR1UD8FK+xjGHlHAOa9Gb4Iv+gkyuTrtrht3oezz/3Lb3hdt
iwA7l4V/8+JsV2OTsamgrKrg53vJ+C+dcjly60Z4WP2Yc3RK3xnLM2WN5QNqywc7
BVY4gSCLuX7vYuiPek47kIECBUb/OsxPgLIURtdiGhMK3L25Mo0bDTC6ryf+AjXH
nvtEhGcdh30xujhI6dqbr+0W0R9Mfc7uqs2lI+W56KVTl7EUdtRW9iLBjBOK13Rm
dCCJHEtesjhm8Izg08hiKeuoNIJ/ZgTFee097Ccc4Ez5Nh4/pwkBxpcf8Q9KSKwh
pgLqtskBe2dKHYr+3mkdj+/EC6JSqGdrJbAjGCO3GmjbPBRV3u27yACggwcz5ClN
PciY/RWFNK5QfC+jSEgAPEoUtNUyQzbDHlpBrf1OG2SVlYiugN3+m22FvB0+y6bY
Lgl24D2HtFbsLA8AxL0rQhRIPFmd9VvnrYh5sbT1bLTu4zRPGq5jgGjG5z/wjW13
azL3IthiUJrkHo8+6qrPI0mbDNkLeAW3cxQhXsSryd2dQFwJDKtu0tZvvL4QCoBJ
WApE42GS1dS92jlDfhvBHmiVI7cLgAjBFX+mB9NyxbnF8BLi5MIv3BfDu23pQ015
5Mr6GQivVjfW4vKe4oZuZBtanAUUFl3H8GfLI5rzh9Um1fCcumbj5l/21Etj8j2L
w6HdXagvzIWBgv3NmLj7daw5PJBmkd2at29Ct/LK7g6HhwUlnd8TgqMHkBYXVfTF
9o/cM+q3OWNZMfYaYC2GCWwVbBZRJthx/ejT0L3uPEQkHC92jgkNTmfwdcXBVE0r
Gb5x1uPFoQjIUNgDV/CoUwmuFomEUQy6He5a0qTMAoEhaMhzrZPdv1KO9O5HZDge
uMLc0Th0nqcwHlMhvw2bfLEzvR8YADthyXpiPBt68ZdpgFWzMGKGr3nMNCOpIx+Q
iELD5nmkKJ/x+Tnmyoy3lWOgNxj+aNDtAQU2tLNQ9gfVJrhrHyXOy51j85mhrwo4
kl07XWao3oIqofRTldj3d7ObJ2M15IpfHNXzcA+zV+UBmwqLOiVlYv6oI7W68joJ
r6GUF/aM/eP/5P1gJL8TAracdrZ9WWr+iTcso1tYfyKzqQ8YcZM1JckbkFfggqBY
kbyim3DJdTNQtIhxpZY5JEw3Cgnm0HAOIKRCY3ehvfKGjljISLdhLuAUmPNx0oQC
4Amlwre8G4ms5c/3XdGvLg7Z2oHjGStx4/tqezqzbQD22dSxW42ARabLVoxw7YdZ
MBRlBo4wWyars/PmdB2ugZSNwq+XCrkJbyfn0+w3l8zgkfjKDFcCSxAkVS0M5iGb
Z52lS76XqG6Od6Jnv5faubJT20o0UWy3CSB7FGOcLkey6CmNiPDQjAn5mOOb18FP
Ri08IfPGlye1EWBgX1U0KIjFj6+h/TtCCD5sT/j/DvuqB7qwMW8Z6AaEDOvbPIYf
1/UfsCZaAUeRK3Nle1aGn4A/lquLPun8BtA1m5D8LRkcYV8znvl67rpSVC8MB1b2
/c5AI+/HPqFSGyVGeim18bA9uOy1YXHWLyKCDrhxBRaX3SD985l3Z4j3hVTEGVdw
gSDje+lgB2Zx75eHA1pOgkEfbfZky+1+ToaQRbX/sdk1jyv+HNLxAmeibDhB8667
2sxDkg9wJcvqvZdl+mRy8ug/YBeT7FO8VF96F+529fa6sajNcml3Jw5CrpHX+mHf
AmwLDSv+03Ov/U3d4dLmI0HG+3c0qq4+aLR1K/HqLpIIGMQJ+UX2vArqktX1ey0P
8xk1yal4HWrSogy8t69DvDbovGZpSHqzLa7W2ZTolENiCpUEqjdn2arid4AK0rK9
cw2vouKxN7oHHE5VF+f4gd6WF1F39ECnMD9bgQR2/pVAJcQmrIfNFtgmOjeWRbG+
1KQIx5K5j9joSMEslvMys/Wta19gT3OY0CFrUrccLzZCOSGGJWg68bBIDO3j8ytG
wSLqoyTJg5Cj9ANBTUIXK6BXCS82NbPHDZYZzXoEK585wYLuG1w74juiiKL/dnD0
wvqJbM3kMJuYk2oWNEB5Tal4kDcAAaWqvo3oZrIRR7QyVMORyidj5HYXOFDdpXMu
bg+Aekv2+m4XteTqPW+MRDCfDIy3+rVAXSbrZdcLbToZSnkm7uFnCUEXQYDlhh+c
d54Uq5fL+B1PPxwuaAUVB4iM/HtLIAUnAqzCBpXDBexQYxMADFEHd3/LvrCNsiIC
XA4BXdSGP38ZJebAy5WoIcRxLTZc+26ett9Mzs/9fVCanH828z/gxjPaarCKcVXu
PZ/Y9/63vo5iTW89l2qRXEbtGgxcDxuALvQKGSnZaZXwWCKJr46GdPX3CPsTDJ9g
fNgkMUQo8rS+eQjG+m2DtEhyRBDBOyf9OnTeS91NuyG5H8kEVb+g4EGxmWIPyAD3
36hujn9vSo6quksULEucpIsbAPssbAH3zczJHmzGEdTy9xHjMqLy1bh11SylETpf
2u7nrNpPxdaROJB5SUoUex3QOLnW1aIuu3DRLBtQXQzd4ElEoJKXI9NQL/GDTeXx
56O/MRrYBT1lzxiYNfASKFZVEym8eur8Kg+r3Gg/UqtN98rN2KtGVXeKcMHLHdut
jdwdldbt/Xj9VKnhpfaJ+OKVzyOOO8q0ejBEIisk8bBrXFSFhyVyzgIsC5deb1Gt
2leVr49p3CEFJgDjMLhhMER/oLyqm7y42Kln5NF84/lTUI1wBF8k2ON6ChGQb9gR
VW9oqKde5tD1SvLPiLSYQ13ixllEQX1BN7MMYNLE7mDVIr8CqJlBgGN6uX8VRTLg
8UqAghTGDonCH3zih9AWdOPqXehFNgwpU+9r0HcPUXDq8fFs5pBZuJJe1B0aTbWY
Tu+hXmz5RPH1xWVbsCnGurHiCpN+pkPSyraATOFvROwmWrXJINQhmhHInKnbAPwm
dXofvRNm6V8N4lDqtbR1B1y3F5vcIUJUPd2SnlxBswbu5fIY3tTVMicbOPopcAcK
rjuycegvUT2ZbgumGtfJgRcPTM7ISCn9/AHm4aqCTCDDQEoWAY/Z0xUbPSvtoyZg
1ZEIpVknRDs4PraK4YKufh5eUcmW3TGRADQniHdbOhs3dT3GUoEItQPlmT5hSh6Z
92RVkVWdhEzMt2jA+WtVG1J26YvOZe27NGMbopP8bRmSzPrEEQ5qYcL9RQ/Bo55k
XiIW6xaJl9mVLFBJb3bdbTG0m5/R0rYJJhhwA90rMPxIfO8DIfJkX0JSyOzQxI89
xIBawhbg1iXqiR8qocN9Jvku20vZ4TgZ/T9TMTzjzYGToJxPW9OmfCE4vYnrmCGY
GurTG2yC7hJXzo9nYZ6K0YSrpJkcBjSWVzTH65xpg4HeiUkiYUUmRaBxqPKmUh9V
n9o7UIB2EaaXzQtvhs7yLhl3pXg9Qc5lKN8Hn9CiAx3GCdrVFJlrwKnSN9XxbRyt
vQ968nYuJQrXh/CXAhp+vmOGMdZw5ZTQie0GpPue0oV1qfSf63M2iyoSzY/IGhrB
1LMmhzreTn9Dt8PfOg7UJCiCAtQbXRIGeimZdBSbIZoCDt3DNFGZsdkNCtVupFPw
o98S0CPNn4CeWCb9lWHsGNyZ4t31622bJFMBdahN44Pv89a1M5Qy1eTrpffaEiKF
EnSwbfgAW8XFN+cvwwr5zGsbOrSEcCkw4eNyDfWtHUnXAjlIGrevYWG6AXQ6WSrQ
6HeX2zmBBt9Ouj9KfU+1C/b/rM/8QVVkRhhZ4h9KFP+qJ9Dtrva55O9CaJ+Z8d6z
h/u9tKH6ETxrjNcyKhqNrqlITmX5Hq+Y20879P4KiJLur89Ki3KcYRvh+fsd+LAB
FOyT8uk9+ItSdZW/f65vX3xX5bRmQMfb27Phw1+Wv8yCBZ/0596O0luoQclQ5Psg
1qwaLJfwTZbLaGmdknbvegDe2sJ8lH6Q7rxrVGeV8oTlQxw7tMhTTEN5g8sYcfxL
RHHg4HyYk6DDh0IytkN6xl04Izyli0LwHo8thGHfan4pm4XDscJ5wOcMiBPp7yZH
/mwQpGjgAAnofz/fiwS67zGx1TIty07tbuZC5frzcPDWtqlnD+/ORUP8PlJwhGjT
1lDKuGOBhUXGZAQN0jtrXB2drs18uvQtc4pTYuf7hfzT/d3woi47VAQPBi2RkyjQ
0pHjNxiqHeALDu3kKAsNUxJ1+OvDhXmo7/qLFZvxxyrt4Itqjpde0hdGTi8vvbDK
ixF7pcQtNaG6aQjn4z/hXsohzy0u6GXEuVOCnvAk+hSD0EekYS9gyhyjZswUsqau
LjMK3KKEnSqqjum/81rvWBGVIMxt6ihsmbVX41lTJoF9HPc2BF4PY1+ySsEIFXH9
OIe0spIEyoCbg7kZvL9MjvC+3XjzImZo4sXheYkBaUAPBkst+wacjSZ+oYzRlPI5
y8UDAZKyWWtxjzyAyTdr4GaAWJXWym3+C5gDX+UKWpLGHv1kQx/YvaNWFej7VcDs
d4+MWAk5Wf9zsRVQ1RLJaUnFU5h3TzXJmoFY4GrLx3A8PlzdabP64KT6DjxPWst5
AWZPOB/dplJfhshT4AIiuAIQN58/uV9mDZ/d5cgM6Dk+80ltuuq3+w/ISgsmSuxX
x0rC+VFphYtbZxw6H0KdI2XYBW9ukUGdpSyWZbBJ54Q4XZYE7UPvuy5pwznXGOjN
HKYlni8dv7Xqx4Eg2B1YF/S51zNfIc/iNt+TbFUDBjI3jSz3j2V8RLCt+8qd2XJ1
6R4aNs3MhX8i+t0KfBWJSQWk2GHSGez8SvEMeIbnndgZS/eYJKzZRVIhfkj0Vlrw
6Xvy9wMfKjh8GHkNi6jOi9oBt+O+jIlccmjEhGHhzjGm6jWWaK8OA+1py5MYBfap
6fBHkrQI1fA1sizywsCVITlyhvM7TvBqybxxp+JaVKZhLEC++OzR9p5QitJu3B5+
vYONCJ4WUl38An5lIN/BC5BL0DXImcTKt1Kbz4QPzx6mH/GMvabNeu04gsQ/j3hB
9KfrkvJYgkUihZVPTVq1w24KdvXmoz7xeyCAed7TsJnMFZAHw3Oj5a2c2hbAQNHP
l1LKuMK8nOB37DGeKmiDwFJTRCdCdGoCNGO/Sq+MVwlTj0PzsEczHjpK8yOQpe5f
NibAlLXFZFX3twrwLu/ggfhwIjgbWMloVLeKQ3DDa5RUt5+iG5eRwGRkY1G2OOc/
b0bLdRrYXauuIk/t3xDknxqgPLJs5XHiPup4iCmRVu3islzYPtxC6wpfQvDa5zDl
BUEXEV8D9twvmHmBIeiUDlFLyIgU1Z7q+rnzDrxqxVB3tp8/iXHiyiEA9SUPSzhs
OYgGaxvI3MakjdjFqQUXB+LenUa6TF58HuCnm4XTcTX4/juTuNjgd0HwhzWWKSQi
PSBt6p052PykiiLk99f2OrcpkfN3MvyCGbr6rNiNq4Hxo8HS7QorI5/eFlSoHd/U
Al2MWGWeFMACkzL7RhhYoEXju7q/gRL0gzBXSiFwExPxy5uwsyEC1555l2EEOnBp
YtI0sXds7FpgBpkpegMoB2M8XDcgLouAEjFWJI1zPORbFAtRQYZJ27fiC2Uv/Zty
IVITZO17nfqOcxTqQ7XbROyLnfMU18SH7w8+94I8U3QqxcZDO+8cRs4lQsQcuBGj
grrG74ngjYiBjqFZC0hQVGU46QY0mjhj+/DFOn0M8JrNaDbwIEDXUZKXbr6B2ENF
24uGd08pdUbXzJHNoaXlzr/NABFLhq+7eKi+hfxSvhsU5+WXKUCRLS7Shc3U44C7
uVim/xsyfo9b3gPH2SA1YYx6qmaq3rKDZkbQhC/q8nOAd3N5JTXQzVO43muZAKD2
XeyQmzO8aml+W5YYnFB72jAw1af21i3B4pb4O6sZ4DlP1pD39BwCiRj27Iep+U1K
cDMAG2MlMbKfKzcqa/Hp+W7B8zjisj/XsCN7TFBiPxaEvWePqVmHGoW9n7bEqEAY
IJ31TczcxrquFd+IcZom13DWEwt5288CIJFJCofSOUwvZ4Cbdq54P53ebN44NSWS
MMWi820M/KLbyw3RNE1ogw3J1YYmJ3g2aH2jdncfUQuk/pxYAlY/2ZI8woeYlmMw
Y/z52fojdZQ48IkY6q8o3TDtFSrZdUkscI8+oL0yABXTXvXQSlZJ00eejKilpwZh
+nPQalSISwjvOpKvRh7dKHTuovcm1IIlf4WeUJ7Lhl9/97eVPL02HW3bPxcj1WWF
myeWaMMDu3JMvPcGHJTNXKqKXqxYl5zUmanFh+1SDnLf3Ofkk5ePwORsxVscamNc
J/Um4oyFVJ5fqah5SBI4Hsj6Z2Xk9UUDOtIzPMLzz88LhlrsqORuQZE0/P1h2Slo
IUsZ/2pa7a2pSAkFXi67+Uiy26Gs+i5A8JHGK0iyRNPOModS8VxAdTV8sGZVDGKx
NenhZ9OY85W4Tjqv6gmXcSmn0iyK38pqlLaZOPHYdVnWQ4GftsLSIFf8P9rVmmSV
kgPHK5FBkmpB3YS9GXFm/89VB2FGjFjb5dJQlTAM8XbihQyAARVn1lmBPKPYj2ZI
dP06NYITRAb5oQkAL0/8DVaMN0B34PtIm0G0hu8BHf7xqnmQ5bsrphDoIlGlDUDD
IenV1RLdEj9ADyj944QiYldMyRkplLWY14+/QdW6PBRXZ0hsQ/rnR+YG8jvKoYCB
IFoxs+uQnR90ZMFYuDlb9g8rFrWMryFOl/ON69F23TySaxfwcFjwfpecu/Q4aiUt
QLGP+EnwF78ZLgho5BbmjbiIMKYGltXSCILLZzVSLLsAJ402QpDZvlnLGrlNxh9C
6cZ/lsdW8iLsKCKJJW5sK6P9AtPYbMnSAgiTSpTPr5Z1+6qnEidm8kMX8cJ1QlCN
7tHgTPMF2KKfUt2YPGC1CIfTyt81GxAyHqif5/CO4aPz1yRYvp2Wfn9hSLKik5mt
09EfigXf2f43fC93F+YV7FlJ7Zn7Q5e1c0F0ABHNEzxO8O/EEKAV5gGDsWZjVxKW
Wodvw9ztN+lhJ4ypPhir+tMJCHXDh6IM1YKs0ljau7DKaf3p2vbjWVoAsN7ergqy
RDyOkzRAlXNtH9hPFRRDa+rZJtORpkVcEDmam1iI5nypzon2iydAV4cNx5HNuB1H
PTky7KD3x2b77jbKRG26XF9UrZHEPMAJFmbgwSZiIPeH3Ml6ohVt/UWIos6fPLp0
26uVJPVrcA1Urssj5hidjq4nVYeKWLvr7OQc92cDYeNODtou2TkZlN42d3WYkZ7b
ZfxE5Vv1jq0pJwxJrA+i85uIei7mYiaAvKwiOBMSSnv1aSJ03lmop4MbPqIZ2nyj
V+LYbEESgiH28wFY1SEyWzgXQWR/noVwaGtdkOCLS00DSK9vb+nSdmH5KnPh8EqU
/4t9hp8/QSdothImmOIhrzkxEdiwdISgcfFUKqlXrkS2COS5NaZGemGHuDh5stRp
62vfWIjz50jxbXooQnKROVH101d1FWUqd3TJwzxJy/vCrRGI/fLJGEzLsJ8VKAoL
wu/5ggRW7o9TTXyj9cwQ2gAzf6M2hIQTJJaZAFDQLWi6pWN3lGwHcq1jWNk+FkLI
zcmDFZb+IQ4rxFtWAXKaxh7a1GlffY3cnXIyAjm4VuzZfkhOCeFLIAW3S3xSHFUv
ANpn2siTsvPixP0+eFgiYUogg6q4L38AuAgbAUxoRJcJrEgl1zTpkQ2KunojgI5l
hWMB4oJqVSVFaD2+tysid5BvcORRIZZMXvupnC1Z8UPKMZdBQoSczzR0sLh3yt8D
No+lodU9jzqZTOSdPncTgwX29KMdHPQr0ar7hRPjwfu6OQWmNQo1WColteTsXSMX
EEqsqpPKL2cQlX4WYBQgEK7G5aRGIrpFtkFa/blE0MRTXGf2mhzRMeT17J+xDK9U
OIjqE2dQsVQ52G7Op2Nf8+3MwNoQEj4Tdtd1lzrNCg/ySlr0J+wq91SFT2ZvVRE6
og169kYBXwC2LVGx06Eg1lngTD1j1q7BDiR87PHQrbYlT1bvbfen5JgGTIpIDRER
vTSIr6n9wr/WNaRrQe/emavEcrQ78pgaUQ7a6fZUBocIlXSVMpeZbITFSyExn7yH
CYrReEXQw/2IHHh6ofuG7Njyzh9bmZ0QJcri4IvJRjpp9CamQGoWY3+hG4TkfjYh
I+SqfpT4twnSUrvdAYiLARb7/T2ItFOqmrE34A2UuYGf8G7ejde6DFvTcPwk48OK
t7TryVKyXXOxjE/GyCD+kwn0uOsDQXtHWtdyW+2aKGqsJqwdtCXSFE3qdJMQJUBv
o6Ip2F9mwp2jN3sbwb5DeO2CHfAFU8A6EXXFTRDwU5p4FyVpq0Hm6YvMhEQ2o2cp
++aBdQxTKi0Ig6aN58aTfragC0iqHYCAZXhA/5RVnW37gnBwzezpu70fTzXn74ku
PKsmZpxr0GK5ga1cdk96QTs8VOUgzzkjULjRMUH2pmMALcpyZHOjvdxCglBT1NwM
FpDjauwBON00qZdOuZebButPBnLU1utTnbp/d+kkFHHSPj+JdY+JkmFeU3P7J5Fq
+3/q65waIQOwhmHICRE/jajEJjlHqLLMqDqg3iZHxV5cJUuMGQ7eHF0REr+vrHL9
Q4qwxL0MrLxm5lH2VvQbWjqpRsar4svHUPabga8GJNpAYp6P/2svUbQySAiZX1j1
rJ/2TRGE5SLtt2oH7hZYBPvtuOOz/bfYy5iEI4ltn+EVXF54NnFNJBbAYDufO5IU
dIA7wjOUZ29LlpFhCYv9iJ9zOTkNEGpVxGlVZSbecznBqI9ywFo+knADIRgENYFp
qWlxbaiCk2NstaQK3tR3KX3ExFiHXe3W1SWFlvpeyCFRoowVnTNmnnIP1I5Y5fUq
YVeXs8059ibwXpbr42ym2D9mpBRSaotg2NBprqSFhS/IRk0RmYdaR5CRA0ppKoS+
fxbm69Dy7zWUqhpYcRoGT48rgb+iF/1J2hYMrkb8Lrt+gyKMByM0cjDO0Kdsy2RB
r92qa1uaqLbLpRna+ChMR68vVFIIBo7Ur5ciL5fYLIxugySeOU9InyBCwEFAtZIx
J4G27238BHF2jluljDXkqtiTqraQe/onDpGfEtd/Enxw9lSyztHW4LY5cdNdcYUm
2NavjPxunKzHudv25YtRvx2hroQeP2n38YfmsZCg2mw0QYHBMM4EKi8mi8VDNXaj
k8oea3uHp3Ixe2lKodixuZu00E2uLxdjMzig53mqfVFi8IGDkekCAu4IuJEoalZw
BjHVuX89cawmwIYjBQIOFfiuMQZxElLulFy5MPh1jvV9UtcwZxemEHNxrRzF2A+V
EKmd1r2pOLwCuk2OKPOZR8/lEtzDoNzSqEpjQa8OZMJBE6LYVvG1cH60m6LqJfdc
4bF+OIhse42dWbgQNDAYjegU4NFig0OoCggvFcUYhcEfvNgAFd3EtqSnYA5jgpmO
eWkRqECjCIUjM7hviv6/WSCY1VmSXf62iURHnlhcUVPXSv2qeZVHHYOePwfO5Tod
NNiMmetMjLWZbbOPBRL2cg8uQh7vstUZc4g6UzMunIeuGffylQOaawTXpbS3zVQF
FZQCchXobUDuXjnp2uQ4lfsJTuJfmwBalpdm0+ypiGQ7/d48yS9axebom0gLEBg3
x4c1NmpQ0P1a3YoD84r17UXBz92wFYxnqhIMpzgratYGv3gy/eaLgP06Z9O3IYMh
NqdbutRcN8jHGewlu8dVUOmtRezWOoTwrd+w/Iaq6DMvKzssD6ZDq9ogeUE/BILT
KaL98TLEPfaOXkun4cUOs/QbchiCMSZVJkaSuF2Zi08R5dfHCfPaeiO33fGX/GQK
zDyM3+NtcNz0ib1sf9lRg+B17zp4WA7y0pznVCTZrdPz/emxV49LntEvf4EC78Wa
dkehKVr02VM8Smr52tCrQdUIO/5XD62+KejliLGMqn9w/yBMbtxJpVUYMJXj+F+C
jQ+gMS/oeeCGz4W1iA+iD3txs+zNyp1aIzM7eeFlVQU3WFctFciVfRUi7+hkyKZH
B4UBpDb7BwTLwHwyHKKx+FfPJ/XWhX7yQM5Zew3zSCJWJk0VFG0ukmM/dxeNUzaZ
TiqJzfeReznSMIbkxTBb7o4bjDYRbctZu9HNdM72wRMHh49s0dnbwEc1FpIFUG51
PH489f7MuDT80qqFvIwiHthtGNr7DFdaOhs2+9HxQPm+anVxsDG4MqxdKjQM4Jtb
HnpCxYNck46qKTrvFrHqmfemaoy5f+MtXVMrv6JyeOyhVnJtr1M6LBxq8kXmBKou
KVl+fVkDDpvA/jhfyVEU4OZZnKaUqmLTdSsAzgpuR53CfTYN3dqauXpcxgC1B/Iw
+qp6ifvA0/RHmSSYNvg5W8xLT3Iig6J/v7SQ0OUuJggAJv33Gtp2DRUisubfhvQY
8Hx+V3Q2TuVfwbAdNat5kaUrW/t6QWPCYp26Ao8hXvJk7X/WCB+erMZHDJGWeM+0
a+VPCJ6U5eX0Fr5Stu9A3R9rpvsJueqZ53R+yAtMvG+SD6fBz8vLqe7/cxfqlGOR
76tlXj9JX7DuAeNYTAOna2brTCpsu9Mka6o4NKGbadWOUqLDX9WCVDrYNuopjhI6
KqUG37bG3jsUACP9SFMcaXCbjdSbOWgmoX0ebjMYhgkUFFqh7xzEZWlUoSOLjfrg
RbNDtqoftXyjahcRpTbvrQFNyspsKs8ISIMfmWzivvJ9/w29mQmePnd7NRM9O2MM
X62o6y3PzvpLCRqy304AkXFUTUCfzlRAKYBafouHhZ/Ee30yk1nTxBytTtPozFmv
nHzv4kQalvLlSq7OrjChxnypSCt3QpMfHgpC4DMsNHBz4rNF2+S3KlffJi1Xqg5w
JESixmlCFdMBWiAbaGCU/9NzhGCH2LdnAsb7+Pa5vaWHCI9uTl9fHRg5/ydURAGS
+FnvvmAADwxGbxNKudMO53JG4NU4s/zGuEJyA7Ca20r3YZpCbLULXE0btfgPoTba
C1m6cFs3G0VvYqC0ReDrdB87KTXgxXfB4y3f5MWQhC7AP8bDVkRvf8BXPi7v++Qj
JWTvGT7RrOx7oSO+Hh5p4Q7hB9HriN93ZT5xcN9zxrmPEFtbRIixxMJsvWfKYr8F
VID40L62uYqcWywVM6+QjUM1DoBqIAQDXLO/rJz2ycVSTMw/UyI4rb9XNX+KWjeG
zJGhZa5ODJhARm9bgBq4+Tq6pmv1tNCLgTe/zrOgVTb/ByWB2mjCmWgVVaE18SKY
/rhD22V3u9j4LQMJb8twQ60908a6lxYaF1KLPP4t6cIE3Jp0y5hT+tveG6bKjm+q
IFI7KJEj+8kW+Ho7pfAjEXya/g6NAtE1xWzq9ap2nMLw/Yn3p6z2UEFy4RhfCzZn
Yk7520+TAs8Cl3ifwP+QG8xG1ZnB+jJ7OMFP4Qs89XCY1CA/2Ea9Fcb13RfWgI7U
OEJF7bluUTTpzFterYVgAeU1B4bWLdROm27fqN4hZYssrNh+H/8RTjmynX3IxPFk
85+3fuXumvnVs74vinbiac1q6GFqAkYoxfFgGlTkidrY8om0X4ByyLpCVq0390Dy
xwLoyi23SnoinD/7MLVzOLnAHN6Pv4wOWeXw6SoQPsXUJRxh+KOAcamAw4BH4oxr
VnpMnOQT1YPUYLM0tZcnJN0LzukMyeieMLdPbLKVXWLSKVWlA3PdnoXMd/zn7eXs
HlHc3bLHbsaH7/W0wYDB2dygxbzP6fSjEkZ3/FYOtkggAGgaEO1k65SShcdxZbQi
wWpLh6scNM4jbNJc/vOnJs3TUuNFw3q6j/ugQi8sWLGzpBWuwPhadQ6G25jet+II
hfsbrxcjGFd8F9Hp8uu9r0rzvbgxlaQULNYQv+TNr7kD5Xjr1THDi9y07jRnviYz
TDqJeMR2/y6UIWT8GSh/5KBACsF9zb7FbtCOmAjij8mqSDQZSRau94NOPcq26wlZ
S/nNR7fZs5tSAF/PPzNP9ix8LqYF73a9eg7VBGXOknGzYHvjRtYccid6WkDZSE+L
tcuxblf+/zHwm2bmy0usxDCoCtc3LC72Mda3bAik4tInHQvEszH11WkVZW6YKKhD
a3YxGeJFrEgVd9y2i4g29nI1hdhKHMwSCGsNajW6TI3/ykpA9YHccNoyPyHzft7d
yTfOHz88su1M6HSknIRszraQskafj4RORX0n3nMRLm6R/KuASXJ5bHvVSNW/ndFq
Qq3oSF1XYdbO0QscYLtww4YJdcp5IW5voLj3l49ImcIhDRutsdbZWYKjxXx9O6by
O6TfZBr3yCL4nY3CfZ8TAJhX3UZCwdDAu8uvbbE8UCj0bsYn7+3rtD9BNCPynYEq
APn5a1u10Yl8qnDeII5p8svkqTBH9C47KWM8C3o6PYvHwehwYAbyGiLc+Sa+eppW
X04mWR4lKbFp+ejzYNIPNxLGZYRgoDya51+68kOG/ThCAdaNoGiX4hLSaYkXRH7l
G9ZjYS90uXSeD0U1cJUzrVsZl3VK8znl2TYCHsXgbQOTUoRYSMoqIRETR0WxM+Zf
i1BGHrPdn/XJ0yVx5/Bf/lNLb7+lvWUVLGeh8NhgoskHjO4bO+oPpCTSoSnbzhCD
wB1vs4m6j/t5wzbGSi8qY92r2pd2XHltBZavRQjKmjd7A/hJtcfdlamalbaxhTSP
ZtP818VdK0n5HUhTsJ4L+24mydcrK9xB7u62I76EVi9Cq18WL9xD8CPca72rggqc
3x4Hr9DNvEraALi5bm211i/QHFz7crO4AVEbdvlMBKL6cnbwVenmqAp1Ok2ipX5I
WasxvHBVOPseBuQvYibRDXQ29AhYNmNggLaofK+j5m22SdSTEU94Y22Uczh35kcf
qXXBepNgpguFRA1dznp90uKgx6Cb29+PX5cimI5CyKha9V9qjdzjW+i2mJ8Yfx2T
+2q/gCQBYPAn7gOMJrJbMdEZNcfJj4rI9tHwTnNWT/zOX63WqzpRum/jYhD+une5
PvwZHssive805nevLRX9Hun2A67tlpuWniNDCEaXM4+4AP0F/xNKlfbGWO1QiBCm
1dRBhAvDeLQ7Kzfg9nZgt1KzySp7uxt1jZdveczWLxVoGeRp+M98z/M52usmelyh
OjNWD+u9z8AN/0BxWqKVLb2yhHrAfG2AzTAxOcePy6JDgCiPpnP/9VSMdL9hZhvd
9kdoTuJdMQyPd0aa38bCQh53XNOxtxvjlMRWUq1JawPwXW2EEI0WWHIn/NOTydRJ
Wt7EhECSw5uwjQYnrJ/UUumLmQB0T4iYXsJwcgkvRKMb+YcZWmgp5MMy2MmhIMpj
Trpl//jE1fgJ4966dycLPEcFpS56wAENyLYaslUO/vPwlkUwx88kVLjUkpqw9lHi
GHDbs+BLRjHZhpNncar/G5HcsgZQD66eAwxP1IW3LVr7PRtvtmBsQz8rbceEHWya
j/cz0Q48iDtvYCdhiPY9hOBE9QEc6Swb6bU77lyx11yjLm0z9cOwPoJExxZqrLii
XLGder8HIHbVVNU6Mb9dg95UD4idMaLsU0EiT1Ka8mZabHeNvrYX5NS4QQhC0nZ0
QWdKXetMdsf0RllsX5QQK9SYMrq1rD/IDdc2kAkjpXSGBmJpCklwR2D+ytauk1F7
bpeO065pz87jwixAP2NaV4LZnfiwdFt3VGj2Lb/kfHOjiJxCzZ5wIfnzvYq7Ool7
MjKyVjbNbVYugePbpJNjqmguyZw00RcFDAPxBjeOtt1QU/GG+6qh5+sGDDj9Ekg+
0+xW5mp34oYRTrfbModfjVD/+h026Ep5PCck0S5xUqZuw4xbnga5L3atykXDy4lx
Jv0hx7k0Uo+UkGhF4mkgYUJSxXqIqbZ7+9qo92gyP7Yq57ymwGp8yZ3vU2IFUrlx
sl6OU6Uz3Kl+p2lTeFaB4GROKV8a0kvTenbHG4YePNktmBf+YM14lLtKhP60O0hb
S80nOHCAYWSaSrQw5SrK8sMqjksZe2lwRifKw7JIjmoo9INNCd42vY2LfU5aSddf
od6jcI8Ie91f+x6SyQ94WC1TWt78/irU2w3Cauoem0wDPsEoCgY4ta/Bi0Xk04tP
D86MNbkXHyx0W0HRHSWCN8dfRJK70H4NQrsSG/o22bmQ6ywQoH3rCATyzzgCL9CN
T0qtfbMq07IkoiBvf20jNSD0OnFsb6pHRBfmrMVeMfvXai9rt546W474PSI0HJb/
U36Erh3zFFQwpkZXdsoFPEkKODEXGZAtxlZfjRsy1IKUEKlNIcT7nQLIQ2vKXU8V
+IdlqU4IaOdJa0m4mJpIEYb1v7jpFZyzSLyROdsovY3VWlFnAv+BL192qgYGDNp6
I4FRJIONmt4RbRjLcaxyN8qcfEeIabDIJwdZ6cs8hdXoEYb3wPTfp/TEPOadgLV1
u0C9LuWCgDnfZk32B950Il3EBx3tpVfb5Ixra49bQ4ZLEs0EIJuzeiChwLbmd/wi
Yh09hyjOrPn4b9MCrHfyFD4XMf7dEWkGcvd3Z/693TmjiwnFiNetKhaPO4ojsk1V
PVRGRmfVYdu0mQY8/hqOLfw9Jgww1ggBOfTwxM3KdxbFSQyzwqoTlISOL9vEUTmU
yEZsXTx/zIpear7QECgZzJNozrwEqLzuB2YwZdfX85ZKE6HsjVKnehomnh2btJxh
iTeZHoL5mWpwbD8S4h+vYFiC55Py0X8sqydklt04oiQrfBQI2SSSPkendqY5+8Hu
HJsCHkt4ux3MtbnUDDuFCYuvrGsDR/PWLyzyXC4SPeKG42pmUCQPxxfthARhw9GO
hFaG+Rhn82z9VI2fM/8LFRIA32ero3ltFIR5X+JhN+qYIowIy/rTUq7sNtShsEjD
bvPdDbldcafca7VbAm7w8k3Zh/SNqpxo3rG1Sb7j1/ZfPOYlGT0UnQiynxquZqOK
i3Vmrde3P+9r3ih7XYkc+bKCXh6L/2UTBa+LOKCpjXjCukQyWs0EhUVXIPR8wNUj
/H3rZ1rLUZL2MFBbOC8XrQ3pRybeDp1NwEZ4BPnN5ZBuQf9MIIknkAsg/S6piRwh
1zru21b0aTACYlKMN5dSg4PShO6IoTQpvb0C5yten2ktFs6Ck5tQtbgyTb9HWaEm
2CpAgx4H+5c7RS5NqAXJIg7eN3J+v8b3DgpBnJ/L3UQ7FpgWb/oq0wYpa4oMICFr
BzV1ThXK0YIls3yRS6hfYMHQxrhyqQzHdbLfd/QVMLFPwf1GocxRz4GYh8NBzy3D
WiXcbQ0SQb2tX/7ctddiBw6aYGpeFC6b3+eK/9K4EcM22J468x7co7KSX+ChgRwD
F7ckB3UcpsVNGtZS3x0yVogmRv5RQovinTHoO4QpuSL/CdQAh2tN9fSsWhlucISk
oZAI04Xo+S+xuAlSt9/ZzR/C1W4BnHUQSrovay9eERhsa1lLDR7uG2yCioxrnwFU
jMTMmRW6vO7Quv9RNmF8V7w6yOXArMSdumQaIimGcwVsX6NXSv5FH2X6DPEhakF3
uCSr2Rly7nbfj2PdJcqwMceEPLvWGG+UMTpg5qKw6dj4WFXXhRSQVoVBN5OtoAMq
5yjeWem+ADaO1R0INdtFHcIHzg37fy++s7VTPDrIBc+wZjDT+I/bFgXWcVtPTgh4
bxUU7kgpRXLrYOVPTa7XYPsSTugStbWn7Uos8ntGuX9joA/7I9ITP8f2zQMFxYCV
sU+sbFBa11zTPCIUv1m64wdF3bkXiE++eRUkq2ld3e77eU/LG+ULppZvBVdK7ot+
ula32MnziIz6QK4hlE0Lyxch4rmP8sRDMErErD3xGCfaCef3QxDgEx1XkdE7Vkss
LJt9+A/l3llXQdROXvc6FiEVHCMmXk2k0KynQ9MttIvL9DeGiAO+51pWSJmAPL/7
wm3yR/1jCV8iFgTWihdWDiTwEi2C8c3SYSbWamyx/CB/LYmK2L9zT3z6YlD9OO9O
p84JaChEUgdeTg9PUIe6GoBx0Gy3LqtncNY/FglM9WHVuheEyAJgNddhz/Qzq8zh
XPqP9YASr9zBHP8dqp9yOCwjo83PUBQ9QUPWWTmhvhbdWUbq/je18dzQ40FOxo2m
Rg89D6f0MvqdvvRme3/2imlmQO7UKuQEdTuCAH3QhilIJPyl90NyyG5Q5kAfrc4P
VjYp0KdhBWJnmh/ZTt/911rN8TwNXRIc7bEp4Agyzhzg0bR1nDzapNKXj9npXZCP
JneuKrf5n7ZlRKyM4SZw7k2mt9sEbWvcFEZMDxBg/O2GZBt0I6wzEeo4+wBbagFc
sWV+8UpGMsjmcZCR+gR1dlbOKQuas0ENHPnwT1IgrA//AlYnkDZkZ6qGWuBoVDEL
fOb772S7Ve5R7a7BVGuHThhEfed5QFx3HOsfkv5SXoszADp9HcngL9Xx8ZPxH9az
gBu4rd7XTKhqkfpgvcHgkpWxmTSz6iBaNwaLvqQWq2wUBcBnuUZyMG1dMYZ9+YIX
dfk+moJbOiyFdOlSabmldshupwfd7nKuDZX2cv/Ng98uyukXVpPr3ISKIiMTruJ9
yps471Ba1AGc7u0Z2qBgXS49PmAkyhkkLCoYwlhSZ5vqV3fsF4eFbLJ0AEWaNNtj
LqaTsDYp8VnUm2M0U+kVDmyPMYKJJKehm9qWb5DOjQeP28BE7dlL2LSTImeLiYhM
Fw4frRdi898uoZQXhUqQ/tkMFpl32lpaPpbRx1y3wa30B/3j1MFam1aIu6vUKyiE
3BCXFMfKPDzuBJpX68cUnv5V6UUTBcxhZFbmO4lKgYdbZrNUQMs5PlMOIH0J+iOB
ZblOahLwx/GxyD7k6ygCrKg7TsJjYU0IFojSPrD1TbUG8wq5zRWxalPodJ6b75aH
cJ2+dTIEENoJsP2Qykk6KjJ4H3UlkbMl+d5djRWWt6IEQTwnW/R5AOs+GFdpZbp4
qSynRJBSQnqb0nM/itjBVxUvCYwsfmGK3myHK0cxWvWZr9v60J+KrOPiGuY8aTB3
kKH7pK0SPTk6cw8vYVs3p4FLCbQwygGNJCLpiG7rCRkjtWtYQuC9oQ0vranFBh3G
y1HR1N+GMVWDeswstl2wUeqFRDdB5gigZvyN+dPOy7al6yYRtxgrWlxbASbu32vZ
iJAy7OkpHi7vCsTOVMULlqFuyPbYCfD9ODXXh299Gr3PxYA5MVDE9jl6BIy+vG0g
BPQYEVghKoPmB2mjNTaS3k/teDZhTVgXZbjNZKUjVWgaeDHiE8CdUDMxD58UPj42
T6Qj3jQrPNpP1ggIvVYWow6gd0RvRHf0lsqheVVO42xI+4ko4FmecZuOX2Od7k5d
6g2aajjl0WFOKkVlHUsdblBqyOvQFfkzsadVJN3hsRj7vXFKmWTe+dcUaXO9sOGu
Asy3Wxl8IGX5F7763ODNUQoYItNM5aHgRC8Llrs/XJN8sy4Wost1JrL85hIIUzKW
E0bZp/1sFjBCbTZHejUrvcf8vsvmgX/DoDnCCARJ0Fss6zvmR7dSC1l7u1Qd+WEm
zur5jRrNNoeRelU/SnN3Zs49mDL0zS9m4qhP3B/zaYaS5GGwdBGyGvyWkIbAOHCV
tC1PwmTy6X+UkYkZ5AqIyLzeyTZhwYkLgRZX/EEn68D5hJO6D3TbGTrkS2Nw0gGr
PE++X6re5KhQWgcgYm4rt99+7cql7jzENz1M5Ycce6P+Ee0QqpBT+huzw493fjw+
XH6lDgpKe8rktdvby5rg0mj18vCSCgw8422wuSHivoLwTCSZcegmqqREHeanVcYd
iYdyTcOjLYB/eqoGKLQhp9odafk+i6sTi5b7aYxGmlTVusjeDHyzw7G8q5+SNOSS
xlPu/vGW6fIsLnMGjtiz3fzgn/lhAcnmdUgyjesptpz/JKfc9smhKF1WLsmQAAjl
jwF78Wj+0a7hI3ElTvNCzjmoyzS2pYbJxpnbmfzpihUcdq4QpLJsVGHMRLtPQPcp
dGtj3b2VBQiqXnhPyiEXfKpZQW2YGM18zEPBO2iLbWUwyySGbiaYaqt1a687yQb5
7wr5fVzm8Aawf0l0Drkmld2nkBfpMBWj5uXfI8TEdldUVQf69GP2UFbbnyTj9eBN
el0rRhqp+ftIdtSf1HdnI7CTO9Wv9zeeQbsIEnCly50zVwIfGz2hGT6Zkgv4w3nw
gaskMoCcdsXp+6U4aK52v5KThr0MMVjelGerO3mDKH+SFccus0uT/LtCwrmIOG4z
iDsSFUyHt0vMHsqTYuBOPTuByVHRLkAYQUmdENqIiO+il0d/BDWPqCaigY5g5iX2
J/huvEyW/jFIKg8ZHUvDjfOBNYjvw6K/uesVHIx8UsAx74BzKNagE26+FH6XhB4o
d/fwR5dQXjSxjoOlYvMeAwFHV0K3bk5BCn74zwU0KiVpm7YXSorC33ix0RLSk1Zb
UxIOGQhuE7QIgHJwE8tn9lqz2bTDmEXeM+X6Amndz5MOluybHPfHGXGCVvHyHBak
3eEWNBkWVC3Irx897Pb+DQOp9DVALS+8NidsILuZN57X+MOkqh1Gmc1h96ilnJkr
BeLaCHRB4aT+iiFQsbIJB3dK8kA0srFhVRMboVetyfCWTzVG9hbCr2b1r5sWq75h
cdoLx46zb921Hi5jd31TbobnwWdvqZIh/kB5d0LH1tt15PTdBZcyYcCUUU6LP5xJ
0aA6xx/c2fvJKKSdtJYzy2wcsZ8+vje07v5f4xC+MIaouk9em0Lwo5LgcCV07cyc
e6rvzCi78I/MysDM50UivG1YRgsv1FBAhpMT8DCVRoJq+otLRtDANcMj4ikRNNbg
JucRGj9klZWQbWpbWTmX1wgkE+R6FSfSvq71KeR6sHevzygfDemQR3KzCUr2w+7z
8E1m1oThcEcYYI18E1gDoa/t9Ytpzo0PT/7sRVmZfskO7XrOzBWHiTAs+Is4UXFi
cLIl2wMbZRasOpxX5HNrDdCCrjHIbxoC5qyRJkDkxK/okRdNHX8L1DfgFApPhO0y
F/QlQ7Wz+QQVfRI8vDPX+6UD/JVqxQ1dRqW9WOhptiB3k1Pe41Iewpm2gOnR7Zw0
x1yU/GKmjgPeftDfy4bB9NPRj1oUVvffJ0LdtBu23I9LYpkvst4EDuK7icdD+iD+
owA/cID2+xOoB5WntuePPD2Br6zJ2S3GK9O5xFk8F1cpPRp2GY1PoaPtbMf0wCR1
yMOKznYrJm8H094mq14edh6DiL02r5VsAojFn168GuUuQEeExFapc0edonchzVPH
TMSwKA0ZZcf3Jl8Cm1LK987Ve+rIZbeFG6fS3mSfP53RBCVfYSjl/9B8vuVwoi9T
pa4PMcNadIa+2pOvoAVNUXC/+4PPSPCVb0Gkv9/F8uOjAd9CMx2PLN+eyhwiESSN
6UIOXfgr9goHXJeWjrRZTf7Vn1/FXB/F9LosjQm8e59ee4+cVASHZOe3ba6epYaf
mHe7IJSHaNJUuD0iRPrFVucKvsvUSZDlIS/QXrXWEQvyZmK2iVa9krMNce6kT/KC
iuxQqQdhk9Qr0Yljo6tguO0lcfEfNbXe3jw6lIUUH13CQpWimOvwmXlscQC2WDfc
Se/0BTd/dnMbLRIOwhntwTZXSo6NgSC3gAcvBrdLXhJwG5tGq0Et46AJAuJQ8EYb
HZx3lPLU243iWuHNHxQAjQjqXKmKD7daNyMHn2/lw0mK9+/C7CAyI+FXEcvk7wiM
3kYXh+blRDPZPcTHpgc/GPkV6dYoJvwdJWZJavrvK472ERVUmRKXBY7g1/cY9I0U
ujYhLSZWCe0aAF/kZNfPZ+efvf8x+NhfojsXoOG7HFjMA44bkfbAIVvv4Jht1a8v
pZBxgSBImqnOsbxIjgtlx8dpNbcv0Gz1oe4FjQDrPKOILbsDoogE7hLAWjySnOW7
k07HRjXFIj7xNZ5V4cwrmXTDLR96OGUKUdzmwaxgJs+EimbOhMN6uO6AHPpRYTHw
k+lWZwLBOF8D3IzGHUARqiL6CvPNPRNj+2t8HSyMM0w+/HhDyxFrBmmCx+xn8Uez
AY7oO4saPuLG1iiO8MvzzSVpJmtoNL/dbzWcx/OTE/61HKFvF4P46QbEvZgLhVFq
ld3s8z5UVZm0qoab5yABsXRagiybqS+tIrhTWzcs29L4n8z/QB2aPW8GBQ94hrUz
MG7ELNIx5VILL1a3OLHVudi9t3C/n81J+9uXB4YD2jvk2eM8SAAGxJnpJ+QFIQW/
Bq3LQlwC6ArQjq72SbD4FoSv2vytBbjr54OxuuTKzMTCN8urWSxko0yoi23Kf4p1
MJNyYj/bnUWXUebgScIfZ4AOEZKpEwwOt4FKT1RIBBObZoZLbswbOBqJUlja1r8q
LG29I7Uxl7CRgJr0Be1txPVs8xkXY1TY5t5Psc7tb42h9Qj4QaCRPNLwCI5M+FRv
+K8f3a3YUh1HnYu4QVibU0K2YPePngCBd1rr7NNeHepLt/2QSKHu9l549/r76lbY
7mX822xIgfDM++Nd+0KR1VRk2pYIlGR95emXtMunOPT/dEmIo59wZP0kXHRhhO1k
ipjDL/D0uISDOvkqjLqiFTN6e2XT1vcCsT92Tv9xg0R8QPuPg6MlQpq3SBrfMy9r
3ew5lws3AFVvgQguAC8ozDbSfAKy4nu2FEs8FPi4LixnTc39Y/Zhlz5oz9pFsp/8
uVq1x6kmHqzgadjigv9WjgOksOGiXvXRu3Zr6/wZq1K/pL8hO8RlsMaG1KfcIJ+q
wb1f/NofAtvAvLk5Pl76bZ/02K11hYbO12U3NnX69R+Bnz/ACC/08Mo+QldLiFfa
CGhVxxyrnzW5yYvfTjveOwIBxUo/UYZHjCQ0VYnL+FrC4UtIIQizdxnBILyaOWa8
vMr345Nq9r/trKF4S5K1z7AEU6GGIvQy5tFjwtcV/TXQG30tjH1d1RyjfmorQrZL
swnCWnjZurioLClJOwG+w0+GvtvBguZ8OKOs99FTlyNnBtLXho+ubBNX/KmDpTS8
2CQmpf4Z+jkZO/6vFOhGHTiiGCArWnLPLKcXFLXiComQmPp1/q91Ot8YzyMeKbg9
hBM4jF6bM6TefO5p1RgrkahlUWpw9d9BvV7g5RCFlJMC4HHn6CDCTpCWePTm1E3p
9/jWeSrQOb9K39a6ly/D77tsO5jLpj/rq0QLKIgvWzKuUZehf44leBTKw/U/YN23
FvWFrRQyPaxx243PyjFTC95uUaFJ6OV450/4s5lCPRWOOk9ie2P9hGRcl7Itprqc
L++WGLm0Uxgd1YA5wwuuPV4N9ymyCyQRwgJzkqDZ/ElehMziCFid0yY2h4Vwhuoz
7+SP9TlyeCpGUXrgu6imWzNoo1CUOm56jJmZ4wWUTULZJcj8dU3fV60BIICApWX7
wtIWxDC+nGL/1pyq08KX4CX7zGZ3l+yubdX4s8c7zjbonKxWyzwq7yot5qTxwnpX
Njz6h12Ft7ODd16bHhDBgXBfSJsbToKHH35wlGwZYIaQr0ICo0yZ0eyBeKTfpGNJ
vleFR28GWcx1xHDqzNGnlzEW0uot4jQU913vyFy/K6ggQ2ZAlXBKcLMhZAF3TNfT
6juwidjwhObJnjW+To6gmZ7m/glUtfSjsWiZCeKSA6a5mBaYKnOPk+Dsb4WGlPoi
H/HYkGB5nSMS5hbXeVPfSJU27PRAn/e0OgJDopeKHkqMp3u6QrX5vib47cth8dvH
1xYAfRpiiuMrWvknBeRj3aFj2RLmm6Dx/KVt4Qx2KoYotCBRNLqhQZYFE4uA1Sep
GDABGqUx5fZi6qJT0H8cyy3xKTAUBonKGvPVqRGCDAg/m8auvzZJA79d+fEk8jE3
dJOry+3uPCuuuT9gUx7v0rx3oGS2RGOBAlrY/zUz+fuwzBctN7wTtvxOet0ksfbs
8BRn1NpIVcQ3eEMbY1tF7MzcMXhlGL6dvDJC6LpRo7EG/FJhFcZxvmLFT9tk/R7c
S+Km+c7HZcfCNsFpYlaAY04zu8n7jHI6q7GrtyeeJUjEnID1V+yDwA+voGu9FevS
66HG1RRM8W1eoLiHuVdu00PDK9T2XTQofdLBfVwwxwwcsTkmAxXPPQfZ41q+UwXY
8LH5hyIW/lgd4OuUSxrZ29w8dKuIqabZYmH+1bTCxNZQCGXDU/dD0HQvz1YkM28j
EG+VLJIFpz0QVWPdlx9Uglum3CDzERfQxTpquRPls2xwqYvG57tg7Cvs5eh9Dr9b
nYZdqihb0aLoRwHiLqNoisZ27ZEU+zTiJPDaK98Z9Q3ZWqDYutZlNquET2jx/05+
Pu87RySkST3rt6GdlUMEYTaGq8M6t41wNllamekRMA0U6cblWTNRam5ePFPaZiTh
woe4HSDAImij615rTVA4hcqxX9yzFY5dabdnq89lvGioP+UjTPsO9OoKzqq82DeW
kpxZ2c0GS+/SHCOJ2wKyhTsvKz9ddEKRNIsNfQ6XPVeN+H2IMUi+WNfnjecwlgeI
ZTkf7IEaHVD+wVQY3k70tNGDDtR35kVas0YeWlHhInixFNiT0CGtsoFrA05C+YW0
VuhIlQKVPKRHD4v86EsN49J7zTqFE2mIGHJ2DoISwC9ixh/vdZDru5uv6SORVBD1
hxzFBwyVbAMTGSTQ0CaNNGTBQ1YtzAKq3iJTMZuNlD7oHwjTkQFVpBU9x0m3M6bh
c0Szy27itl2//6kH5h3KohmRcLnn8RFwSesfjyLuq42GCCQ97BKKTDwwY9vAp4pM
Pg5p9xUS3adBlHeoKISdKDrQ44WnOmAKgeWcg+Uz2tUyEResV+vr5YXAuSdoqjSy
jY6uFTmOUs+Gl3Qk6nn6lZcM33fKQz0AAjwLKMySsybWbKYC9qmw52TDmwTt1Jz0
fQUO5P/cwuGVcYuvbTKpXUUP3bYSGCZrDiwEoSqlB0ESacXNpTxfakrz2MECweu6
Qd7BDjBSLqhpqJCkGTqHFkfCwvo2T1UPA6TCj8aGe8l74lXSrCaCiTNmZQf7JvSq
NQX205l4bnpeU0cfVqoIkakdM4TqXMjySUUv37egQ/mJDN7V90WYrOzu5X7G03aQ
AHgSEg+XFVt09pe5V4MrWit4h4fmMYLQob52TmVTZkYcrX9uIh8LZOdtB6Ev8IdU
TMmAiLSNCWGQR8hXCHwGfmR+LNFyc+LkyassJmc0uf5vECeGW4rlDwKae9f67qnU
1FJod0agcCJImSFn3yJOAW6J6rk5f4afkwgvHBU15JcrwvmQR6f5RGzehzM0++8J
JRShYx4KCLeimTsUyH9R3Oth3N+0GXCWbx32Ejitj3eI+3IUn5d+8Rqz6aKJ76us
ZCseXwucbHXue9dYund9Iot5eZaN+wiRxrzJYrBLzpF46zDVMMlNUDnb4ia4/TKq
hzAp+KooisrROjRJY9Vq1xLSvYMDz4GpzpXpieu8Jq6oLtxIcmHa0FhAPLD+8yty
+VygyuzpxFLXngBcBwQ05PLMuBVVjvFUrQM5/L+x4ygszb3PFv4fJp+YuhMCR9YB
tQ/x3TsZPzJwzpm6zuJN34bws9HhGbnq01v1eqTzbc6DcRWvYFs8FkrHYg5aND6z
YGvyjXwGH+hctUmIVtGmqKNPuxNi2NF6XdnhMzBcyPtQJBhPuPqjltWFI0YUeIeA
PUQx4CzwL2480M0ua075OJzHj4LUBS7MyZOkCBDFBfkCmyp3JDLLmOyZ1dNjvLC8
i/cn6ZrOgP9ZaCcV1rGplFNsf8bry+za8tZpjSmtKetNjLhlhCmdxQJj9nLSm1sJ
sI5fRvno5CKMoIItrvDH9btsct3wQNIkldVYCT8pcuCe/58NSrrwR6pYJbh2IWbF
6ZmfwK3DdSk43XqaXBw8TVsju1NKO/N2CRLZN/TW/2KVqh3MufNhg6GtOiBkdPC9
D32WJjAtlhLGcWsTK6qMND5EKlTn4mURvVbxcZo1QgifCnyzZPCxK7awQs2qap1r
TGDSKZiGadMUhm2EPHSPqjjKP1munyJ7LUZ8D9nfTrqAs3sdl2zLcldm+JWLvD8R
SVl6swC96kfE4ah1AvAef75ZTZBkzEhynTFLur55K8fDhPq5bcW9TgGE+HrkXMse
FJdxzmyUiiOrNAe3Uh1fusJfArE6wKTRwHsYPDo1LHXkBJY2KyrSH0h5YxakNFhF
y2IQghSj+m8NLtzArjOmzbLhUBV+hxhopXZKYAZXEORM2ci5Z0PuEW/K/FmGLUkf
uJOwE0LzK/axlNpYS3SoHxjkAmWEa8qfbit/ooB/HkNo47EmROpYrk+PQ4DQ7i4+
kPOAD/l5Gqgftwg2x0Nm6J+9gLtQnyEMz5Rtz3R2Bn/I659oPM0efjkZEuUEYwS5
I030XNdDlIXI3I9eIZ+sNq6r6R952lAa+soqqvHS/tDeUiEcRK24gT9HxWcc3l45
nKXj3mZf09lQzCiUcnXec8hgZ0ubw2mycqJ9V5IbkybaqRHOKexrVB7UYIW1osRv
EvFVGqEqI4mNVSCx8jSGcf0rphKj7fiaZqCewHmbBVnT9FTDnBnNc5CdBYp6qJeE
/xkmExxSyp4+IcM+9MPYPU0xek3Hg03tm0Ky3K6JScDG67g++geB5kL1gwagrfGt
qu4KvBHXJ0Dj8+Xgagm/kOo5HnaEIu+aNuDF1x1uJk8xRcnVjGepQdXWDv7GWhU8
FWy9BJWAFOg2+plL1gWhOtG9IdvANdLzflYDcoBTqCg+qi6DCfGwcV09NN+quotj
hvp4vVLobaVwXnxWYJmPwgAcpqdCYzwAY+VM4UwGY6Ty3vdYmLMJwRQN10+cqi10
6uHeeE1PqNRoxh4d6wsxmvcoD3QiIGl4arlQPR/J+5yt2AJEZKg7H2rq6+uBB3K5
fiXKLjtpmaEUx/N05wXZe4w1gByL7MdyXrJ9sWEwN3tvdblDp7Vmb4RRGu30gT+M
RggOfb3f7HqfrZfzSp2b5l2PFAs4WCs9ss5q2wnAXopYjIYdYrtuvG9II5XrWCtd
aALY3v8ZolCgOta7UqTiVL+QqFmEp9/F3PZzpx7qSXnjvxHpcfikSaEn6FMqDXOH
kAshvkpNO4B7KItGvn3aVF9ylQQuWDQ7nR5WpWz+FIMHy94LYf0GwQtktmeLapmm
FqfUIVGIsaLtpXXgODzKfnK+/3A58/ITojIKYj36CRQFgUTuTLHze9M3ZstdjtbY
odROXbdvSnScVnySvqLrN2VPXEVda6FraiYihvuhCUK0ltQHjtxJObhZA+RXh1Qj
JIOR702NvuufECXwZI9Vb4b5Dfk364a3XbjGL2m86egS88CVQQW3mm9T76ErYcCG
uEojYzA7uVYKFMDs53YS67+8x3Q+63bL9Ig+T0POMP3eo/KUn1EDXAX2i9zJxyV3
kJu5sKsJZ6WxX5yu9SjliTijv051B9WBwy5JJDCi5XUp3DA7VPgg/KKTfJKYsK2n
nH/gx/Cmngmh8WXULF2UsdGu6p34VzMLpeovciObHW16f2Z8nMMqpDhSuEOezNft
kpYktuwNoZuPB49KYsJw34X4qe7d3xhiZEJRhEBF9M+ClHxq1IoErUYK0prT4D3Q
Os2pDcIyWbVG72gLqT1T48LuTcPwwoVEOYSxX63rcG6/0ukifT2eKycfOKi4sBpK
T/iVy2QKiDlMm97yq5nZPWmXzDC0ZmBhtPFvKfKVzQFETMSEXU9+0fDUYidB0C7s
3+gQOU0OMpfpOeZ8t8jk4JRlHOJ+G3WGgbnMbUz8XIiDoa1t3u0lXD+/pXoe2JVW
gORPGjcB1nmfmj6ukXQUTBjd4GZ53nz8KDVRWZihT1KWKxBq1U8YIc0d50kJ1olr
DPiCxN1cImtIqD5SKPicmCfy5n582/4/RUiaFKs43Gqh5KdRf8D80B4BjS/97hrX
M0EWEZJgG+jzPq3Y5dcQR/nu7OFh98yJDhC+dVM239KpfVjojTryjYlefqxEBKmr
TJn7QxyTddx8iZvFIvHpzHw2csOj3e0fdtl8AtNdBzq5NTt6Z0OCb9Q1zujdZleA
nJWHpzuzslwOl7f+a9i/nivDBu9qZx8c+Yt121Fw9rSDGhfD8CJZlpKgbJKL6Wkh
jcirjxx0M71m0As7/OI0BMc5Oe0995jI4YOCAfqmUnyxNg312NR69rxJuJDKS/qE
3Gowq4Q4zMXRZg9Nw34TVpQEl/zHOgkSJNkRtFBR+2JsLGqg09JrFdjSSiwQICUo
O+da1ei+5Tx7U4IsroOJpNrBgho60ot0XhfmNiB73A/37vnk4EVCqEkiN+gjogJj
eFQvps8YMv8EN8SnVJrJ/4rCfXMytQD4uWsY8ZQ3wRZxVxR3ozIm94bmFtIFSsSA
LJEGfIBn3pgc2wnTf+c8akSiUTckdbAbCTx5wBC/ysHzmSSz1IDaf3KsrZ2H1Llx
fbZohImA1swJiCbfjr1wDr3NZVDd2zkL0KqSvFVyTpT4RBkVD2uyjXKTDT3Sm1w5
N+vazkHzEpLCyDpfp6kjA0GuwqvNLVTcpoJ0B1uVnCIfp/ZA3wz32BOfde5cljI6
gNDew15qCGOKfAK9o73mA6OipY2afx2EAPGGD8TdazVBjRGY4q0jzaKXwwy0Lf9W
tjnli+CGF4A4kWzqzNZ6PHjxfx5frGC2nfnUEIHHzUuJGUE4WGFNtCvD42QB1s2E
yv9n+BUUcLCN3DA+V53bCJDor+Qcfr87dj/6JrAOmKvPotuI2+rOcG/Ju5zAPNYc
KHJN8EYr9TORdKCYaph7S7T7R3PJviXYWjxvasl/fN4M1BmGZxk7nAaEctt2JMNX
D1mFBpvS3vyIGhlC6zW330DAJmVUo7K5JBalHg4NH4WMO72cLRbacIcS4KbOWEPL
kV8ZCuEp8j+X6Lei3R8RsxiDWNX17hG8HtG3OAPCUw0TCuhvlnlupnZ1kDrLsG1T
rdUB1bh0K30Z+rr6x0/YH0ctrEHQsodJtncgK9HhR1FaVbNKglFTp+HiupQ69qWe
M8OSxawFdDQzDHNekCOvi54Maj9VElpvad4HwpKkQiHFnf3RHXUZLnRiX5XpHwkL
NtzOgqX2XtWTNYK9niNFPdIUkKvS5oUqA9hdtKdBt8TiqOBJk6EXapiTmzC9SbxV
lbCP9A1sBWbmuEqEaOWP7RsB9rVYR/5ZmCQq6+nHUBHXemWZpTEtVhRSeTTOfz4+
F6NWj/DzWSw0tJPl9JIGsHWfrmTMFucc49JfW6j0HRIcgxgSEy8bitYAt/gXDwOE
Jm932KD9U8XLUyLwna6ogrY+WgfNAUXh1CpSE0i80HezkE5zt1BF3utLOUNxL0F1
WDOjMAoNdnajGjG5NP1oFPFPV76nvAnH5zIyLMS/NKOlsxk9hko2+lk6jRMvtg4Y
iRXB2o3ooNpPXni5aKkrbMwSqW8NAt2ybVkP+f4ujr+pMbwn1QqTymkjQ/nhaYZR
j1ZJe5VcF76u7JBatQTp2pmxhuVsqtpyZMSRO4iqx4haAzM7tmCyZrc0EDL/9Nuf
yL7QAdV3e2VFR0TQPrgl38MXqAZ72Ed4/p7U6xZTSHthmKj9/fcY0sRVYcEUY0E+
ZISYM+l4wvzpFa6ZeT1snzNFAlOFLZF3WcShffqhLWO1/9cpcz9S9hEe8olZFtk0
lJZ4zAYBwpHYpCwky1TeZYuTLNErbngUh8hLuo1mM01yrN3cB62OPcQKtHGvoR21
e+tjsob4dhpdY7nx3m1eZ1nYmsagyee4xZRNWPP8e4rMBsblwWz5DLo/ulT2obo4
2oMbai08+7gqZvJEYW54s6za9md9vBzm7qC+dmFwYnR8/2vCkdosQFg5C/Matka7
u0o7akJhdzBnzmtChfmQmfKr8udARkN8vMzWwm+X1l0+EJIU4zMFXLQ5947tO8Ik
XkWsLJfwFptb5Gm4HHlD3In6a2XvVMBnnouEdE3jSH9hecIetHzPIrdYBtnuC4VX
pA26Q/aDuyzIOflXue3Gg35XWFgeW0H2EJe6ra8rChKwQl+FrB2tHNsRQLOjrTRl
o39SH8A9C6UIoWLdehXIBYZu9UKUdRw02TJEFKQ/ROGhOB1tSLxblLSYa0/a2zz1
Jg5/j7ibaqQKY4A2JQ8HLapwvgmbbYKh+1NF/Txhb49sTQsLvzUAfgq4/ldy+UJL
ifVpn5AVtq06eALyk6NP3JRmTVEzGxko9iO2jy5HDQIyRRwrvk7b3aGryQxzn2mi
6iV9044pJj4v/s8mQHMchKNO7c//5fr4/SjBiG66blphMhg+p+JF6ChiZ+hnNNDm
RfhnnXpaihXuCG1sYrDBaWcPBgBWGFcXPWwEHz5NbiBdLoI92rcx/znXt/3PUCfb
C+AzkS5RC8u03bsmarHCXtgRej/uPTgJtD9hZn/bt87g/MLDqAnxlGTZ8Dvz/my6
bsSiipMAQgakohpW0Ws5NRX1g48CDzIYRM/BXidTgM81i/WR3Z7HfE1v95hxM6D1
TMt7lmNr1FW0ro954uZpnn/1MHgftUTDS06s2goL6tKH65zs1JrP/mQaKbMd8Jt9
T1VLurxD4P/9SuyQfW+Jw4TnBvKHT1eXo3S3GB+pe3LgDxLDDAx4bv84pow54bK9
fDz0faHTzN8mOHSU7Xx94Wn4gbcb0pN/uy+Nr4COECDif/7WYBLmWKdFfMHAm72K
E4rvaYAPk4GexBIzpwVA6YF9zrWJNNl0HHv8ehMC9IHqpVJMiUcGR5CLSuT+IpaR
BNZDUfwQ2Zt9ZHDAhAaJvBrryz0GVvc3FrQHtiHJFtjIHScWGwDmUGZ5t3aFBpC9
E4c/L9Wt5Dq+rf9aojXHuZ4a/sViHukRVOvLXDyivXinEqpFTCAyqctvwChgxyif
/9TfqdeFIu2rw9ZWLmsxdvrAHBH6H//d2FQsDe76dUvuf6yuy/eseDHeSuwp7r4B
5Gc3fQ5c1S/OUOpOQF/vLR35S8B7Em2B9pNiw3Q+ho2TqzjXGOXGn+h+GIJ8v3pO
otC48W81CFiYV7PU3TN0O31loFQp65SsQ8eI5DXg5o0JJ0EgIe/xqYlrAPAr/Lgo
vE7f/l8pKx85S6bUhsXordik1A9OurvCabl5TUoMoXEiYV8QaJ/eQpxjm8Tlc5nL
b1VH6rDxQ93nnPZlvBR16GhlW0XsD1Z3NIVi+qjj5cUIOoVPGuJCITI1a4AKgVy7
LstUinRg6aDtPf40oJRmcnr1hpCZfZhTRvyWzZs7yiAwz2509ho1YITOQI0NZ0G9
gCtQXBB5s9ZBNw6BNswNXvwh7cO73m7gTuKYgsNTLMLOebxQ9eDIY3YmZRYGvp3z
4n4oAD/s/gxAeI6BpR2KPk8L+T/PVRDVH+6USP8tRSNuAMQqlNMBfuOLTGNyNwcO
I4/MJ/8MjrUIwcqBE0E1RKKrTsF5DFbP/va0e39H/c5hmPddFski6OeVGa30oAGA
bF2TLMRNj3f8fRVaQ0phcn04sl4Fdl0iopULRQxTdd0BDfPctf4CRjTGof3isAMA
V7WStVo14bqALW269hRwnBkyJCe23x1EX3MjqTwvYlbesK/YdEHuKBBOsWtN8B4g
aM9Sh6vmckVoWQQvCW1Q7l0vqFzkGHQG9PSp3u7gWY9/XXIEDhHsbOv6EzjKjTJu
pCJVizSISQr5+KFX6lgP5CB5IPoKGySqw4vgtKacPtf4DfDi92ag6y+2e7DlLATs
/CUc6s3Pkn3V75mMNK5Bea3jtPfwi6YxIznLoC7PPZrhM+WLLl5mxUbyEGfOOQFY
KINHo3zHeADj1+Wtm6WhJaPCEMohtT160ryOBLKIlaImLvgbW8tgkOHPYUU2kv/i
mYGVLiMcWr6WzETcWzp+KzgHyf1/iIZs/Ox7SVQ6VymKI7mDosFjZw6NleEwB2dG
5tJ6yj63SsIFMLGjy4tM/LmRAPOxAY6Xa5INREMFbC5MUhn6x0qvhbLPjtSDkdcj
3UviNSPoOFVHn617GUdhvmQGY93J82Y+mrKQGLobPIjm/1MizZmO5oG0Nq2dS5s2
IDVhmJHzm4ykQaT7s5xqD9nPzBL8ekqKmSX/S73n+m83oZxCrSHwi2a3vsJxlbKc
omSxgUOX+mHBnbPVRBEdxuzF0huBn0+GPuFC6o90xjSAAuCCMtKYa45FWgSHovQw
1H58/rabKcYp8SQEAavSZTxP6Hv/VzPOWKuG+g455AR79mpWSbyrI8Ox1okFXhmk
a6aO96uPU1Nc+/HJfOW3xG6I5FzwYu3oFybCdde+2Y7AbWZTVaAKsJO3xGQ9lUcx
f2Eu7yIaI/hlUc8FoX+oGWhEQ6y0EHSrELuLdCwH+2pw1kaf/sRnocNV/mPAA85X
i1joFK3+/pxEt1KSmmY+fYH1T2d7Zg9tULHGMIkVFgnkNl5g/Y6RtCFD30d5A19o
U7IIvDfrAwoB4kdZ1KCD0OqZYqNV5JOmlL5s/4hw6Xe/DLwRRHNlROSmx8eUCf7x
ChajMFMkQhBgz8/wwrpM1Y9wwUVZ4ZwQyoWS2sgHQB2+dcazrfEYtDc09JB4svJF
QW7gWSHWMjSD9OiAV5VQXmYWvy8eL5ZR4FK6mod/o3oAhmkcY4GVXdgGQXU7JhP4
MQRZzOG/81IshkRphDnwm+K/3LUrYgscLkUEa2qLmYra8UcT0JSOIjrgMPz0fFkY
8u3bUIqWv9vqHbAAVhZgqnhl5PjJMjzg9bJf7TMZO+gJsp+oZ8TawqvydarbOmPn
PEnfa0yIeLIXjHvUCU1QZSUUS3SzM3de3nguqGqvwOMEA2+RXNiT5OwT2jcp0eHg
HpSe4vjQ8/3aw7kgYGlC9Giph5v5p+5t7XLaHBVl7rqrNcdEJli1RI1RRtSFVTS4
BFfhOlRIxe0DcDo+GxKKNb28Cr5Oh43c0U6bvqXEOymtjhiAslVJd6qiH9vaTGdj
cZzWuJpEfPJ2pFENrNA+fX9pAHjysM+h8y+1cXiKiyVeseZ6X/wpIHYx7sAXqUGB
767d9xSFTsCKDC1D5kbSi4IcGVZYXRUKhAcytw/m7GjSdEezz4iV+RSFXAPxWGvR
apcuGF9iVK6mxSWCE2N1p/sPdHCl3lC4T44p9RjOmdu3rd93VFBiE/fWXOZvPXFe
aaMjtwCBgV4CjIq9ELG+iQRTw8M1c8edJfujbIdt+BQgJkljWJEBKA0i9zYMb3vI
DhEtf625Zqkxc/rLcQ+ZU1xYqn7xuHAdiZ3z1DcNL4vx1a3tl+6yCgbbgTP+MCeK
vwlV6ocv327T7NdTe79KUTXdcESmdT0FBxmTQueYds2NspArbSvAb67AY9Q49+Pa
9is0T/62f1OPnRALvEMtkKQX8vJUEqC1FWDbgjJQEzPKBybA7tmwUKiFlQhnCewf
jxOiL3Fr3Ik6htfwSTnFzTbl1uMkLM4uE1ibKEN0zONTiLvVoVO2JlzdEhxDyEsH
jTitboCZTVsV1Bw04zcMqvMQtXeUr+C+UypOaA0Mjvxl6AF3wmni346bks0obwO5
ScdqnGf0nuYmbqCxDPXkOi7cCcs8EFixD/bNhX2Niy7yAUqdQNmvmbRZV31DP7lO
HFbmFYW2Ii18qQO22Lr5Ov2/sIixbm3gEUchKKfVuNEHg095ooghZhcX8O/JO1Os
cxt8C5Bs/cDNiHFW/+3mm1m7SDO0AQtoeY6mDh15r6mJ3gptjecMc88VUKzQ/zvy
K+6tj8NKmumihFEmaqvpaJgeTeaEyp01VCGhJ21upLxDR6uj3WcBSRc/m/g6XxJ+
TwXJP88LJ2rmQlxeKXVcDaP0lg65rP+DuHA/tKJB8DxWo78d0Rez9d5Pa+UpVRGO
I3Uktbx5nYlwwaCqEiuaFre7XqJvXlIO4+6ckNr8EX9ovCHpTaQR6qzXfGcRbUL7
s+t6Lf3F3I2+RFLWoSFBQ2ibKiBWY6C5d95NCnr9QCKmQCCpppkMWfSbdF9DKkdM
rXQ4kYszBiMZqhKpMNIi84ZdFLtnO64CDRczZm+8LHdFASqmcfX3veXKFYv6h+uh
iB37m5a09KuGv3scwLmD9P5oFJVs3N/MKan8OoPbtYCJUAKz2c3oqztF6XqSL3hp
BiVLpGRsCeZdr90ww9KgLfcLMLVlbBili4f00tkZANl5gpnaF2yMaW9FNST31F3+
CEkaqciTF5CDqiVfXpIO+11jXdZXHlmtkRF5s0rlkhVH31JH0X2UbUfnb/8t6VCt
+KMxUh5uRDVWH9MN6Kp3yrbXsLHWiEEA/RjEd+2k4IMV77ItsCyJJCS+1wVBo/C8
xteDkNGAeGntTVj7u42mbR4P7nYp8EzKVZyOXmctlEN0L/p9Gaqa8qkfntpjvz2g
N3OgJOAyMoUsk255dtzugHk44UTXqQlndKM8uUBZjIdIxBSeIks8u9ifHaXx5iFz
6rLW+nNwjFax5Kre3pXtr80w0RoLMMqA1wdd1YNHkzmzWyGZFEnPDZynlVboee2R
hL3uLh5d3zf3PyG82i9uWfUMgjflV9MgJwpv8cExysMwxZYUepJXtP/G+EGA3mJt
WM93FTu7ie8prteHuAwRjN0i9kkwFoSNwkxQj9KH31xrE8YL0gT+7ZSTlpjFsM3a
6jBJQHwfau37T40GrUAUWVOUd2R+RTz/nQOhdT0uLBpbpQOdeyXzJQnHSUh0FR+f
M2E6N6Lq+g5JO2ujG0ygAVn6IaDhKg7/GyZehIuODKIvGD2ygXJ4ucoYrKcHfZyZ
taBDs14Q3/LiyadBqQGPMNuC9YRC+XPl4TqbWOwst9O953IIZ3ar6O+KNiCT5mJq
ptkSC6XAPjOCGE4+GJN4KqfaRFrTZZyiwRfQpB22GHjJR6Ls1lokMNwdWZclGH1Q
YN3hMbZHlmTXW6z7b4PUyGSoJkCZSls6SoMRD8RCw8Ec04Wk/T3Zelqye/3iL520
1b4AvxNNrQTTNRAu+yir174rj4Z0cW//BQdvpgVGI9u9qhH3PvUO/72r3O1h93O6
a4OqpNOGRt2GbfiKf2VO34svkEW+/w+y/lqDBrt3i6HfbfPzPei4qPL3MG1enmlw
7vYKY9PyEQrN9lEn8irCX2TJb26Tci4sUZfNpsswT3fdiKeqC6Ur5kPLgk6z+OI3
x9UjANKfCn2FERXaSGaO1ZOjxyemLDm0QK4eb9LLq+nbmbPCOR8RJyoKkGkXnpfQ
cPPZTkZKWHXerkgXjde2Zr9fa795137W526cy1EZoFrPex8Z4Ku+gKc5jAkakRHR
845MWyT0+gZUDIekF4hyv5cG1LxArmDhHUIVz5PIOc9W9HOACXCX4uNtmBqXZwZe
KWAodh3KUAyKqEAEjlmN8bpq6bIZpZcZK5Jl+9h3LrrgWpqcJUPOulS4BGzRJd27
VALw0TsGAEOUJVVd02yNVATLDVR+qKbtmAChpmWKcKp/XiGxXvHOrd8VJyh/jCcm
IB3v74ohzen53CEu8AkcmlJ7XPajjBcYRJzXZQoLeU7tmeSoMQ01VTjdyPX9BP9O
+znZRx63XXtKTklZDqQ0IntpHyF7ugwMi8JNqC9K2UM1vlqNJNc+WarMh+egSpBc
PAS+3yVUYH/qQtIqFmZ500YYyYlPunSmqawSe5sHsbGU1nVwOgLJdcUYNrNy4bBI
jCsS0YIk1PDJwULxcx5IlPYHyaeGyqf3pHX8HjK6hKIdrTHzDSDcRQ24hsteECoE
LOqi2ECD0nRqzBg8j9q+5vtBGxO3Ku5E2EYU4OGqh61BOL7myxMKKPjociwqMDbr
lzByqeVnKT2BRmBu7ryQaJ21cif2qOzJMdMvPZUMMXDsnbv00YcQRyiCckmVCMb3
5ugHpZ6MPhmS//YoDAcs9J6GdQcuNbMrEVRK1NeI23avzj5MXT5UkFap/naWl6Vy
eKfgr270dTpgfp/kKGlKB1nDgrz/6VHqttcju+JscpVLdeA25lwffeAasazeuY9o
+uBsWDri+FycJ5iK8LgJkQymxvoYNLbsJZeu4eBY6Qy4HoQCPl+fDHTYlGXhN0sQ
sSkPOjZuofeYFw26vUHVcKikKII65QOyAUJc1IJYEEKI24Xd6sp2GBsIfiqNAXpb
Zq4HnvWb+TB3ANrzKs9tnjj/og3yUR37Prm5ok3aIUCLyyPY3cr3/HWEMqt22Kvp
F4oPfmLs8oAxNGXvzwOKBYcxE+LsymEFCSscW0ZEkDQVlsONiSZDbMksFDvc1NOl
uvYdMFPvnpwj4FGc9rrcKBvwuFKs/xMnChdBWhS3lDquo6IcTONpVu9Ad2PxnFvs
q1tEzr5FV3TWYKi7ucNPbYkNg9CDEtop6fWu1kMFReChSqwy7rttNx4xF/xwsVmj
wvXyT7tB7z+BKee4FS8npQSCdJDV4wYjrPqcOc7auptneuPUzIN2dYd+EXeIw34T
l8DOPcX9tRSFuGn64yaE0IXNM+NlcMeAswgZFQRPQtztigL4xgx96S1kGqU+Bltj
VpQ+Balfw24i9n7DmMJ6YrizS3raBejmgYenR2cCBQKcxLACfb47pg+MNCGBDWJC
Kh3+D6FHDmSnYUf+kYmTqq6Ed/yRLDjKC6Ub3ZetMijM9Gj9IzKNW1mzG8QAzviq
UHXruys2Pd6F2z3Ny7xD9pSK3LRgmbT43fkmb/NJmeosc6Qx6gVQEndq9UUk8QGT
jht03tIMpvTLoretHhmC9rYOc2TGtMuMAqyoi+etSRWuzGfcXJug9qw8DdmVC5Jj
X8jjLYvNIelFgu8qg/C9GPI6u/+AQFJApJPz9wFCPfseqmG+XCvXqaU0YIRdmdn1
Fdk4zNIRaJidLvW1HZMznEoopgn0UNfFsW7KH0MgIMZ1jeLaS8VSzBJBjpFuUkut
nCfmZEJMjc8a8EO+SnzbKoShRPf778FZOgk15apT8qpTOq/+3Dno40JAYdL3tfGh
6DQSZZ4esB36kjHBtZ6/ec2TCFd0/9SwtK6z59ZLRX6k8toWPo97gXi077j/i7Yd
nSP9mUDGtjw47XhgiP66p3uJ5opfcZsl3qw4clUd0HWQDjp3XU1P2I/ONfIEqBUI
h39ZG5Y9n/Mk13K+yqjamncY6Nvcsq59XCWqkO3sIV+c/0VhNEZa01GGet2uldjL
osfJi1u7RPL0pwpdLKQEavOnV3JxL2tW79x6vmKBv7QOhupuVMhhJhCu+vmA41eZ
4FHv8QjuFwSEunyRyh7v+DU+2UwOFyUPk+TzCZz4hTQngdI8uQNLHqCX/L9UNKPt
+oHsD3h2m+Qy4xnaSY2Pf8GjDlC4WRmpQ08RqcmIVLJS92hDXDqXeBMVU5CthHcR
20yx9omUjIkvTHIi6wSomg00O/P+lvYUWLbp7+VNuzoAhgHc+6iTjgNHhpKrWS59
z3ln4RZV2Msl4mOOtklB9CB9MaYdWSjCdpNmLh0Cp+9+tfOS7nk9WmHRtJsjV0LW
yQHepBXIvgOSETjTbreQUEd8Z/CQscqbnKeBqFLz1ARcWS9aGC3gWq9D3oi+q1CP
gBBE5NQfi+nfjAa5jeVPvNnO/4I20PbpLoGhod8f2OmgiwtGTDzB+bZvq2WVdg7z
B5Mj1SwvoQ/bSJgjYcA40LcLKIFrIqa8YViD36GETYpLq94xvMrM/Irnk+ODBIvZ
PL9xv6hOjZl2wgqrEOXyTpQ5+dkxN9pDPvX7rQrB03ElLu839dzVgR4rHQ360KDx
pB0WmmjW7/fI78l1fgxO8QM0KI9B5iO3zJiyAVhvs0eUqiX2PrUINqAfHD4kB4g7
igejgeVY5zt4Nh4Qg9aenWZu5hTl0KNZO97vK+Re00ZNRFyhKtGRmU3lC990xBPU
eSWMP6rtOIUuJKO1YsRkovRL0WK+GkbnDvGPcVA3xSFdkXRh7Dzt1qwlU/ZAz+Po
ECMTAgADSbNqWgn8rlZrH5t3kKUUbizOTbHeHsNqYIKIQUBAN5dHy6fJtXGIMQj/
PFRZFGzqci0HQAendzEyLQAbnR20V+fBm/YZZfBdrVHoxcZKqJsPmR8AXAxPmrp1
M1vue5yR/YPw6PxxevGPwXum1Z/tZjHR5SKC5uI9DVDJ6Hx+KOuCWEERoot91k4g
DoeUB8q7Z0EZLeEVOUdHNoQiEEXdpcO8gwc54h6SOItNpuGvqKgxIQAB2khgIDWW
AlINlw6qLIuQYUq54o4EO7zlb1iWRQSgX6/TC0dbMBvEt2V6bZn1e6w2/fXvXP6c
ofG1JUbOOZStWDZ5uYy49hTnpRVB1meXR2F2hctC2oyMEr8lfqgr22kYkidjy9Xe
PdQR30DkZnLFEA+O43wG/uR9pxqGis6PnLjpoI0UttGegA7znYxv01fLdZxgH3ZP
bigm9xLuUokQO1K9nigzbvEOLdv/Pd3gNoyyqPiXMYSxDlKSWDpdXSaTqPxd+3ga
x0zsHrD22k1knTAkHOf19/4cRyoXSfcf0lzl5WK05Yo7cPaTM0ClH02BtHuJ40A5
anwx+vk9vhoeziK44+oOVsrYUfE6BgtaQW2XfDOQls1kQmPizroRLcig6wZEYcFt
uDzDjyh4VfMl4jPihBFI7gPCocrrOtUrz5+TWjEIc61wFLm2BDGv7zHcxd6nMVRt
7uiEuSra0/4LtY1xm3QOcAB50g7UuA7gc1CqdavPj17o+ftK01jGBzt9iciovh63
vlCO8bXojgMkLJhmFXYEKJPp7NDdkZWd/owckUQGgwXCPTok1Uz8TFwJBZ9ikGOl
dU6hocijxixFGZQaqfde2AQV84ysY8RkAR80v0YUAUwAM3bOoUR/K0IwYos+wzis
UOzclvMK3AlkM+LyPkVFx0WcdzZD5U9Xau1+Xt/jUwkfveEpEq3dj80S427POqtb
AxAEi/X5N5XpLD4sVqGXWu4Wb24Zf9vsPzKcpeI0fi+5uJpTV0WT++ymr3fkcD9y
pkOo6j68f84uwGmQItv9yDiJpiyp4aOsZiG5p3RknaW/cRn5UGuXrR3a9mzX2WlF
fUWNdPVuwc+Cg4UP042NBAjiS4N8oF1oRBtI1hJwv3HqUpyn/6a+7gi674RcQ28I
1TVYAradx0uWxvRpoyjxSmUoQEmbijZ5VyYKebkJOhU3tjusiZ5Mzj2oWM6X3hU3
57DahHjYjisSARPGiLRGDUI1wvAy8AUgS2GNbmfJ2qty+LnsW5WUMvlkaiBU1Eg8
AFFJvhu+RgIWM6y6QSST4cCT+FS/sEOKf0c4hqtpEEssmbugtlJg7RvbjBxCtpwU
L43o28AvJpgSFLpgMvOJbsob5+qaP+dwEB4niLos7X1X67kb2151gMBGzySrQXEe
iyADR7lfQOctCO/yCsQAVrGIQoYOlV/AHoN58c0C3S8xJu9TFkHM8o+JmP7d/XD6
kWXwB4iHTiUB6JMPDzwm2Nwrybr9ed6bIUnZr9l+cbSnaaA8swEZT3//mq0V7rQ5
FFqJIVF0XVFrWVvESHHoELEFOD6eSlKQfGIdMCafL9/qK2wzdft0gyPcPrG+xtTY
F741xyllDPcU9t4Com1CZZqmr9I2s1+PJUs3Xkw0kJVzPfK6tMVTrEhbDxAfvrUD
QG9gqJr5plkTXdP1GnM5qby76yfMtw+0Dybi/1xSt2B94jEQrxAHkmQYfVILalsH
Zu46HzXlG5I9D+QswMnk270TBQbdtIKZ+t5EpP9qK6dCQMTDoLnygzPzk720wKhO
Xw106kGerGOF9Ds+ZdBea2jpWEBQ0pvqTJwQmktQsOcpeYz7F9A+caNSag+ZHIAU
NmBAg8QKOH6oGTz03TH0LOCisS6YD8Xq6+aXsbwoqgBmdQshSg+L3Y6/7LEEERhh
CeJ4yOsf+PfRWx+E/lW/ucRrZQsSIhAi1wrHCkXOIfksNKHTwSPLoexFAGc1YPSH
OCC6dDZK70qEaEkvKrjkd4B/DA3QUBaQWoTmUoThIh9szw/ZmSItvqYHtQpZAOm+
I7No3RNGsiOztiCUpJjJ5NauR94vYeC84qL0h7QnW1XSeTdYNn48Y7RD4giILOix
g0GEGSWJ6k8S/0n/OkeqWvMpUEE+KI5Q9dnPpzNOoUdUphFZX1okkMVP0csJ54dz
wj7E4QoEn92O/gbMlM12oTaVBk5fiO4dtD7WBu/E0ExyLgHMT08I6M0hKj3bIku5
jAxPk41IEC+wTEoYNWMSovuNbDbF8DXZPAc+tVgbctA44At5yXnvkliFu77N+i9h
uvSQJf5iN2W8kY/TviKKKm3ei+seo64ckBWlhoj+uu9FCB0HipHbsX2Y+icvT2Ix
hvqzrsqhU38Xmeq+37Ei/uTb+ltc8sZ/Cl/7F20B/dPKCeamp0S0B313euz8VvKW
SQtbDvmJv7QU0z1ppUlwve2HR0lQ2+bTNuOs70R8INcCn2AG859VX10y5n1XkCOh
imZYzs4CDI03Dx5Yr9w0ZdnjIaMqgm11J6oluXubjThaA4XF85qWB75YwHQlMqqn
OMgXfElJnkIWsW0EDQ/jVq+aEVr4g1GjEFoyb/PoMqkF1oUZoy4JqeA47yesWH9v
PsMOokZbdcmxnLMk+/Fp/L5kQ5+NyqwhLFZukpvQkAGSTOuTrb1HEz3PlJm2/oy+
jzLawYg6f+zBqFUWuCDn0oaQtFO/6+z7ff4R+btJHpEfyK7OFcEjMcUdrqLDazg+
KEnRUpz64vBG3eFaOFvmeFWYvAeMAmFHxFDGf6Rm106O1eAQwHdLOURfKK+V+nwy
4dTDr9kZTAFWzQii2VM+1py51mEtA/QBfNW4terPbqtgV0BczYDGUW5vZVrbUrML
7po3zhY1YBJHnMI2TyzboMdvV0inFUDJHPiO0VmUyLXsAkFwQsN+ASnVFT9xMzbc
TYAmMGOeKgALBvh2ZinIRxls3g/8DABo/3S3bb8kzPHeh5QLK5IpdZbTm+sWTIu8
Wk/RvWqju4ikoZGsFSjHKtE9RlBTkbsqx9laastaofrBocLl94Ivk7t/vo/Mo6dR
qT4oO30p+uEfNRExbd3F58DLtiBoW9+uXTPGHBFE1nVHWIZcq+2VtxGSDrBn3iAg
QIeThtNsy8mnG2kTOc5SZYaS3Z4U4uoxylfjVOOG+xwPuZC61VEp85MohEylnVkv
pX7ftbpCZ1DIBYkLIVkuZT2K2aatCXJCTnxtc2rsuFngoju+GKweyzhh/+dMxpl2
G9nWcNThLtO9VzRaYm3kvzTgN555F4NQ+YQ/hzzdrATjuhsV00/aVWQp2lvLf3hD
/oEIN9IUaMWI5BSCRS0Stmki1XsOqtmnnwVcBeLNzai8gjwcdcNGpcLTYIVFZWpA
BL2HthkZNPwQYA7xI0laoIWgNwDaBafAaW5frRDacg4nMmAtIJS8LCIOiFv1BuGW
+CI03WszzEDAH+o97dRu8KkySoVNRy0Xs/TUhgbI3/S+qzH3TGqbpMipxOBfrKGP
myFqGRpB3rU6p3nwooZVvdOfa0lGgBBsNPz739neY0pFy5AXm7wDydn7UddTb5qs
YTrihdLyLNAkOexuD5alRpMxIqNii6tW7jZ89kwIsYmT8cwl7xQYT3j76fPM9yj1
57eyU19rTZI6QXTHibrQLHY76VDsDV34GcktOAiDY3Q96syBF1LyFJOtL9LBmMh1
sRAsY0Ff87e/HPWksULYItnexcvIvgBBUu+NSMtFP73LicA47T9xSGDLOdOUgylF
OcygF7S4fj0lLXKg3arlNsvat3ZMk4lFzays5emhK1eL8vFIDzofRpZ4r/mVbKnZ
3AyTujtJjjvdb8imjvLNP7osSuHzf40FDKlAPkf8uOzxXn6cazkAJk4FMC8kljpb
rpGJegpg1ec3aSK2TwmHiRKkgxxcVXrABFJnCH+XI2mUc+BtwyfW+CaxGU1pFIY/
M9rfNvAeZbim9bEKLCNbsdreEcRfrGNcBTVQgz/grq+RV43uStqS3tOuNJWIfqoQ
hLLPQp8c+dP7TMgkvhg+yxV4w9Z04eXwoKxiAsve5NMAfpQYSi2Pov0SalmkbJ3O
GNOPXbgFAgriGuZ2/yp0ELRmJTlGnzeL8mdSi5n5wzoVhHbrPvpR6O/ujhgXsOGC
EezObX7e+EP9gKRQ6SYyHEYxy/8LyM14SbD2fEiiQFEEG+vX07A3D2FSUVeEkP3f
o3Ii5d93bpCvcrZCLjegFYu6lyvTxXw4hcSltcM4XfFZF3nWUQu2N/teypZuvzWx
70qoGtPg/e2t/gby1mJidrB+uEKhmn1ku7R4tdxhYvT2DSaqvgiGmi3bGgicIJWd
247BvJH3Zd0mHSfGK/woQK/W29aIFdRZO8WYPJcAV4qIE58LVpBN4Su3lNb2QsHI
B3YNZo99kJqElmloPCkSKVHumAFy5sPTYp14MHX9VIbuwnKvvhKtz3lUYY6eszmA
qnr3j7uXRBn3IDiwvcR4SHwvSpQrcXjMiQwdY0FXYGnSdq3pyAyonY6coaR81QVx
vwpresNvUvTcgWWcTXqYiGNAGpEfywyH2FVd77RzTkum/0U+4oFZagMQchF+HusH
pPEbSlCzWJtnQYQE4v6vZMEZajTfY7G1LmTxRluJ5MTzmVvRXwDq4y9DYCgqI6nH
mlgA6NXZpaT/TB6//5PdNMEeWu997NlSSIVlxcVULZEP2X/iN5OSngmjfwWXrRII
OFbBxkRPuNbuL8PNwEXDv68ryc7zeOI3ZCEfhsPrhj96x9D6ngeIxc9MQ9ryt9Sv
mYZjAW5alFyMFBfnUsQwh7L0wxqFFxCDrpm19BJBtHb5JJYRhC4eFSXSMjZYQZky
67w9pidkjahDNfocILkAEoeWA4ZTm89XpB0eYquc+RZsGx+epmYMQoYiFR0MllXl
LcJf2qG4VrvaFf8hugUStkUyvSTPB9iER0a2CgFTrdWwGE5CcRm2Jior6vpTcbeB
8h9eQKu6h/JSKfC8PcPTOh3MIyWZFnLO8J/FqX1H4/ESw2azBxeI02sVhSkBFN+y
SP1hYm0IIdWHyvg7NRseXEt1SBB1Boav4ZGBZDb14SAuhhcGB8NQ/6U6rKF8BAnc
/lD77ntavW2+a2rC27Jvk/vUq194yoNjarVKpAKlW5mNZV51ShhLO1MJvvzQNCqi
qAxHinMgxEbEXSHxdZpoPYzIVU2T3L/c5paSs6UUKfWh/ZDUcX7FC/GCOrXfwAON
kd09snJeh4mgyUolArLndSffn1bmsMUUrKPJqDynqfKQKx4PCne2gowKzYatU5sd
J1BH3U6saumxPDPlS/shZHKa3ENSpoGvrpY7z2+MAJHKmPw3Xodfwd+5cBE2TZs8
zSY8XZ5Jvog+vEm2cR5od/3jqKzIFvZZes12nc1F8fhbsQrjSXJhqmIORSvkNPPu
sabMuNiwpWZ7w/vdHYbb6g3FHxTmvbm0TxAeDHvWRxNTxdiir47LTWMH270kQHa1
0biLSKBQXtW3YSMJJA0SPNtdK+YiHnrqDtv1LyT93alw4eRKNd+hQmZulRjw7cyA
1qkpa8ug5zjsx6m/QltOPW4+eQ3lTPmJ0b/+ScW7muKZ2VImDavSyTXwWS5MCE+8
6yor/Z1u4f2q7vcLfx+INqj+eeF48UBJ2z4evQx8mVEnQRp5plOlKfa4XElDV8YG
qNwkm2H1skza4KwAlxUKO83Z4BnOXfxZNF5OzroZknHPg+xgCqnug1MW2ITey7jR
MbJKb2aFLr/oiCoomaiQ3/sTJ3Up27GykeZWdOjkVR+fjeqNsds0yiwplHaQyDRe
9CBYtNvgkI4SUNdGGtofF1u9J1XYlCp9s9fKv1eWpSHvGNxDECqM8pG8WKZtv2u4
qT5EpNJu3P2eCndAiFw1Hp+HRc5hpcmE6wp6wb6IACBW+MalEVH7cD+by9ioBdLj
9YG0yt0Fb0xa9XMtYAGCp2igy8sO8VMkYyvzZNzZqsWHGCNLeehrnNx5r9h3lj/k
MqKMV8cIGw/QwkTps8C+Wo2SxI/q/lQurfVrQegkyiUNO8zKpiCVuCx+LdNmzkfd
a2Rq10U+xrfR1Cpci869r9s7Rw3kFu0iLEeBrY/qSfvce0CxqKv9o/2B0wJZEJ8T
epA79dtUrrLneGSbwDQ0/qusQldj7NgM6Nqg+xfP/j2J21Cgqjeku/9eTMwihCiZ
BU38IHvAlmWIkxvJMi+R6wLh5NL8ajqyMvqDY+YPzZt3vqC2U1Ea6srobPTcYgOB
fPZ1fI62Kwwthm3zicF4bLGEcUaSo8uMEeft9Niz8LypiNGBl0v4vRgLcgEy4ayU
eYp304vx8qt342eM/J1KU73JhiU9NQhXhHM8h4GHXWR/hWBA19wG6cXV29jnmpm2
IwzuwiOqajX8S5rLUnasgqxWhACIh5N0N9vq842AsnH71ipna+pQhPlsNR9jTHXm
jJ+QCLoIxgf5yOWUv8+sw4AcH9mqMT5wB5xgS3o9PhFDI3Nr9ZkGG5cglNfH8gXA
AxplHXrkNHrqgZ7zA8595gz1fJGwMAymjQrScsbVlP1/OoP+6uQX/zHAUwE1Ivc+
fWuLo2+g4lphijnmst7NCP6hXDubZz4lOHmstk0LLV2Fj3sw3Bgcp8dJKKQheVvT
lDewMF9QUUa+nOFlaEsHUN0q6m50BTiqIURok4dHW3tzF1g6yBtTGWPUZrIWVX3w
92Q3CtvMQP1SRgbErXOAunfHo0PLXQg6lGBtXleKBhcisL66FLS5E/e55pDy+Ljf
QY26It5Cs1i04DE0Al7o/Se8zsM/pDkWKBTQB7rXMJoJeMqxwmYMVPKRaYBTXfMR
AkstPAj7VNBVvs+uaNVsJteWmPTJR83MWkZGOtyCy9pjOZCc7+y03YClmMI/wWYS
RmaW5VGy+R9aq3ZgBXG+VC+RQXRKuk2FA6UjnsATjHDIDYl7n94LIEHRhLpRpmyP
4qnNU7LbglW5iTraAwPwZE2kVaKLrsMJPlCbn5idWzHoWH6nDi4C2ra3iX/TWV9c
t4XPZ4//y0RLLqgn91crfVKup0Q0nUks/Ehg7KuVKuM7ztrR3wBQINAVUXAWEFbw
HNlSgQTVRyRw4UDHkeE9tPXcQHBLkFmjzJ9UQfciniXcQgvVVvzTihpa62ITXVi2
omSn7KOSCKqcDjdXb3kDdj0emQOvTY/E1x02t7/m7+fVvxc956Hr5piy4FscDFpI
sgjz7iEjAFp3+hn6jF/dD7b6M+CEPqFGQ1XXT+W3HqpkrmTFraaQx97zVOzT4gra
ski0emG5/qiR0nUy+Bcpr0qJkQuXbZeepFN9KOD9HhvF2FQN69FFb+0CMdEuukMc
rUi3SkK1rVNDlzHsTGI2zWppO22o0+hQYrF9WagCSsAL1hJQDYdXnT/d9rJS0Elh
yNF6GcWNOFs3U7X3/S1Zol4GHk4FEdaDqHCPLv3dyIPjSyvapx6unu9j307Rs0Kb
ETIgZvbQ/txKMwVL2MKG6GCUXdcadnmAr0e9W0kwQf9kkuF4oNQCv7iX0CxmAj8r
XgDe6K/se2WRwx+PHP3TatmLrBh62vPMOTe9Bmrbo0ee+NjjFaqw5B3XHDomLc5v
OOBwStW5aifWTuvpaUpbA0fagCXaUYcvod1srMdnX/CKUn7rrd5FNihkZePItGxU
B/0wjxeDVzCT3GTtjOKHcdsPkF5FPZBWU+Ti0u4hPzmSkKgayd5eQvU3Xwmpa9LE
w3LE/6ZOnLP/IimakjCBdvTm6sZ9qwnNyyijfWfenAmBSCoIpGXQMyLI4YDIgjIq
c2yB7hO2Czyils+awgSURy6/XAfGei8mc7uPNJ1aYvXrnv7XJWYc8PjH5BpOXRSr
rDL6bqXIeb5n3IpbhjBv1lXSWlUEh0+u4Os7nbcikxQ8a8SNrmXLH9sc76cA8NKg
JmqQM1cfvnBrotZnYvUyxQje/NPQTP+J7FrUZz+KpCwysfwxGvqrrki5Ea9rtXww
7qrSLs406j1jjVZFFvCIPSRnuUZwF+Pw2KDQ2tQVWKMVuV6E2Cr8ibwz63T853Su
iiPFeQKHWCu56Mft6eCd5D9U+WKlChAqmS5MmcQrEKjpa3gSbQUUMGCYorDTpmfi
mnakExEBAL+PWXC7AiRtIEmEQqyScvNYZFlP6HTrn5Iq0JuAOoGBxhSKuyaOj7OU
e5hQHCpQt3ecGFVxsNmEzpt2ltX+4k/htjJ6JQpXT0si4zx0YIL2lUsnFm/xL8/n
CbOGyOkhDkFbhgmpjcnqkEgYIOLlk7hvnZePAcnEn/yjRuPwnfkXBF/thJQ4nJ6Z
dPYQbJauK8vtsFVvqYw/PXxuyftiOIPX5WVeCalff3vqC99Iky+DZUn+XppOtpN2
H1hqpRkaVD/84uWIViR4X+VH+/xFv3PGHITFnbIIEqA2jkTLDDATJde+VQHt6lRS
AuxXDB2SqFzcZWvN246ox2tPTu39KyT9KoIPvZrs+rlP6evfjYe91zg0S+arJ97S
6fOLF9rNScWErE0ssRszvYpvtBYY7qrzLvsPhO6yZXskPylHMxMV6UvDhiJ4aO2l
tzAoKwTE/RBVsB8+VGh+vhczUg1SGht99vNYyqp2hqQjSggJ8pJ/lvlmEYPROkFb
fdPl2A9ZYFiHJOTl7FSoipNugjpg9e9+ua8AHoyM7B12Q5Xo0lMYj4dOSc01Zy11
ujuFOzBzdadcUc2PDobRsLicd4phd5zDw28lk5ztutRGX3LzAcRkKpe6jEDwwEIc
h5ccUzpDoue5DKgcetvY0uMjFozOge6Y8bwyC7c4X0y5Qy/DIIUz9BvdJz50kScc
3UmBv8UB+Jc68sNFLZw3ZW8hNw+P6f9EaUPGJey7WQOhSFWyTSjClezGembNxNgK
C41cREbJZShQO+rEjK7VJorJgUHg9sZRffighr8DF4yIDxBE7gY6rruT4TRLoOPg
hBwBNBjgKj7fH3NHYNG1gZaHjvfw2lkVTqwudYcqFctFXD7zaxao5g8u6mV0cn8K
rmEaN8AS68qtjqa7vQa3+rpOEYgj1vm2kbvRnrB7zwlXEXMB1KHmv8Ms0ZwOxcb/
ABCQaEZYYz9sBOL1rdx2TKzmXpSPEhx64QosIO7ZBRjFsVHBD1o6ZLE7AcrM50ka
8h2WyqeGROOvEYxzyOgMDOQ0Cw78FqHG0YaniXvipSqO9xMSe+Zpgo1NAcnMrglJ
1AsIaq0LvlxVBTjPITvDfah3//FIOdmCCM+sgukZBPQ4UdY/bGNZbrDzqNnNukb+
WTQVIjoTT6+wAEfu6PJ4fH+ku5je6I7K8HpKIpDGgjunYWpnituF55FOWteW6s9F
mOdWaYqiMcw6Fjts/GrgnCk1tKi5661Q00qDPJhUVokCNWlCSUcYlxvHXAp/vEPk
4ReSMh1Y9OVB/c3rBcbIc9MqzyX5P5SjX/TG9Hy6mePf/sw0hvZ4khLKfZFtI4XS
bMtZ5Z+PhEkGoyf0/+A7wFpNeyHsvMjDKVIh413XENczOlUoJCc6zpgo2VDXFbSU
CjUGGudKxXiAFtFRARj4CguSyMWKCs0l9zbIlWEiLhHThg2UUHMylzaWTM+maf9g
FxsVnEok+celjmf2Y+767A7/xzOnwc6/DKIT2KqkkYzzeS+trOdk3Wl2yOs3na+s
zC3Sa7cBmQEA+yf5zcjeisq1DxGVbQxu2R3Zy70vLbVeuP1GKdzYCbUevLMygxqk
I5T4+W1qBqm6r8gUHyvGdAJTPALUkM5a7vda16CIW0LCHGSJe8rm5hToqXa04VxT
cPP7fM9cZgyvQtwr5F3F1dTm8XALYSydYXe8UhuzBU5upBpfi/359tHm/dNGzNWH
Q0NTMR9cQTEFVDLNqnmQXaP7iBEVHZf/d8bKE1V3yE0HEtIE/RHUjQYFSDTfu7AG
/WmVPIexIAKsof60OC5UGJjgWJ3OsSdkbh+viU1YvIAfN4teXVd6+1doPFjmm1Cv
ENBBcXa0y+piZaEEvcJVkcC5o7yuHHs0jQnvGl/86B1oEqsYNGtjKfgvdCZhilVl
n+unzgYJxIbNMCDmBhlPr8u4JNFJJxCLsvcJI+X29uSU33CkJcNQKDpCM8nQz5Z3
SuP/kqoVq5/Sy28v+OA2qKVJ3ybmFvnHZnAud26aTJOeUev3mX6GgfR7qrpL9AdW
oJMbH9pPyqj3WF3VEciSiyIT1PttDVpvwoVxpcbwm3HSRQ2joEySc7uFpDKTDHPs
KWqjjcE70FfBgq06aADTaRpQHO0YhrcjmRIwVOWFbhpwuAEx04XtyTsIi+z2LHPi
FaKA43SXhbeHmAX6IqgYhP8w5mkdtlwuVAKYeOSuPfLjg/iKuyfYmtEIL0dyZUvu
+dL6ZQy6VY6txrzj5r0lZWZUMQGRvFvke0K/PrOvMwLuPplF/OowTygoAKcCskOj
ETAQnC7eLqzoBq7nf1AX4GC7rNT/brveGlU5uQt27V2/l2xhL9Wmsc0l81LaOMFv
yHGmVdXQ8oEB8m52T7DHXwRGv4NumsS7suuAgWrb1a+LLn2EwrdVlCoE+TnS8Cb0
Be5z/wZGIPwmDRJmDGGOJlrd38zVkLbYxlTCM84UnaTUCQSnWq1SQU29El4WiHz0
CFisgaU6M8FdD1Z4XB1m0QcRc9ylZlPvRWB8mzABBkFgth5jQw0Pk2GiJWpCIHKD
iUJw/vUl9ckAAzqPJa5+Tf0fZlo/V6SD3Tu1SwIM7zohuhSebVDpU9yQLERrIvZG
HeEq0z/d4UMnvuMdoixQHZs43KEd/mknP27zL6ivesltuFGU9vsr0y5UxRXkz4KI
fUF4OQSG2op2L5rhsvOBkoLPkug65pVEOEryzW0lgOrhlfmH8xh+aMvdSgOAYblU
oXjA2GVRji4jBYqduGMMHYCKRy7/q9FbZP0nOC1FSIgMwW+wH9694lLr+d+DDrta
COd+4EuVpBvGC/+jdQoyG+w1NNWCwthjS45CCmUbD9eJc+yaeQ/g+x57VBgpmNzt
YoclNNv0h8lHVJ3g9hHO7BN4rT3SuGLVNm4ZLsSDJw+h6r0GRb+DMW0LgJ2V9qly
JGZWPfoYJxaCiV/xzdDAT8v5tZa9vRlEUf1e6Sk1PllKfzCOX+iYDYO1l4bKn9Xf
mhLr/5ObqDL9clxWG7F1C69fQU3CKkRcaSdh9uz+kR4YUhJWnYIY37MXyQrbE2ZE
ctVZE9mizAuHRHdHP2VqE6u7ovyHdpSyYGGmML5gtNGnH7JoPziE7TL9BOrl0Aj5
HMYUxEbx2jil/Z+abdiRz4QCcDlOeJUGRKj2evD4ODo7mwozegQsBoPlLWqHxp6R
lhOa4n2b0+Q0mu/H3TUJVgc7WKg03wIUetod+GRtUdsS0Eb2SE+uIvXOoBLzxpYY
IHqJ0oWLAfkVZAnt2SFpMJwTVR6yvZNJRpxWzyL8zNTONbjETp5VN8od4eyWEn+Z
dSuL8ZGMygRGNK/QreHX6eBIcY8rS6ioTVYKNiACD/BKgrdHewChPtXzt8sVe1ov
40tl9kvYXJzYFhk7D6nDVSVtt8jWrfrKL/OOfzs2iJQplHyHzXRL3GY5ClSVtk+u
hw+pOzjEqvVz8fMGeIj7rrZV48buvj3yM629K+kqJgpvRfj6xHka3EFi6UswGFdi
eZ2duZufq1NqmTj5+lnek6sM0hDdli5OAT7ci/dmEy0WkuznrYrBhB+rydFVWpFy
cbCoTPRlCvQJ/reNFqJsXFisVyOhyp2gRGcB6JFBIsrSKsOnYG4T+DcE8GuAy/Fa
/XpSQmFpL6QrPP9VgBGpLGuj9Xg98oSsFpOJCh0RZOc6XqAPse1DBIeoLYiNUIdd
yMehcOtGDj0kP2k7Wa54iHInhFrD8Db3upDro+XrSrRyTMddgZItJp6hw6/e6yyD
ZyiYpkuZHYLIfGr/iVkTYIq0DZ4khD7kpLwWJ6gK0BDKpC2w9bQH1/SvZsHC5ntM
94pkfcnWHVxhS4cBLSJLEw4vD5vsY+DZza7MyW+R/V7rIpChk7ruyMemJ6BCNLox
PBD0Kxqve6ALoZJKSWD8D2g01s3QnIfwrZgmbLKld3gCeYIXCBaqzz1oev5fc9/Q
Jwt72uNM+ORTSd07AQLR2TZKkdAf9/+MFKStH01WUTDFXtxddi1DiiPQ00y+Bbqq
gBzs/hZ3iKMj7XY4jEs5ySk4GfILHYnXSKIvQvaRoboSoAeyYuioXqL+VCvi3p/I
PT6Fa8OCJvRP0pOnozJrwH7kKszql0sIyTB1QipbnYrAr11m1z4l5tpzTVcGip3J
jO4V2ztqiHG2QSh9gzQyYX5DAImE54wxPwKsYiFFZxVMpYfuDak/Ls2A2b5NajtR
QkbdIQuel0PG1GDZrvvmWWmW3eo7qCFCoL+nGmST67q8UmOGp+1Trz4r8lATjARD
+ZhS7hHev1LHPuX5Pz+IygyN/hnjooQ2Mgy9em2uN3BUDgikVslb+b8vq+UkhdL0
so6XFo4OO9tHrpWcXu2H6NncfhhOOmkCcrtj0lDVOmG04jEfItO/CntCi3bLHpih
bBf3n1pHiJYC+oA6FNJLH3EjhiULAV0jHLhvTz/2/XsuLX/YjjrXDD+maDXeUiqo
Mp+M3vC0EJ6pAvAhqT0oQ9h4Z7Bgmt9ASSrnhIhoM64o0KBlnODPIOnfXJNrXddO
4vDl0q/+8ngsNQ57SCovmNkGKDTBCmxqVkGTkYzB82nrQ8ijK068pfxjqVNDBuH0
v1l8xLz7NNgwHGk+5MQdeX+/mAsi+f4vUFJNen7zpAsur1/JQKGbtgl5456CPm5e
Y5IUYLPMnI5widLR56dgEsEa6cBawmii5TlrYZvRmuBrZDrvSiM+TSw//76FjUQM
6ck5it/mWXKtGBbgmoabmXp59FjwAY5h4+g+3jsF7VvU04H2/K0z2QsVZLU7TLhW
txz5HysDhti374rRPMcVvcb6VYpAIZzv/mOxNNsZJUsa817I9wZgQ5g+BTCUEX6+
OVM1cq426FOM/H5Jb5igOLvXxv1fKdlqQuqyo90KTjz1wtgaxh17FJTOsJ0xJ21N
xPg+Kg0LD/is/jaKkfTbBWnZyy9dPwRLunMpobsp4AoP5dKHdIXUsdi41MlrEKy4
/XNlT/IZU/Gad2Sr4ZN7qP8UWpG0i0zainue4JHQ5pPfE4hlsRsZOz3p01Jr81Fm
n8aG4lGuLfXFbixHH/4kgqfXW+fWMK8pWzMacQ2sRl7WhHuheuXE9K5KZvNOPt8d
J/PnKFz3+JD4FZ9k86uPjtvNVFVIVcX5GmgVyXG7izKoIormw0DtI+E/93W+dI32
2OPdKghwvGya9YVmSX1u3qU20twe9Z0ssiqfWTHlyiGElzIV6DZc7dS/de79sU8b
JE0KNR+epaha2ERzq5ivMx3dk6tyXh1XbpzGmGtdpQ9nYk4L1ADY7J4kvezOTNGk
TOLhCUkeA6WFNWuUV6rXQDj6Qn6WcigY/zjGBfcwhx3RWJsXySOHxcaQiTsoFqxl
07YD4SxqzyaFnIIieK6wFc/eFIvuqIWJXVLGM6TjIcRUSLtq70LVqRtEuqKiN6EU
hAAyzhNR00ctfKN0lBvJYcpMM26/5MxjYh8tuFvfmmRtD+tETXVMnFr78hws4MJV
uo0wgsXwy+N4c6D7xZTmU6dIwGKdbYxymYZmE/L5G3EIKZRvzSWNz9ym48vHr/Tg
0kb3vZpWLrMYAWepGkac5Xi+3FZU0p4w6NuaZ9m6JNFh6Rv+LYOj8jn2XDkLF3AW
XMbnbU8a8uGJ1CG41j8be3wY5yB6XEMKWSs4wV0GSAABp48gP+sdGAdwr6BCqJUu
oSWiczjZA1eHhXEZ2ao9C+IwJH3SOZ6oUCWVcrsT7nNBJ4Usl0qzUHX5eaQ1hvvl
Amskf2Axl724Gnb5IQd3ywGQEFfG0+ByjNki05vpEcFF2hylhGaq8kE0t/ZWaOmr
KEUCxJJsdF+W6a8EZgU6RvsAiI3C9fs7jzLDm5LjcwJQH8ZlnTduWHKuEzZQpP/A
8/lZWX4R2jdm5yvKtO4uOUE2DsWTDbUj96kH/n2g8B+CIdKfGxfa0MmJ4qN5hcLm
Dbn20LK91P4B/mz8ohPBiNDOWSYpAmM1ug8ZKvJbNT3QKu56mPx70M3grYNYcnXr
cazZTfORdek+o1WaYS2MZaEiBE7+WjNYgXq8ZVa3wH9epFbEvHDgHPMM1SxDXXl1
aBzR4wO9UtPy+y6NTfFZXRCQdBJhnx3DUctKXiK2NOAzNXIDphwOzLHvkyCDN5Kh
ENnMBl1JUM+f7JJbZO27/4xRDFPjY3gIiqEcNKr1in5rCRqF4Cdx+4n9HxXoK/hy
ORbqoS2K1JI2+uiQLRO5Bm40zABOdN6Mn9dT30RrrwN9hT7kNXFj9YGCrk67b7pB
iav4feEReSYAcMMfXhfh+T1ZUrCoskfeWTtMMgYeYMiStog+bHDFPtAHLnPcgYiI
u0WXI1Ahx+udUxslNV6dzVRDtiarROLPXZWXAqPD0I1R7LENO6vh1h7K4HUy72IA
fvI0fHI7SsHqgWFfaIh9p4oJu5mPIv7x3MmvQ2vqXa8ogU0fse06FJ7VRQYcqteC
rQs5Zj+Y45pnoUYmUDZSbI6VVW0G6n4ynmpyUJo0x6O+HioHOk4KQ+pdzwsPuZ7a
vS7W/L6q1hrSuxGgKDo+2gyFN5Rdee3OEz+3DvQlHVU53CAyQgPb5YW1BczTwdAU
448vu7JtyUWs5j8Zq0gR5OYdUGKcqjb+RblFM6JCtXqyQS91JWy6lbASHUSzWMM+
bvYFyaauhRU4c92ppJQ05iMywWhNujduoeMYeyr3eG3EvGmEwW7bW+b2s7uOKiJB
NrE7ifAyptNqoP2JoOnua9bdNF0bU0wT+XPzzo4GX+dLSoG0aNdB5PjCXp9ZAoX5
iYia0eQuHPxlHymK374M60hMRjzzR18uR7ZU5/tjmdDWW92a5wjZ/33fIHKoSU9Q
CiTPUZVOpdi65GPe34ITnEdrsVEUZq6Lp1zPzwb/QH4DMSyAsT+0nGyX9mVEa+VJ
vRLJ/YDU8UgTppoaL9mFPYzf3Ni4p22sCTq4cGI2D7tF/sY08UYFsWoBOMn2jooY
MQQHl/X0sBUrDGNyQeHHST1SGXjmDUH4701qNUBA+MqA5BeZGAXUsa20kIAmqBBt
sHJAatohiDLs4b0f3kIW2QBhbgCIfmu8R1ZEdXDqQoY1K6RzOqSyRLb+ru9VbaWf
91DRRsXy42LShSsIm7xcMtLvYc8kXHlBQgPSKk0XVgiZTaEfwWnuokhtO59mbsc9
UnXeLXbLblkfEZuiD5dCPmNLgpqNxFDfgWaKlwar8p8Tfr8t4qujGnnjr6PBqi8B
t+RSzlcteEeJ5M8p4AvJK7YMopmE5Kr2oydBLdR0nuBoSdT6UqTNDn46iuIEEP3r
KtGDZcv8ebQhby7tAxxZ0SONcwfxHg2SqR2O8RB+yTlIykeN8Kcvhtf3wkqFaPZT
Pe3fmNBfPapjxdh6/arQ56XryL/gSHGh8H3HsW3p/+Ky2kmNwnUPr0d7NXGJuNce
wPIwkjQm4G/rwaDil6C8kEn9TVbrEIYdE7of/XdOPof0u2w/bJr7j3lvvM7eG82h
fN5hwu5BIav/jP0D9r1TQwsG2x9kzxRZzIE9dR2WXcpqjMUSzzmCWmjqRsNuzT6/
0Pzf3WW6L7WXG2fDpU8GvJDiWw/YCqhF6H+wX+noJE1PIYhoT2+ETCv0TXrUuVfa
osSfAXvwKggxQMejc87ithP23Wcdq6+GOgrEixB8326R6/NzWzwfDwJVGffuBQle
asD7rFaC3zSYUYK+LTq830xwolMQeZYcdYdC32RTNrH27d8013qAjCh+6wXnzHoM
PFspBmis76HqL+jn53hlQl8YcAx3uss4ykyYCqkqfvDYW9uNY5kP6/QvG5C50V4M
fPCVcYjZ/pHSXePsr4hFDMpZsaoMQWbMAmjbd0elfSW2rfCLYw61EWvuD94gPs0K
ILy58OwrhmJgyK6YKY7XOeruG0GLilPggJcmgKrRxQoNFMDUOtw3xVWKP/EqQXGa
RG/IZslKhCpkJrK/++ypl3infCk5vbLF1D8dNO53ZzZs9GpszNY6vQJmid3Se94b
761KYcAHv54mXvA+nLhAbZknUC64KUXbOV51bn+IjxNw2gPckz4y1j5A3tv3+G9n
CLjUXKPyrE00pdC2I/IF0fyAuiqPoCMRg4qbb2Hr1pLJKl2xm5ZX0qdJP+70Cw3v
GP8gkXv9b7Pmcei/TKfr2a8Ywg/u7BBzPE288wwuxxAV60XoCShRwaxS0TaI8MQj
Vr0LiRHv0Afpws7PZ5BkuAMDuM87cDqDE2TFgj10yMTzY9leO4RwMH5Kl4bqz48I
AHN0H+H8wlevFbXVePfGhPMZkIcWK3BVJ66QscGarkxDSa2i2A+1cIrVOzVKA85r
tXj/M7wVUzLM1wxvkdhC/ew8rReMUD8LA8t6/+7+W6zE7e/qDdIWvpg4PhGpmeIR
qPLBfIzyJE+/rPrV5PlXjKFVSyX10AfBrRIqfFikUG1DaYtUibZtGiQ0SAN4Zdvj
nTfuQKqdTfKSNxQcI5wVSIWj9BCi1zkwC7ope8fTI6OkotyTiS3tWQFkT6k4xCJC
PBQ83MUvXlatSq+YkXMHLpajGSv+RPJMMu/qSSIEhk0UL5bwdkoAGu0tm5zbe4FN
WH3W/NdRFfJ5mPhNCP9QhtTTI0QiwdXQBx350uKDRNEW/GaNoywA7hzFEiSzlXMO
UKPATdJyk3PFXMeU274+5BiqM+KJOoWYsubrtW4rdwQTSOld6HwK4AAi2YL2TXIh
gBZkaLoEJfiKE+kezTfS5jFMPqlTKZZzT5q+9MV/3/WenoZ2R2g+de++5YHg4gPp
x3jjJsFn3eDL0gOav4DjF7pzqxJnA0ftsno8mTshJouA8Fak9ikc9dNAUCTHwv78
2Ksyb77t0e3Q4VwZIz/21LrqBZGJAsOb/iYKrgk+P4Am/wp5RupYiRjMNGOrtwuY
NrsyuyESzKmx4j8+E0GtKuQ9QUjvaMb8mItp83q8xrWgNMTzveyeogYFc2ktinnU
7m//iBlwEpua+VcwXHa7/gmp1CYNeXloV6qrBUEfyIgWG7Pp8Lu9E1LebRNKgGOR
T7Y2dN2u2FdMJNCqZsnI0+xO+b61X0WBY9dXeeBTsyo/w58xfoLdRTIf0CZE+wit
jaH6uhbHI72Kv4Pb/eHhUrQh6EmFQbFphHYDWDQMwex7HxXl7i+HuMQI8Fv0VVbE
/rtm+G4rODSRN/HLd1c8RVytBi6SFgw6WWDFaEeG5IdRbWYgC1Vt7oLiMyO81aWV
E/M/ZfaiUdNNmZf2Q67S5oQBQGGwCaUKWDu3FsnVykd0A+CP5o4B50cAI8hwl8SO
vbOda2q2L3+7+vjUKXeEYur12VLvG3jGNarIxOAtxmRXGW4EquSmTWQhB0vQs55A
+c/XVLVbkX4Gbe9KMmXr+5M3KV+OHxzD46l+VIZboYxCCtU6uk+kQNdqmsv8FzG5
OnRGoczMEEslf7jWD1CvsrLZN9rLLyACtAr8cL5UnIakXQr09HghDr/4g3ENM9Fs
pFG2bLL+MhO0o0HX9xTd7AUMSVejAFyVjmva1xLuEEHveYoVuy/GxS6bFVyIeRIS
jH6wZpQn6qbGjdTRLd5Qnp1qq55P/5rAVpqjYhXEircD0gB01ph9/CzR896KG2Gt
LRS+dfhtNImEpVFkxThj+Q+h8STXwzTnD7INWe6LohS98Tad1r0mODNX4Vu434du
V+QoYLaqu4Epz9Npfm49mCLJaBz9f56JEZvMWF297BFmqojtRdrf7FEJW1XnRe6Q
quHfTHxvmNPjPqxOZ4s89HSDkdQXrBiZOvgt31knHsaj9oCM4vlLr9zJ83X6QjBG
PUcQfES4PLW8rABnMLftc8S4iOIZI2MtBxUz8WLycVKY+FRC5tWgt+y8zSb6IlE8
QC8XAXoTZkncDSXpAZkvKUiZ3uaNO1bhGQ6JiL8bS3BYR4IgiKTR/PGSuCiSAy98
Hg+j69iyN5wFjxxg1DL5Z+iK2rRSumoCUCwSistTDANtXuQqy1DA2Wlb4YwGDnYd
Ho7bXXmaUxXYT/4+ebwooG6gqwK/I+kzODLbNU5LVfVgGDLjkBeZNha6vscMD8LV
29HHMwR76qNC8ppB8rW99SWVrf1dxHMerGLeG3G8Z3WEqJwUkqH/qCeJmRQQZI4i
saBIlMxlLeymr29eVA7irFfcve2zZ1TMdkYw0Ff7jwdMjplsATr2J21rVYz1r5uK
v/+tb1N4lmQUev1pLiwjK/uwteJ7OL/A6QagzvxMd3N8v2D0C6hGf84TCXfQnqg6
0kw/guYIdNlsikdYW9IR9tvJxV5k84APVVHXZgC8T0oarGpQpv0hV2USErOhZDeg
uds/rIKt36LBbuUTL/dgq3RqNJzi84SgGHWbFgN4FXS6jmoHy3EQTgZUrRGP8V9k
BUSu+mFsCUzaUkBBjh4yBqvk5GoMHvwinu+JEaNAFq09M195GFQ5MXOLvz5SVtxy
RYuaZ4G6ovUp03oaZg9myXyJbPV5Wjds2gVIQUjOEUBEtOaiFy4JRO6ZUYghpjxS
B2Uw2Wz/iij8L5dCm6JDh9CzikZSixPfuRmN8JJalrMtWRZztxK46gkPXOkW5W3F
nnA/tkCk1x75iNlnLJlKgGr7qHHHoheXt5WgxmjWdj942v+STbWNui5KFZXP4k/Q
VP1TTThUo5Sr8UDVgou3cwDFe4F2ncpmiUPTBPKnBROkmqOsmzA9kt1XgySkyPFU
Y8ET5TDbJcRQFcwXxIBFtRtkG7ej6p3GgfxXWxXa6qYu/Why7SExaxhEuVxA7GFK
cvdgK+Ky8JaQPQTpCW4VWEyz//uj7jfeSFTSDiM55ZW0a5G8IGtiE5TbWPFjR4UQ
kqO6x5tvuS3Z53PHJfYw68comAiTEhfNRxupvgI8uPv+ECTPWYambVK23VE/96Ea
5ANGp2C3nYPQAwRoXBeboiMpzov7+YonWu/JD1EgBd5zCMbGfaF6fXUU1tcCn2RQ
H4FurbiyxFttDaEVqUZgHsnvcsPtxuJbtO0a6cKnteogwnGRAtPp5PHLLnD0Gt17
TURF6DZzmtX5k7IjaQjs3OVQmo5cyRnnCxOhsqSt66iRCMselZoBsKJV83aAEP0R
bjw7JB9yfV4Ef4zQEhPKhK8hI/d+LEjrtPayOrvxNzBdMLDviQgOmKF4rzWN22mX
GoVgvDLcyzqnElk7qSoTvjrEpk0KDHey8RNMs5cQu7gimeU6M1XaBXTpVnh6GJ5/
FadIBo7a/26ZArmV6RFBLPv/ZvmvaI0osgpV1yibAmnbS7YWwdbmdpwA6qb7CeKE
wEEY/N8u72Ml/0aS4tw7EuGb7DWR0YHU5zRPPRqlwpEAdPhROUFItgo0nKbOsSGW
zLCtj+TUX62aMQmVrXXmq7J7+x2k9QA36eeccsAmNZua3itkIDacnSalBw1KLdCH
pCNwAdJvrVaj8rM8kjhd4jNUKKEoaVEDzAVPxKj3MzSfm5mzif8VcvUN54fqyPU3
SHOb+phGonXFi4EVS6gBdmpieGnoUCIC9Yo4B3JKBFfEY/sEBinT1Ev42A5erJGL
WO5f2iPOnCQTKEvAI7qGzFHGEvHqaLYaUmoyJyAHjloEVqGDKcecQmEn+/d9AVbG
oae2845QRcQVHg4z6JiKvWeOWc/gszKDTNQZfBWvvNZCjR0XKarAZzf4yXcWNIAf
TADK7q/VvNbnwXfQEoF+fgXxD/d4Qv0vR1Ba2+Ipm80PCg6ndp5fkJP+BNUl4VG0
0a1Vrh/FT8tCgGxYyChi71uhrjn6eSzp8B3FTHARquKF0UR4mFPJAmaverfEA0Cu
icOcR6jcmB/58NvvcQaIlukya79lXyvOmvUNnICgS3YXSJMlBh2Nfg73cbi4iF6F
GoPd+V+tF9BwVRWb2Wz2/HkIJk/tzbDsreSekXJtPICpbjdY5l+jKe6aH0OTQJ9I
RDGkOTiKquH7/lYpu1A9y0OrTZElTQmaW1pOzsi0dH/GxOK6J1VcjOUzB36zbf3h
iBXc0AHDxqSI3y82hyiG9htOgXmHqawtmorj3gX+huF+1/sWUsp73xmJ4wCXkKWg
XB9A9vn55dc5UkqcSTW0V1dGwBYJCsXV8WmvD1tOQtIPgrKgLXDJxwIfHOzxW0je
mdUdK7hitw+gVkQEH8ctYf6VD67T1+3u4aZdrzxYwwj6DRUNXVhl8w2oCRCoTwqs
hLCoPzM3eb2AT/YiAcYztQQCJiwXNsf41M9py1ZloK+h2vz4hDYNPszgg/o448W3
e+Zk5o8PhnPGpWPXUqmqvJ/PxrJMy7TxbXR/81YXEnp+CY7X9HyQN1i0K6hO/RJ/
u/judYkTZ6tarr4CoaGHQ6NN4xN36eheXy61OKLDUoO2v4uC+2LvSwvYkac4ZFmV
2xxmwxnBpoT5jVTs4nGty7hdAenD0qqHDRZdyiXqFCMkKBegeGHUAWs3NOb9om8Z
K7L645o5vQmwJkEseHMBSaEEkl5pDkFs9B+ikTWbxa/W2S1wwofER/6A1qLr3V+2
u/16s08O9pRRHPZj92TE0DoVDyKf81/Hqz0fo2/1+WhgS51YnoeedHpQu/o8Dg1x
wC1p82Zi7cvdfRNPnwtml1aQeRTtB+HrwrnaN8aE7C5swMqwEYCs/1zkHrjMib1N
jsi8bO9QBu7l37NDPF8BrgphgW1rIuQ9MyguAsn3/DqDnZw+mu/GbE0AbwD2Kxl7
8Cl2grUDi+CwSjAbBlnz1RicqEZxeqPnEic3Yt+o8NFqyHdbYf+LsEUlZsUBynNk
EqO5+OpmKpIRsaPbNRzczbnFYV49cjfp8aKpF421hMrloj9IDOn98PM18zru2iAf
QsiZHAO687dBnzCwAoq53OK2q+fsVA7xka8Z5ToSKmuyy3920CWwvVNJdGIL9Y4c
OR0cjYSbcA7e2j0Uyd96iZqoSdsNnRr/VsVFjd356bleexcAwADYqDmgJP8mElOH
255fiB8uxYK5W5i+vQLSHJwfEyx1sMpwfbhaOu7cquynRw/iZhbI14l9oLVsycZz
+kWxGMq+RyN719vWc3S03J5JLo9/f0PG5LtPB7eVCTGQ84mDDnW4eekOGE2h+Oew
62aV4nmqUNMcR58ule9/X2WbviTf6NOu6O7KaFCX+B+X++5Lopz6MTE/n0rYkAfU
xlLtQzDWRHboxwcM+rh2TrvZAYVWnaQKJbM2uriOSSPDCSlXoCuOgAGgT3V2e7Q+
3WIDof9yn4CfkcjR3nYRNMnF05FGaxkr2Qz2WQYcxbqEAIanpP8pEdrQB9iHHhEI
7/HuAk/WR7DfQTlWlobLjyrOk9pSHddsBlpJ0HO2/aTuCDsucWJUMKVCWkpYvRn1
mxcSUW9YI/8VNsgg4cTIyy4YqNsu0DBOerR5zweilJ667UODR2o3LTufSzrrDHq+
WkglS4+oJidAfP5YGe/IsqyrxQU8Y+3VctyEOYKtaMxWCBJQIMwdW4cZQl1DS/0p
P44zMH1L0PrmpaS+dDGLpaiZjsyd56nmDzGa1/Ey/XDnKaK7odUDCjO+FDqc+Pnd
7IwfJeQibOpkYgjb99ZpatA5W8bXYNIo765yRUFayVj12owSulaW1dGWEzD65eQd
GGRih+2usUC38IZ2YloyYmJatKed5iG1lGEiG68+La3GOEgOnLaiNAQFwnSrxjmO
D9Kiafz26ndiZ6OrcX+wNCyMOXdu5A17enlgyxwFrsQZQUnEviATWR+HtJ+cqZ/p
oreY+gkEbP0NddN/oz+ZGYPZXq8prOvbrEPsnxA4ziEmMBAKS/rLOBU39xGnu110
60Gd4OgWfx2kh9sRjYn4lItPH+woI604dO5khA/Qlxuu3fy8I/xkeOxjl+Y7xyzQ
9QIvV3MJToKGTwrMEsz5lnFYisDtqm7Z/WE8VHwmuPuT8aDxK68OhPeHNqUohVKy
iUT/Ad3x9YQ4OCDe6WsXzT/5xJJzFUzLfKI7nGH/XdMPDHnCyShj3R4+6pU/BzOW
BgM5DMh97vZJUg9lyTOtsJ1Pcx1URcXpZI7KerAARWGcbzBU4vPqxQEvRbDiOUSv
IqGkWCuFaW81/bnrb1qoaiDT5a3N056kOQpulU7riJS1CxFwm8Wa6lRnjM9Bt5fQ
wDek74MT5b2zRFXiAoVCQdOD6RVEuv/3yjyL4gfU8ohU78MhRJrDn1CsWlxVjAza
SckBtz9SdCGEzSFAatbgTW3F2HwnEAEbgrYhyYcQWtxu5HPQ9Medvl6I41aJCTAa
T74tqdtVSx52GE6BWqPcXvEbMeP5y/zovCJm9mveTtXEjlLLkU5jDZVqRJQtVwaV
yBodraNh2fsHtRZ3byFswcfjV58+p0ZeJX2INVjsSnALun2jL8pt64cr4hZHJ+6I
Cy12i5AAmiPhPHFSXNeZAklzQIM9ZCyEIhCdm8BYoE1iUTie/fvEpb/qYgjLoaJt
kkJNlYlIkdYZxrE2Q3sqPfXS55jwwG8UJmNkIBKUbBicFJGkcNvJehHSmCNxRYDi
mS6QAnMuQlAvz9pb6LJ4WghbzI0l4YoXXRp1KIn6WtVvJG2216HeIiBVYaFyqq77
SS2Ee/Y5a2iH7mH8b31P/IL+V0sZ9U4BNZ0BcdAV/rrWeCdSX96/t3vfZUy1YRzg
8G4F8CCLPHeauniSp510gjIwsq6Y+pDp4Ccb03ZZZerJhfTHl27wvRhg7CgZmTIo
8nD0NX4I6uDDv31Or8jFqT8nx1T8pwFv7k4yGvQwvHkafX9GgmlnMNFBTTGPQHXx
aQxzAoljtVEs5hQjhl1yXxUxvPR+ZkdXSmjFjdr4fZlRThmJKQ1J/x5iwUUfue+n
Pp8QePKOU4sB02AuOOZmUbRYosQhEJc4AOM7QgX8a2ZL1TQyROBIVHlEbpdGLY7t
yijmhkFHu/ViOutqAyBjGQDqorLILuzJu0dr1Kp6RgpsTXMwvCpLi/xc6dMLvKzh
EVM+YSS304sdr4X1smYKkeji4HqILujjVC4SyaG/FWzXOyaLbqqGanLxT0zwmeuz
/pj2KsjQ9YwVa3dOSwfofGYaN9WtUUiYIqv1hcAhudA/Wi8sXNi0myBlskoIhu48
+3F0V3veMV23Qf8teO+xIjmDQi7OTyFfkrpwOXDBIihwBRGpCeGmUCazeJ2XvHjt
MC+flPd0gLKrOVQbLfCLygtxgAzyObpKi/pkd9kITlG/OBHBr8LjvR8vRujlbxi4
uUEEGRRxQyH88S26Ab86UXVigbFLXt+3cWY7AZfWPrPUsxKAhi+ndjAnBdweDvCo
mEbBXfflZkDUQ9fZWEWVctCGRKafVp4akECBmP08F0b+HV8MfUQJINWmg8PcmrnU
H4nauXRkX4pV+wpy9HPPL9v2f74SBhuOGUp5EKn9G8v7xxhcBC/MhAL2WpRTeeAa
QqVHwaq5hSOhszzXd1F1ltC4Oor/P3Hk8/K2kIQkDQuVQAu/ktSZFRs4q9FnrA+s
Nrkf4BAvX2BIppDJO0dmhZE40jnbcSpO9b29HEV7QRymx9SmNk/ZSrI6xrWXOkcB
JiaPi68u3oN72FDMo7iw7Y598VR2RwfjrGpmCHhDhhqF60NLr+F5fN1k1NdwNa9X
spwQm4XUONQvN0Wfiii7LzJ7CrWG17DdHGHGvMDCBbimm2yaHSZzsla1gzfPvQg/
HaeoD0uEr3eMQQLmsN3T+lvxHmQSkrn/oW5sPA3YqObaHiV2YmViLs5OoYHEdNJz
6PWba2V6Aotsm2jSSJ11tfm/HXlnxde/ADOqTD4ytuM1gAzrqLuRBubq2m5cvShL
b9m0iSdwBZwhleTt2AqCtQo47+sE5fLhiEla21ukA+QmQG5jbhXhgPQrW2IwSOgK
WflUc6HueeN3KGJHeEAR6ih7EKWY2wnfPEd1Z1DucrGPykMHkh81J5u2IP9qXBgE
RMBqjkLlN8JSFuAGGUwWdzPBRTbu44P8wAv2l2pI5p+CcWlG40pCB5syz+NvOmyO
0CeTiBof/eJlWAW4XHMCh7+MKIp6YgP95rfFV4GKVhYvmAMvI0MK3G9F0Mqh43+e
1b/ksl8oC+h40umeGE5H3aBftq63BJkvAxfQ2MXR49Ouv+UFJn+on4XmDMewoDl8
CBIRZ7T9AK1qxxG5aR8l/26UvFnadlchi9yoZmqEmLrTmm/GhAD7HWweuJZjkD11
kTYM5lUSr/PvitKGMfja27FkDSMjv9pwOVaPMTAhxSl3kwtj3KE3DjCflgSM69XG
uc/t2HUsbDQaAqx7rtuNpQDfrAOy4lRKJWjQ18Idc5F8GDUX6K5voGGB1o+OwdbT
Yp/fWpfxHjGkatgaOm9VZ0GnEAj33XOVx7kiLt649T5GjQk+flLIa2D05/qXRdtC
2OflQckes+A4EJUCyL96TWHWE7MuTV7NqBngV58rcQZf2CuFqaItqhH8Xwu8AYA+
aJShPbLp/9oGqLr+RXaPTiNyfTgsX2faPRi9hUGnp7ruebd//llZ9c/Lh6SSPNXn
lblMUbdz9hPw6AciFGz9ZOkyk2X89GJ3cFzyeWX0qYQCSecUk7hcfsMPoTbkDoUo
b7WyoeEodWgPbScbVVKO49QvpSpD67bwwvQEKWGYx9xjDzB8SX5sd8YdlFnRHDMe
QrtaBlOxurhYcL8kbOTZuOZQEQHg88iOX0W2taezrq8f/QSLJTfXRkQLZnJVIcDa
ZVM9wjnTzoVb+XNWU7Cj+2ZW8oYbMsYAe7GaM8rND/ZinQk5hLQ7iqXcxN+Jw30m
1Hy/yl/8A2tMa3y3YcfodBIuBZ6HE6dh5TSKF1whX+S4w5F93iJpjp6pf1TAYg4F
BMFEn2j7vrovlTiEIQnFbGCaaR+lBpxvm0Z5L2bfRI3NVmOoSEn2X7e7mPMxjLgE
jevyc+XrGjyf8KpwFf/CLX6Mu7hFmT/Ww4Fq8kEZpl5lTjmy5bVnIeaPNZAqhLBC
Bg+GojfD+Wa3TIEuiMBFUjGhaNJiZ4Z3/y0UP6kc9x9GqJbZVxr5maIzp+WM33+K
TB25BqT4MEVbmFDFRyOOn/yapTMXMVW6RNRorHkhX1/M4a53l2eunKLADvZ2ut+R
JAcRtKS5L0KKtTbuMmDtvxHoDVypgSgtdy84MPNcxrtWbiq7UlibfDGuHA2LvTYj
vtUrkuC95KZpub+P7zIZJjIV+P6zDEiVbOi+0zfJAdJk7KiAKgGH9uFtCIGcf6JV
boP/auLVNfh8RzVoxYy7/defRZeIIRj6iZWEJOXQyMJJ4QhXfZZaOmjPlRF9lR7G
RMheo0x85vWegMWu1jmstKN4lex7AAsSnowFTW+Rje2om1krHA0F9W+y5x3CEtyT
2D7JeKlLQBg4nnBEmRwuUFBJAtZgKVIj5Af1BcStN/PC0UNqMm/JcoisQxOOweIi
A4mzqMx44ro+4xDis2ZGCDSIHIIzZziTJ7AGsksNgzf8BOHLAAxSdLA3lWqX3BPt
TAiGvHs3JUsSu0cQ2Tm5PVs4CQ7O+/4UHywL3WCD67wg6rtGbz3YoGShzvGasHQ0
D5ui92nk3l1vRVg6T/6mVJETaxHRTeBpYdliEZpg2bCS3CHFt5TzQpmXnBoBZkc9
Im8YUZjR8ijyeE2wOtWWBlxdKj+RuMxa8Uo020PNYHzpFmlXTtVR6cdPl3yjkHFm
nqTWmv84OBbcM24a7ccEwgmfgF0Lv4wN0NtgMola7AKOq7bo/UG7B/I7m7Pca7v6
fkmmotMavhS+HP7DUqA2SO0IdiR3xDpJyzLABvhA1UiFlcwh43eCJzR7bdFEqbj3
LfzZI77LbuJUZTt5IPCOxGqiBWOv5PbWyRAAuYHgIP921QZeLSjj15L3gQb61puW
Omp+SzotSCLKEDlss9BajGbfafFkW96G5IoBuwgi3YUi1K5ZHOQLS6iG84qr5s7F
YP5dt3rH/0yy/tyjRY8kk3nf6pCRk0+dySpEfgkD0WF6wzDi/4J9sW5MJjZhLhW+
v60Rzh9341FQTRcygq5GcVV7gxrluHoHJtXqHgzQHSyy8j1Z3hlLWPgV7JJe1uBy
ghmLPtujOYWRBw2vw7O1tAxPF138llY9CsShpeeADExFwlDFMCWJ5vcmsBA0H/Eg
1dF3Z5Ba7agdseOU9K5Eep43CuUeCFL4liMlKTaoy+Jud2I6/Wa9FjKs6SqC6+/v
Ef3+yxW3H6FlePs8DzNWk8oTMBV7ZdA2dE+LLqH6uxM9Vh3j3x/DqXYWpqVRYpi0
sb/AkYj3t586kVEtSx23Ln0ZYRjsGAdn6AV4yuFbmjrZHEfaWC+23ZmtGXtg5MAX
8ioXvhWBZJTF6b3YRRpH3651L6ZColVf9n2rgot9eqGzcpvL7tm4V9cvOnlB+KgK
JaqKePLQL66WHJNEPQHZwGQsLtVzRxuGT17NLOnQErsswaZfhoGFAnQIEKhoY2gm
WR9f94XgPSIOdzdoF4QIoX1WgP5jsVBNQ6VYN4uvGd8VEmOFiJU1QSEMs2MdosKJ
6m9hNp75T0+EENb2fYaG9So1oHdyAwc6pFefVvNxK9H6oNJfTcHjFag4E2yQVqp3
YIEiOhMShUl2eM5V/+TiRU6RynPBdB1SqHkvH3AupyIanLhkhdmTQP96SlRWpsgu
1mdaOX9BV3DuinucB7IC5Yk5QXTT3L4l/yh8bN6+aftBOESA03Cl/KxabB+UY/Kf
1e5CxdanCFdLEtnAC8TJ7hKWOoIe2eThIpvXELMTsQ82jOwPZrY4J/mT/CeJ5bZM
cAaJcF0YzcxnARfjHBX4o5yl6ZyrvKfLvEP3Vg77WaIXAyQT34hAkNMohGDqUqwO
LmwZtPSs7v3GY6h38GeeEdyTZyq+UO6XtIoISm55C/w6G+yd84k0kFZEe8fHF9p/
ETli5gfrRIS+BMXp4EYfHXbk9AYE7Qr62A3626JJjnndTe8CM0FtpZChrdjOWo14
jhi0wIZAKN2abwUmTy8YnxSHHv3LGAUJB/TFqGk76ont1k7VExonjKw+OAzLsQO6
X9HblpB6czXCwHnIc0Aj6Al9lx9f/f+eP+J+aHQKeQEg4tjfYkYNcOD88XuEXiNk
wGMQHKTipft8UgU8QAZAMNID7pv/MwFkm3h7oIyka0xZQQ+/Gktuh8Z65JBgt0EZ
RId34zB6NDWFU4M40PevnQikjc/eG/LGYZrHb2Q8Y2KggYZijxl+Gp/um9eJ5+fH
mmuItnw9G1H8Sh+hse9Ogfr1JsQqj1AOqZJq4m19v5B0LOb+2hhNM0AS3kkGeUiA
5qmaiQCBtwjF4ujySo6TfBEJUVnU/+Bw5MDU0JelVRZXsfbWqtbmtOci2+pz6Yej
2STJlS++K576JiE1SwYM482oldfu2JK4OkclhD918aXKWzVLIdASBpzhh6ES0Fbu
TdLBzfFzMCwzaFf0jUQQ+jMlITkZYI2mtmPXszZxyDu5R4MSzZ2Kyy8nBTdyOdlL
gsEp/FyKPW1lG3gDextzbIdY6mpoGxIVxYoL2IfF1kaGfzXwUbHwCMD3lI4WVj82
vcopwdmEOA1iKT3/7n9vadgrae7zEDntWBLySqkJrJMbt2RaoASnnFL+NSNU1vY8
51TWY4g7y5jjgkrVNiAVaEo/V5bpqIibUrTtsKqMNRV3KU8S14aXK24hkvDEGFBE
nPVsF0M/8veGLozmj+J4pARdNm/SVwhs0Ve5yYznxmrV83JAGsIeNzPV8ftk0NyL
sKppqfmHR7uRnNIChkKt03s6cirbZvxoHPXASSEHt+CfzWk7/XXTkh/U64LE7rcZ
w5q6gaUhJvYfX5TsiP1FbnVwXlIV6lu/fl5+Z+UMHu0bg/E1PoW57gKmnaRrFr+b
u42AdzmEKhObcyKhLBrcE47rT9i2IAQCDwV6GQKF+13OpqIc2ebyuZgIdRNKgJc2
/m568dYyZCT5niNxXHG811vvC9x/yv5LS8M2/9G+cFYjRSYue95MVub4Xa9zi3nn
w2YfIiKYJmlS3fgyAWZj5+a0M+2/6+x875SK66y1OaY53hdFPq4bEcNpQQKMo7nn
uwSTKAVhQ4F9er4YcEH2i3KSKpirTduEdUH018La1uJ66wxperCZCl5gzk347wYs
QJBXeAtiWs+gsSVU+EpbXhYd0pDkcvcRm+s3diFNjJHUWHw99iw92lz24kcnYc/2
OoHLvdtSFMdfETKIyQ4EAi2YwUJCm8ppZ8WRvIl0jzd7QIU5bw0KLraO0FeVYs3Y
rrQGbwIkjcDB20+gDjEhkyDPcuLEe2+qg+U6BfPJmIcUFWS9mAMZjPiPylD68T7R
9V5tZir+1Jh5ybHRDNtcZvA97wpYoUhWXvuqPlxyP0YTk+mkUwRG6vVYLpq4UuEl
BkFrVwoZWnK9NT6O6HwExLg0ecwgnckfR9fh544mntqwqWq7LfgUMxvaekGhK1UP
LOOkkDUauQOG/MkWbrSHxNkkCYYq9OgcpjYjosSdqYD1R6ckuXGbax6eEMrT95MR
7dXt+ZGBNwxSNQuR4k23MLxB4ZyMdEfh59rDZA9tVr1r9VMwzmGXJ4lcZEJj7Q5K
+k+Oi7HCsAGBDGm0kKkieCOh8qC5gmIy8JsMBFhXfS7os5KPWsqRykUTLiOv0WD6
cXAV1iITQqVBcN04PyGATUOCmWr3gP+NZHxfWt9/a89vEHbWqvSkygXLZ6u7ukbQ
GaKdFOzmROIERYwHJWCvpKzndic+dUzMFWBJsdDXg7Jgn37xacMyvpyD72GyCTux
LlFvZgQVL0cq1QuoTTAlr4Uv+HrbjuyDRwkb/JwzQ1/VpuzRoIlFRRYUZdhD6f1J
OSCd4Wd6cKZZkyIFWpvCoHF5fXy4YMVu7cLJ8RRadEmQ5/OMRIMlFPRCY++YamA9
kFtEvx4tQJZu3Hm53B7j2U0LkEG/VRoSTPDi4fgayIfIIu77vjThWIB1uguQ3yNn
IrmCHdcPbVvC5PoKWPVym/qJ+VduwjAuZys2DA3Scecem9xmUytGqROwmOcPbH1g
R6r0yAD0a7SCUijtbhrL7L4bW4nto/iRhBUhqrqakCjFs/mhYsdVhil4ucwo6QB7
DloQ2U/Z1ekYM1MtNqyvKIzPEPRnfurTSlcwJsN3iDWoX/Jl+6TMFx4nOvea3VOW
cLICxB+VvtBH10BpgGFZdoaRTTx/zosWyLlulnkXYpfJqGA01j4olSXLxBFE8G4H
8w2aRUY/yXghFVtPSgAWkbrRBOhm363e/J5xmdaccCo4a4XKVaUVX6aqCeBb8LQI
RkfUI56c7fwjZQRYoF3fmumHNuMaqRJzqa4cxLrILvOoOBFbQaGWwltAsRHZIEIX
ulRZ6PfqiGfWU4rT1gNG+J1ypNIUDRi7cVHyhCD29FLkZN4987TIFLuFzADBKhLy
AowP9Y8h0BJsF9SA9aYUwsLuA72sX1BYnRrKwJYuiQNVho1vHleMrmgBHPxyLbUm
150JBKvDkmrcV0JlMt4Glf9OqG9Q5p4K5ztXw++Smh8wm02fqtf0LRX9yTvV0zqu
DyjOjNXXTk0DrnTfJjMSyrTCw5jcNtEAf9DKhV5yAD2OhlV4sE5bbo65xdrL73bs
23k5hwitRTuzb9MZMgLOlfToNHjwtLybnFE7CoRmaZUxfWDZkYTzFxwS2WalfQa3
NODJ9Muw3ZmAX4J/QkSF49dQHa36THiGuHIYExIM2gJyhs1NBCfzyTBO2DTPKNcj
I9d+tuCy88YhcDkn0DyoiFbZSidVdNDbM/Gdxg+lC5Zcez6NiBTDRTVqycZuXLoq
Q4I4cndgz/hQjr9CAhDv3pMB4MGkyQGLMWjohEz1sUEXmlhzjfRlRjeGjWC53ty9
cBVRp7LwO6LN8uEtTKJg0O++PsgPXBKETP+I/ZVC5QIOAsVuX2MjL/LULbhrh05g
iDV+6Ubygeajm2U8OYXtYGuPpxzP+QTfQl3EDtDAoF88hFjCvHtZwl8IzWaXBB5V
Nnu2OzYIZZs3rksuQvZClSG5eG3CjcoPLuluNT33Vz1Jqd/u9RLsaTj8o1VwNmsK
4cgNfnIijmeFPdGVf0QmbGDHSjl1ij9/JV4+vgP8GhqXZErDNOuXrUiDSMes6rN6
a+SKHJ1P9xX8bbFyUv9NP2m8qqpxOQzxU/iy/uMzl0r4cZn0vaj2MM0g7sEBEnPI
7WXQZlZXShawZ/mTwsiJShHDmgo6vllaWWB6/VLhCvCob8CBWOHe/2idZBoYUQrr
2yRVB1jww36CQQep+YaZxYgMbFYVZoca00Nq0JWd/5WVxyQsAOoCe4Q1IAzHjrRm
YMGXeglhw8AhSrDd4r42oA+1o2SxFa41NE6P6gfJn3Iqu15LgCIQbELgb/rNtgO9
2Yl32UcZlXpSEkp6Z8HoaO9htkUYFFTlj3VzU3hYl9hmrGIxQXRLtc1AJy8RK8ju
+JdkEav+ROQIXGtDpA2wlpU4cz/ozEox67TQzLXQZoBvoFpUJpHoWZKalzYTZifj
V3vchBToqwZqfsLx9XGipC+mvk6FmG/AtYwLRj2salNdtJ+tOC6ldw2r8hX2jI0V
M+3zGbFJBMxjJd65YHQYamqtdFRYn7GchvrdlZFcCUQNeYvjLp2fTiq07NIlVUnV
j6WKQfuRKYiuFHzqD/AAuAco+4CCsQlTywEnIeCvwL2wA8UpSaCfiLiyQNkUIKSI
5CXndrBsRt5lOmykhiT9z35O95Drv7QAf00vfl5gZPN/y3O6RxWmJBXQrREORfGx
oW+X8D/yUuAHACzCHf6xE0wOITl34NAVyP7pEeuDZvwZMs/8COIFkPOrrcuIt20p
2Qu0QAWapjnOQT34K1Qj0P76owmeh/jljkipzb52ZyDqpCo+9AOtIu2/6spdm+oV
5JxqdONwV472vXTHvlCqtbaDQU/KYi+kKkhRwRjQMXLvz/gaErLZyDrJHOZa25pL
GQ6WBbqR/TV3Ztm1KDKrrRQfdR9eed6mlzIIjseWMtH4ahlx7BQt+ixziuLiheAg
Plc+wphUL2P713MEINeUtLFGRwZYHQVl3wlhMqs+R7g38+KxriUp8W4Jt2MLKKrM
shvMpl0ZKVu3nNA7rVoecYVbV6eF+SFRd+A/JzoXZji0csMMtsV646caDNgXwcuL
pk4ylKeVVIBKlRt1ocAj9JTfgFpaTipB8p+OdcT0pCPMNjlBWSfFI93W2L1OBl9t
VCFXXwG7BgcIcXb0AcTy9DNKQB4l9f+l9Dd9XWRe6tZogbwKXGTUTTrEvTMvQEJO
6x1Swq0I+/8qNieYsLt2juFXMqaxEw40O3vRSyeTFQQuPQRnOQMfuG/O1xwQqC3j
NfgIm3okSI5nUoiDpn63/pFB3Qz9VvQBDpEB17wUlQooCnLj7jpPqZ9+qIAva1Z2
UAU6us3X7o7LPA3+8OJwAQqWJDfHjByThlQmUrthev30+oSGZaWBOLR1ZSlpIbOX
DoSKw1WGdkUyP2qpgQPsSGn0v52FFA/T0fCtVzPAxMq0MP3VO7JIdIhaKW48gCGY
iRJuAaWWrt611/O/wYmSaz1Fs9T/4QogeEFSNhZG+mppobOepyC7EvB8wTuyLEtl
WlH8gPyLl9nhmcOhxyVOWAMiUMY4f7wIpwH6gQDT9voP3f56ietHmqgdCoAfXgNf
zU4feE/zvu750x3K6Xt0txeOluZHxS4IdzCD1+gG9VnaMliaCxT6rnw/bcj0mHCF
85PteHgP3w/BrgdktBhroZ051O0ytVmDJuSVcTUi3ef+dLrjPt5NYoy9s7o5ktMm
kYXJQ/kO7jUjK5tYk6IeI8HOuye6BnnAcPsCLRusQMiqH4DwMU4yUF43xSz6Gqzt
eTfxyUbUnboIJ5ZYeQBKQx8H2kMY7VKL4d0w4HhBisyr/J72e8HcY+Sic5PlaAgV
66VMMDCdiMGCD5NAT1NR1K/fZvp+3xXYarXx3W3wYEeqzEkPxafGIiaYUZKVMZw6
wZQRuIj7ph/ReC8gm+meJLxxkixmfB+mPA5jxOMGJxaFmbr7Xr/j9tHatQThBNMJ
nFQr9mx2ADEtFQoH5nujqd19B0RPQu2b3SM+YIl0FqFeC+kLYeH2Q9XQKIHeTvEg
953PuYY8AH6BH+liICj+Q75/omuPg6bHRqtYAUheKDW3O34AYu+0qCBiNJb24z3p
JjpVpHGZ0s85Cnu3bu7/1JnnLOdCy0GXFEhr499b9YN+xoZrLY0PlF5CB32NT1/1
+x3EYJ8o4UOek28dXV1XFw7KQ06M8dPJIyNYtvp/sYAVuDqcD7jdNdxzTlgAWEDI
17OQybiM2moMPvJVB9P4wyvudn6e+gAhmi63MP3nuXi44YKIjIWeGlyt6q0RHniz
J4B4P0onHn1CPWB2aE9CvqSJp4VdUxRbG00pKweM8Zb7h9Bj7hCR8uWyvauAkCd/
VxZI666YKNSOUBeKZAlQYYfudjOyz9n5jaGrzVDAEQ4sustomTZmo/OwOA2hxnXK
RTJiTfWpI/kfBZtoSCE0wPioJKOoIfY8K1JO3UWE05XPhrIFYUmCCYP2IEgHtUoc
whOkurRXhfkfw9iHW/PSTwcjmskyvhyraUx9Noezf8YofGU14qE3jaKV6ilRibdj
gchj8Hr+JtW8TRAQeRA9194Kyw4aVufGLz9bPnbHm9sOunowAK/mAFPu23frzuGG
DBd1y3dF9i08xyQd/6y8ydJVSuwsGv7459bS3HtkkzU2rQhA12sHkZAXQIm9qJ+i
yLuMp/rEO0HYL0B08l09SN6wqpycnsuzPzNSCIsAIPH3AIAuQPgBZzZoVhKTM57q
yPW5YkpRPMdBbEJoTn2vSmYkjRvGZSeJ4XboRY0ih9AkK105hXYGnmh0tL36DqQy
hOsKGoqod0LJ6sD0d0Y93qmjjcFn264829XSpDzwuzoo2kCVwUMrJ1hMuoajMGHZ
/HBrOf2JYhHkh/r1TkpUov/oxpBoOPAYGesBI7j5aGujSmd5xxI9N88CwrwIFAg7
YZTqJUsJ5X6VQRUeAkrYry4w6BUdQ4HXzDK7HjWHQy6VZBU/waBSlpG0C1e9cHCd
3xkP1xQGy8MQhjhxNxaKrDDcfnIA6p1bUxSE5FyogSZYsby9AONRzEXw5QjayWt3
XvAalSPytecqqseQiLlSXpzDcfYROpZ1SgwPFVsHHI7sg7Bzdi4FjhixsQKdSmwf
Mj6JN8DOMZE7Jk268Nv/4fW2B9G3oL5PdyhIQziQcxqhhEvoM7DvoWdQNwD94xlN
5fnoSXek9XrkXMdSDxgJhf5zJBB5fmEycUAfdOR0IpeYooggSah7Hhmv0SbsTj/a
qkxiIjI6FxSG23WdILDl1meM4nrI+VZD0N0I0VuKZQw1ezCkiQB1gucmAuo8YTSS
MbxsonezN5A2K7F8xtodAL6450N3QFe0O6IawfuejWCgCDvPnwVX8pnDM5lcgUYG
I3+ALlslKcnRu/ZZ6liypXQl85BHJKoQzjK/EYRN+ckgMfNHgVElZAn2BOowKScy
6DjuZXqaLyQZ82Jj/FfOVEgkyRgFRUJHAyQnKQKUjYAgdiBLd9JVpK+O4hJ5QAps
75zJOdZgLo+k0MWWBWOvPMQveHOTvE+VJViO/90vEcWXdY8zJc6QfoGwRHnMARYS
M/bx4AoDBcKSX85LVMl0V6qrhpYJAsPPrjANCevD1sGfItDQgRRdZwqHA3V7JjtO
9n5trM1s4kS9Xi5kzACrnQP5/I30F8kqE6/pA1f0v8uTTY4SRSfQ0nRKSNpCEP/i
NyjNfV3M4FMlZwP/DBtN5nkXJdPza4jnPIBK07kNVtw/hz6mSLSibK+CTu2OesW2
niM3GT5OaEmk5MBcZan2UaadAn4YkM4vdXJ11DMq/FvItJf3E18hParqt038gufL
QXJ/gv++j2gPe9IQNfyIVhh8O1rNLFW/5BeMU++L4CIV3RPCeR1Bk2HG6nPq7PJu
HVx3vfQu0K6JYlPK06IDavNTD6bGeXH6Nnbo3sgHY+IQFt/HK+6vxVpw5gJV0Bwj
ywCzw3Rp4Fz9kgt+eORLRIX8CbHwbnLISZkRlqz3Ji8KHv+QmYh2dHrIONUOh9FV
d/A6sCg3HAWTyyaCzhsSP2bz4yAUaIec69SzHCTkaVFH+qy3HR/4IIY07xDvm5kJ
8vzk+oDSqyKShbRrQ6scgW22GxOkrbhpB407W5fjmdSJAEwkpUIIOTyox8dA4b2B
YT3vvaqgtZjP+OqVjRKDfqMwMiE0ahWxWxU6JOJLL1cpmMqDnTdd0UjvQZkZ8vMZ
UWqLtgSK1yEA7Rm1XJ1QAX/EC4L6JeDv/9/VycB+yWOpyvXJLh4LQ8phpqFh2xS+
r/aG/TO37cAesDFDyvGdQqhcME5QgJGyvcWsQYBj3fEBui5UIQOByIQi7iv1UznL
r0/An8Qn0FKDCfrwpMvQsbgyAojCU6KkTvpcBJ/U38qUphjNHEzzftDhg4R1LWs0
DQrf0kDEkqr+iQuZIxQe/ouunlv8pD8j/XbhcglCgAuYVg551heSyzx0xhyX5CmZ
dqk2NCiY2TsNJWSbpFg08e4NDqytMWbTLpvaoGln9OgGYaNtDv/Z0XoCIMnktB0o
/1ji73XHqU8sqqqAhF1Won0PT1dpnGM4uL/pme27/j/P7Zc2W8m4OD/0x2MoCpfg
x7qqnCCFWqLWYawVMuNW661yecWwILc7Z3cXiH1O3m59wk/YVisxpuTUpZuJZWu7
aeVF4l1qVnPqmsmVGiTJ43886Ou7J9dUWJohDrfYr47SonVl4eXjGV80kcUttMwH
uaZeBEa0e9MWTi85S9a5lloWP8RA46UAVtsvP5Pu1g6Fg8v0Qs6nmy9KbTMrQ/FF
IzLoH2K8EWImTuvZVBtFex5on7yUITDY+/QqlZoToCbPPF6yt6l2ViWhlHs489T2
3rC4japkjB8Y+MmWNbneoVB30yAwHu3tNxc8aaxDObl7hxolr1ernzh8/xdiNvL9
YweQ1K5wivp4b0/20PTk3cNqLIN1sND1zsDnQBcFraIocA+GV4PNFbz/TMNxlMH+
LZEVgA/Fnaqv7/PMYQS8F4lS611dtBY+aPE3NH2KM9OfeBJnEDS8ZwrGif0l5F3r
BeJdYyM/EvC9MXNIo3vGdfeGPU90ECB8INkNK+Asw3SDvHmV7s5rA6+MF1/Z/Dbg
2o9KFfHeBCU27rCCpqagFg2Z3y81es7x0K+hxAdf1vS7MJLjMh6TvhONE6FaUQyK
06JlJorZ8VShzcpC+1TU+zocNldCLMziiE5BMY7iSaAgTS87pwlJCpL2Q9TK0jSp
yq+f/asqCv7/ITy7brocMKf3ztj70ZssqnkoiKKkEmOfdiWA8GhFQ1jtX6MZBNKE
3eIoBT4LppHsvk2Lp0RxfkP9gRsQy76Og0fegtnvOWx3IMGCAX9YuIVWV7UFxvxx
+Y5IEYRfwZoQ6oGtjoop1Y6IpTKnWnpFYeu9g5DxlUKdwDqZV5+axSffM9HSRZ9C
ptLFUebMdlx8UYylA2LVfT4En8H98OXKmjahbsYh0IhvoHzKXHm0/7/73ztaoY+z
EWJLEy7XJf9dGFWebPWSP+m5ePAZ4d3/ZldXN2rNE+lMSSCgO1nN8mt1/0NK8PCl
TTSFNvzLFo6iEKi7TjqG0SddNX4JFNUT7Pn7xvonL2D9Hb0EDzQw8P/Xg3QzsOov
k9kBiQauGL3aE0cD9oq34JI54Cjm37qOtqoxxz2oZDHCcmiHfkeO4M39Dn2aMoTT
Y9mT5loCatN5ypcmSrG3TruHAGqwN3UJqiukGT4NqyntB+dLJfvtuYGe1RW8xG4C
0KdygQQq9F+b2b0KiKLb1/mhE8rScJGUXYjT2elAxWy4Ar/kC72yJr3nwgywoTY6
+Cujo7uOdZ9fBJuDdnS5Y19xIKkgzdIPmg4XIMnNdspQdfKwwfnxo541uwU/m+Xd
iFOZHvIV5+imURsJaflr4EusbJb+VWm7QRP2sOnQZT4nMgPg4IJge8/oOmy3yASN
g++/iGlWPLbEb2pIR1x4xsY3dN/06EI3jSYXSKKousG+CfghO7aXYzM1Ut3omZ2D
npMFpYcUv9LZP7jLx5+RT41+41R+6iTZwot/bRHz5pjfl9cwOnhdysUoGsFpJbiS
u2hu01LejUn3b1zKGQKcDZeuH8SOEUAl1s1MX7vY4F2ep+ifn/RszjGQz5HET1zA
Up9z57sad2KJluCjqdqxZhrG+u279KD8uLMT+/L7tGtAghUoDErWFa4pKpO9Qc9z
wLldssdKTLiYY6EcJQGcJbyZPFVJA4+9SIsc9VpWF0nZ/GtKqqjFw3YiRI1FrStI
2Cwj0KC7ptucRFsWHGdMYmcMixmHiwNMO+dFe95P6q2+jb0N6aI+cxmzYtdQmfqM
vBQunhYRWkmUrh33FZeGIXlJqfoAzPAFDfy7xWTaBnPqtjZOaMmijlHYKFDbpdzs
viuyrUYO5/ugnR24JiSgsTud3jiqg5TYlvFJ8AufF1JX0BhLmtH65vnXpmLNATiW
vcl2F5yM1iKyGMb4sLBixoe5s+aoS0FvmA+x68poVaONyIwnSmgPqgELiqJeJMIn
YdpdGZMEe1ErpJ+F2gbxGlB4xY/JGDMLLUrQfRH0UPOk74QNW3lS6gx9HofvDbv2
IZ0WCnz56+yepTYX6HRpU9bQuomTjTj/Fkq/CbYZLTrPJ2TSucEWSUmBGymYiUR9
is0CFMZEQDL6hzDT+xTe+TpYONSPRH21vdWO+X7hsI84NerDlnAJFewvKr+bzKNM
fukMw+bfwjl5cUDp7OO7yuVTjj5tQaRaq6QzwzmW8WIFVJOWNIAZnuWxQP91f7dF
pqs9ZREktppkD+kr+3LBmrn01abRZWO0Ve5mbeOEAo+QfXrDmFt3LzXLAdYNgTz+
a5/6SNv6FWmcpva6fQQtm4DZhEJy4mrXsQETmM2/30RofcnyDvu2eCcqRPxHr2Iy
UM0mdFyw3NMur3NRZetipltUhKVqZx+kC81LfHg/Z3/thY9BY9X1MRwDr7TacYFJ
o39JLcgFg1UsrbpHKmZQ9GaylvmgjUWd/lKKNJmy4kg1f2c+kF/rpP/OJRpfi3Z9
2MC9J+rDz47YT7dgE6f+hBWbfXoLWPVzRYltDeOb1QmdexP9ZdISFUBKOpR9eT63
CcSljDPZZTSrViDioqidCmj3sUXMcHJFhos7voJ4ofDm7dl1mi6EbB0STpMP6jQV
t3ueO1rjwbX1HP9yRH4WtzS4ptZEgtYGdANlfJtWaOjbpQdBECtJyab2FnxxVTuA
mkr6CSGWPKof/U+Xox0kSrYd22DJ1Xg9kaONIJCjlzeNbKzE6MkKm9/bTU+1uL5g
IXMvEYbjt5AhKvHpDxAB0kF6kQe5PKdHI/waxIaGBU5y5E7Gs1VCbqCEXKJmTz3i
bNk9dyWxLuo9OUGMJ5rEPrNzHqnvNXZH02tGCecx3UjdXnWIjxuIY64RFUWsRF9y
xatH+nmL0lAKbFWcoWelx/PIwENyOwoUfZgSrChpiX7rIFBT1BN1JncelKQoeg/c
RK40QTFPyGlJ0dH5JRXQ2C/xGICGuKFMPbpDc2p1CD3ANGqvlNn9IGu/NpahUIfP
3nBNe+8KgV500glOwBPvaNEgR2UYyCwLlouMFa5UAhBmwH88vCZkmKM9Om4OZDxm
lfdbqL6JU+C4KAF1dD8Tbi85AMhetlnxJGz9R3zrZTmkWKEdoJ/qvtSvYYYg6Ii2
Z4wY3rfD0tJ8UclpMuAjfijPT+sydl9Fy3PDb9cb4elQqxORDKhHgH59z15T8zpC
JScarArzvRL/AySx2DJFtpzYjWpDEiMfR/4yBL/BZJ5Typaq75+ARL6lHfwCipuH
DYcNkh8RzNQa6HdmAq61sTG49eTVmPn7tJ6t5U3S7BtBcXKvrlZ8Sfrw2Wx1nM3u
4r2n6dgiaotkr4iTwmLV9r04nU4OrMa44+Z9SfzX9uKP7XwmolsYj/FKg4JBDPLu
zv18Xca+XLWnKxgxUyk+sbsY9X+y2lmopYFpLIHP+WYcsXiN9u+SEkmZ7I12Wxrq
jijN5Xmv5CwIKUnbw01puV7aaT70U/kFWHOktshGUUJcEzMzhg5gBzw7ivfNe+bN
YZQHz4APl6QVYS8fHv1c1/Lh94W1XhvGnW5MsmXvhT6mBEsNtcQztXqXS9fvdSgz
0BtNEgbNvogIXk+voEAt9h8YQhK4qAgyj0ZQDkN8/vDFVXfSAid4TLhiMVrxXhlG
4mkiPjKYBxrBw9C2MX7OhCYWgSotpejx4SYaV7uHqtYR74y4Yuh4WrUwHWbEXi8E
g+Rx1fBvJZLsrFJuTLMrgQVaku/yrGWvikbCy3cBMJPisgidLrE621LzVHax5oK8
SdtHPfz6hkM66E7iVP9ld637oosBZ3BlsLTFjB/Ayr708oP244KLe7nCzVXrGMIY
J7mt+BxthLsAA3Hy6TUGzdtdkwDvPduA+hNIfr/RoRn80icAPp4qbQm4h4fzIHPP
+r01SDtVUlzhM6J58v4XAQf2Um9BfkvufpxwTmxYSX4/5HT/x4m+duskkwqQ+85d
Ju0PHhoMn/o7SfoCPAh2rywc4QyOzWGKS7jnk7veqn/eVBwvlvQ7IJ1SsKekg7CV
wn+yp7kjyGN+GP6JIbGvWeoCoHM4EzK9k30+fjBCiiY0sHVd6MkVEg0NuS3Dh1rm
jbVFfx1rnuh5MSdgUCsnX6u5NxhqfKKucoc84Ii4aKS3BcDyD+VlIKCr8Itm2DMu
aL2LKuGX/BodVtmGMFifwfvv9Vga1fMeXGyF4iotd3g1orxbxSiNCOO5FCZocpY5
c8wU4GRu+sCcVb9zYW0IzJqheRwbCpf1oibVzsmkZR1o8HC0fWd6Ao1+ta//5xEV
MoGKLwbAoYsbxUsindwuU5eOevL8LzbdlDNW28RsYheO7xxJ85Df+12c7r2b7gvQ
MY7ePY+ryJfiQMO+pes3Jpb4nF+2QTzJ+hn2dwzMb/2ezDLCFrQeJ8ubjXlZLfgL
bLZrQ5PKA4pPPPOmRyC67A/wjsqb6J5KehUTkWrUbnXjXRo+HMOTzkigl8/xxGEu
jVoBxZYJWRd8VNWExM55/F+yUZ2A5pygYPHrfEwkPZtgQQ+8cH2z+JvvMJNJlgUd
71H4pvLVJvxRvAgEYI24gPqeSEiF5Q82ibn4BTVooZj1zvDDNBzBzwOxiZRpxoVk
ZSqLvCosULpkgYKh9tw6braleTRmFT4/o8hO8R2wKO0mLcU6YiYQKZQqQG3Z4gcm
kiJUTtPO9cQNunfqOjrlra7fCjf8CQ58vwG5X75UKsiNsfaHwold6HHu5jDWGnN8
iIZgLLhoEMsipHMhNxfn9psHF4Of5vhkQ+QwYUbp9XNBKaiKdwlE3DD96W92Vfam
2LvPkNmRNPz+uGLco3KT7oOnM6agaAl9YdwgMhHo96PtxuAQsRZf5hfZv+73j5DS
dWEwflw1w4e+VV05sU4otTOtiEraNowxVo2tEnHTA29pfKI5uTxvEmkwvhgyJN77
yhhrx1F/EqL4j6MOSIqQxMhplOmZ8ZvHDbkqiARRt3vCzI78VDyhFDRPoqCVyMv7
3FSeyMWiV4+hzOhcaxtsaI+JPffligioTcccxEcbhn/1iwhM0CBK7J0gRZ5AGmOT
1M3TM2uHp3ZLTFo5YW3aK5MwtMumKdLt7giRk8jq1NZrxy+wDLtpfzjk5opmk+zT
4IDf3PPwpmp/N4hXXAnJx6dl4a+CeeIw/mFap++4ViXYjxR14S3kSnh2yMZPNBsJ
GqvF0WgZ/yeQtM9wIMQLROZYmcLbZ2X1UoWAV6YZPhHJVTW77eaTX/GGOAiPMdNW
k5Qsa5lfh4cb16tdf/YoDVOJRcHaUgc8MhRIYC/6BhKG/EF04Fjvtbi6WUd/rvRt
UdgfgXGqziGPNd7FfMvNq7froRpqEZlQY2jzKvO68qG+9t8gjG5Tm88xxF9ABJFF
bMcwhdtPa2oGFNh93rK1vse3tEeXo5J9uT/4mD2IAUd6Ka7ImQeelUGmL7UtzMrJ
g/DiPxJzgnZqypbcVzAijW8Z4HsCAT6Lw45bf+Q2T8/ISaf5irwD+kiyOi6xyvbj
V2fU3eIdHUY+S82sj35Z3Ympd6AXKY47yNW6od8cQz4az8Xaqa0xD8Eg0yOSUDV0
sjzz3m1PtPiiEDOBwC2xeaGR4sUr0zfyywBHp43U/XXwQXEjvzfuVdsvccDHzIEG
37CMTvAnHrlG9eEe8aX3FGJkvNClJrMXYw6WCo5sWMkGfVB0voC14lCNrj/W9Yql
4aKxRL9/iOlB326BPbQuQPuM09Nq2WNFxYu5tDcpug7ODQDGs4eLBw4XuxpUSvuv
hFirc39I6Rl0Aj6MBHBMmFgMlrtyeiToIEPpAr+hIzM6I3eFQ+E7cEkOWULXxGFI
2M0ZymYfb6WC6QlzUEDDvw2Nqz+R8armhKUb/wB29Z56gZFfXUJyzVKNODQr/pZl
7DggOpNVd4pDZn6ZziAauxMcL8Mbz4KURX6MyU1NTsJPntOenv+wPrmP4NZVc1NY
XpMdzcz2cU/Jb2ReH6vxFGQ5TwZoPz+HsY3+V+fmNUlVXu8drCmiM6e5zbrIKPq+
JfwVZ7Dz7qI+CqKkqvYwwC7wHWF5AaFJRSp7nqS6SmZG1eVEPp5RiWxVP2Jwu+aE
w1xYHWeYR1rNoCTcy62Gn6vxJ+Mq9EsN4IQTIlJhjpVwxlmGxrqBHYbmk/gnXr6f
3dM1IZ7fnUM2Z4LbtJ9TdpVB0p7Qspchm/7QuI9XkDxPLuOpE+FjJXlpqOUjCKJp
o7Yvgz3FfBbMhac0Hs1+NS/EwuW6X5biTazb3ITv5i+BjY0ay/MZsfy5tCEZdC/d
m9sCL6rzOJIwcxgQ/RZzV9mgE6SoyIUeQ/I55X3HictprDjNXs0XwCq1JbN9XCMS
UDipDmOa1k6jIOqV/jWGIiZGVOUbcJ6A++XGoLo9F9WwwKEqT7z/BiQXzr7Ksf+7
h+kPQhxcv2HVE4V6XMeWD7w7FYQJijkTnATzvkztk1v9vvgIDeoyk78wV2hcQFYC
T0+6kc5veA+4oPK597RGb4utEAs3FCD1Ay/tsofLbXJxeWXAUTBUnO35/cAlJopX
47LVxAT4OYI+rSO1IkOhdlhv7vrEQ43pLAFc7BG+oUfLiq12p/8OWpQg5l9oRot2
xbBwNApr3lrHP+SMwuTOF16ueFbe4cesovrKS6ryVVk+aWjgXcdkoGgfLOGjfQuI
91rCSo+AWaFxif6wyb4TRzaFr3j5VCyBFIOPZ9WKcvK5sn8s/HgEwddwlhlptMje
6EsPTlOoYRecZTK01C+lpRy2R3BJApgnKJoH7uvuWRGW6cgvmzOSSO9+Vs5rR8hA
q3Wy0uaXb2YL9UPEFJhWqLppieJBnyXTFWeWupiqSwItQ1FqF0tqWoUiOomKjgQM
gx9ZgEBQA1a/d9J+lD0ONwxhksdz1HmrrMNmnw01N7s85DMj3v/B8bfGtcTI7Fj/
j7dcQsn+DS7j7edvRBfFl4/TFXa+lff4aO+cDJgZFqlPkP/F5JUhfGZJkdqSTTSr
xMRTW/TGKq7VJhsVvYCTVH5CeEYC+qLidyNfZGDjhbR7GuVWSIhvd9S4NES6J/Dq
jkVDyR7LXK3EnA4jRF/m5Mz1LSSnf8c0+pi8y15R6cC+sY/F0F9R059UdfzLUsMF
N8PVcz6PZk2tUUSH9+b7gVIYddrDkFu18W7yA7rtYs/mrirLLOTxmqJKyyfS4PI1
T8AmIaFDf+Y9z851oi2O4PVePE/XSRGVHoSTXJN7/y6t7sT8G9CUdEl3/VzED0gI
uIDnnt0sXKW+nyJiYB0jTvUkqJyjLhvRBXengc7pjq018+lpI1xnt+7zEFYCNXr9
iGgMwVn+w9FPePjbrKY0oq0GfQUfJ6jUnOe0BPr4E2f2QrAAIFuH/Lzz1zKINTzT
sc856EudOdXndbvJVG3jODOCPTxUcbvTYTrj8IRaXIegE0eNFfQJKjLU1uAFgqNg
r2F2jBjuWkeClzx/m1KcywmNA4l8kbyjrUOQBuKSI+BuHuGR+//mW1/2EZmmYO1y
fFB6qfEblFkl8jzzUO4Yp6pUaCogawkt7GgX2vYSwppre4tZOyfCo+z7q3wK7Poa
GILvFqjROCrgDUNDxoUoSP+qi+CGKFeq41ij3Bl5Nsjk8Jb6okn4Ft9P6jXIwUoG
JGeqdecRCgMX/vm8k6k3kQZn45/8bJrLLnqxr90Oi41hzIh8MJ0gWcz0psrYOcpE
oj7wfMDcfX/GYHC5V/LC7fkGP3lcZtwqP0E3lrvqk3PIXZI+PVIP40jF5CrV36DW
vQJdlPGgD7anrKulCb1dPRuqR/puvzdg/QtaYQp6EUsVqsVLuzDs+xfUiFc1vH9D
UHoPLC1cnuRaYWCq68xRW7Ko6KhniLgDCarLv7GJkzbBf6Pg966aPk3R8HnaFysk
eRbpLhVpSs3FH5s3YQmPdvfpWXqcZtlGn/mNbio54wm19gGjdXXTCrJn8QK7IqfP
X/sZknKiilvugpEze0L4O0uec9gbQBwOFMUdyGZEKdhps+4s3LH/j3SZ7JQ1k8u9
OHedZw28mmaPJR42+PLpQm2mSebsM3WJJFJsjXPwlskiTPUYJCOn+uKGkj/vHu3l
kqSFHh+UxENjvF9wuGzk6Se5cEziyKK3P7z1+3TzWwf6foUUneqFn8EJnDWq5EfE
9blMuLhynK9SvZ+E/vl7QCZDiAi9o/XEBx4pVu7AV3bmVSAnJYfMrtI38XLrpqmG
6ZJc5Gc9bOQdOhq9F9eCNNyvr9EKPoDiSiQu51Ar+7DA0VaUb4aUgDPJ07CeRUln
PDEgERdrij7v15vszeQ77BctsDHTmBxa77/2TvdX9nH8AQpd0blue46W/sUJgNIh
6aAYSis1G8/iue9RxPInRFigUrx/Dqh/ezIDDAThjtVz54Sxtq7b5FDLqtHcMJ7Y
DpNGjUdzpyW6xuirG3PBq+hQ831yAInNSFuazm3aj7SHBn06kLWx/8Qy8Bbdr1uQ
/YDt2BIPgs5GxIIkVqpiz8CmbN2oxmabHoVHQiy5aF3OMVkn2wa7HTemyA27Fz2P
glsvhHme3N826lWUZVWRhI2zeUy8ndcIuFN7/662MnEtl4TsgOLtWDbGjzDT8hLO
2Ufsma2fchTdr/yvrCdw/Z3ZP6a6UPFa+E+dPBXex15z0l1owedwnFUnFeZTtOEV
pojt5er7CVk+AGCYBFbhe0/kt8GdfOuFvaBt+NzibB8kd84rgEbb/OM706mT3Aeu
rmRsqxo/fWpEiFJvWQvwrYIYWwsdgaUp39xfyNom8e1Ks2/Y8jWmFnNGGBYlCnuS
rtCmJ9PDT9ffPOx5w2aQxyiuvfj0YI1ngohcaeJtVHC9M6XXQ+w288fak/Fgk3Dx
HV3mbuNTXUCz20CB7PuhINuZeGzT1lbyjisvd3ZXjjc68Dwxwp341KboTML++gKD
sV34ss+DA8/W57zZNMjxDFzKZBy+fvd+c92HUkWr7/ZgTM8XjRXr+/VMBiYF0+z1
9tirktU0Q3pDRoRy6KMg3a5hVKQUTgqYDh+L6K28hUOxXAV+zZCxBE9n1s2Vv3w6
vVF+K1+hELSMN68LsQVg1LV7tIgc7bDNVVD4/n31mDeUPS+cutiW9AbZJoqAwomF
9Tw5fvFXlOUtqGIHsQ1rqMgRmVNr1qWgOJ+1Aco95dCD6K9rbY5KKgTlCgz1OnKS
VXFwmQsi4ZYvDrbNBkwOX6FhGy3tRJzULtxvcy/hE8pHoSOfDLTqIWNuYwxW6EWU
bwLjkpgBpLuJJ+KCPaC4DvZMBpVAXjDcoSor8Z0ZYWHbFJaodoxIYG4Q3TrAA6ba
0tBPfCJeTe665pcIcd42FO4QnsN4mvG2ZNQKGperNT0VACT2iBGSfpz7CnL/M9My
bpiBXhnoz0oUnDfk/B0ZUqw8Yf7JqO+bOjtXCS4an2dUzZkoUuKylu7Awoo6Rigv
E9i/oPecebmhlbpOWisM/ryUMzKPVjbWpBMwsdYaAHFZdMBlBeVMkkv13gwTafwn
Zk1LfZs8/awd/GC5Xq2wSgXAb6oAUzZ51YV4Lmw+Tb6gEzSiCXg/fk10QlPLZVCF
URX4E8DRZiFRA4bzmGqXEHqeNmMm+4WwWPHiboQ4lINcFRw6ZSh2ur6kt1fKeKK/
YlYLrgKjQX5bbLmRkzM8hyX3vQjHNav8g8Ppsca0sqBOyfAHG2N3+yfgLkrXeQWR
4drh6RzCe0NJjVXNrKi4J2HJKT1ExBb/hl2MCtB0EnJOeUq2+tPxZAHeYN4mQpVU
lMFr545apoX2NxQOV2j0MaX5SQyOkTKSPMlx24t0EImfSqIixcwFHNb/Flx341ZB
BKibny9nM61bqrhO6spoMeNJDaYYSx0hD28pTUPsIx6TvijOXpzgXk+hQMZ3L3B+
JPB9HQFVxHIwgOTB4kRf/A6MrOzRj7sGCQ+5izX52uDX/u3aakZ8jFsYzG5l1hYb
ZGZzjTJwWb6/SBEHVZMz7tifcfS71b6DkRwwbk0dU6QqVq+ef/4gnkFzTlH465F8
3eaAWx7ZqfX1oZSP12LU+tynKKi5kOr6OgomgMq09b6SNN2G1u1t11Q7Q+WPMqcj
960e1/YZVriOGNaiiGLBFiBEovuX5/rA2OmYnloHP5Lteg3jUBcplKouSHWMGJcr
WgjkcUYdVJgPX52Ur6QpNEKWQsAKpf+VMnWDficFN7eBQCDEMej2yvLc+SBYJQ4x
qLkTRVl6NLyevk1un7mPgmL/h9mSdtGPilhb3Dns1KXVvT9i9Lj1klpwM7kCVo4e
/54SdspscX3Wnszvz8JJsNQ8B5MVnprpxmbVirXwwXc0qkqpAe7pioEtLq1KDJm7
P/ZZ/YiYCLN3Q+F/ykyhH3uFSakDWgVQ0zadYW10X/FVSPAulLb0Cwrm/0vmBJeU
QEpqx699O6miVAd65tUKhpXIyZ9NBIedYu5kr4Fj3Qqi8WrCExPawbTU1N/G826r
yyWAL23tdeUu8A1CQR1Q+/gK97ynFZojCsZpUfR5qyNyl5oV1CIIrcAr+x++Yf5p
WL5dyGgEe0LKUKmPqL4ARvHWkdruAaCSDtN8MdkhZzdQBUunco9yDJa6vm6z8JMT
B7u2iwaI1FqmTyB2Q0rGJUZ3DxjJWKJ4OLE2PjqJUmRDZlkXKK3PYEhGbzsqppt9
+cRqDuyfTEr5AwN2EP0HWwQdogxL+oepU4b9vL77yG1eWepymjJR3J2tPeCW1tCM
ZdpdNVuu+I3VX3hQPlKz56CdsLe7d2mb9F/ya0UrLbaAw6+ByKwSZcGYiv6gmtmj
xOjnKDIY7edbzLjCRixLKEjDAavB16TofSrUPkc9JNTwQZCv2meEGRP5aT9eqFxE
6ZEne3PBZvN8GF0j1vfq+tOYqT9msJRsGAzuXql+kVDiqu1HexHAlBQkMeQNdUM+
nijAPSBfePY92Gd7+Yh/UG1us2upp4/EbSWOhI/RRM73s6Tx5UE4W7nSc8rFKw/p
/dtVw61uM/FjjOuxMQR44l3XC7fdkHKhaH21a5V/9aL7QiuCoqdHxv8piYODWfeN
qCvxrGzmksq7eFdFwNqVxQTYOC1JpZzFEhOB5W91K0C3Ymq5mMLQk5wt5xemDx9U
ol6XpN/eICKFFv/cg964p/KCOQK0/y5LHCqXCM4JEHa2lmPKuol4M2UCnIlSowpi
tBLJuf2UUfKyZRAi2rbbCLumKskytPscc72JBTkxDJJYBrOvsNN5E/XQgF08iEvW
361YvuUExeN9VL2GOSqKKmV2voKEkJtiaFsTsw26VNzxFNgZjxEXswA7wCip9o96
yN1ikY6Q0IQoqmS+t9Ffpd5Ya7nfqYHzd+3nsgNIr9njo22ZCQ4rEag/z1xCBHQb
y0hP/tWxc3KBDp16sJeBuzMh+44ohpNL24wA075QNz+K6LnU8z6KI6lThv2bOsvO
VCtPCSyrw874Fan8+B2xQOVkBwRvAwL20OP48N0KTr6PIxM+zP79H4uVMbcNx46P
jbeeDBp/JxP8drvGeWqted76xj9l7aGNYa+SfDfBBOfyYx6novDWrQNSP204T9x0
3WzYxBd/TYGRq5kqRtxoAdWqtbG039sK7oUd2nSLnKa3x9u40l7l+skuM4xgLDuG
+5Qa1VqwEgaTFicJpNra13derxsq3Tm/zHGS7OM+CYHUDsbcB+vdOSfC5NKZtv/t
xYKUvWySQCl7Z7LLJg3iY0wasfvCjtENBVjxUhRUb38HglZsNrpq53vA+v9Q6YVh
qB5rUlnktJEekkA8IWKcK9xUQF8NAnGDD87gOaDOnxeD83GnIbqp+agx+sw1n5UY
jyqrHGYHZN2cLbn5VvBVbeuP2b3UEYMoKb6wOpAfKvLEy6Qh+Ugh5pv3MmJw7BXj
pxQCihaPrxpjgKY8wPsHVSwOyKhdIbc/zgZYCJIfvdCf8uDCxnEREbsSXA/oqqSh
fXFaPf3UbTYTldzaif70gws5mSjFRqADp3TJDEM15DVZV5dUammw1516FCy4Gh7R
WwSGwnd0AdTSIpNjSahnoSkUVTrLRPdnsrbUFkIEgRNlyRrAMCDGe1W/QW4dFXHG
KEhArpBcc+8SNs9nH983GKzvcxZPHfX22G4JKgTrXFy4JYxHE3UaI20EXru033/O
UwK0iSUK5MulyN278uleGpvyrYuNxBkQjXWZETPgcIkKIfUBAEb3RfKVGmxXjYSp
5sjvu2/SqUdhhyNTpf6cUnIIwz3t6gPaDjLpUpTX9AeUT2fk+3c6+8IZY+YQAd1e
yna1rkpqC9JMc4R7eIEUZEg0xCuXguVboWVD6Y51UmNv6IZJrrGccLmrEhXd4wLD
2WOG9Pu1DWtz8zK1RSh+iLrsn8POG7AbzII8Nj1ph1RHpdfr1p6LSVqwR8+Vtqdy
3+mfjsLcDcfzdTOgVUAh/9reshtYeZDqVjC3OnseWvZFcmr2TIX8Ro+lLVVMA5kH
Zi1Grxk6T/A6D6OkyzbQAGyEgwAFwlUkNUUTQ8NUnkOMHUlLEYm180XHxCu3tAwB
Lp8QWpOS7U4HslpmS3FreZth9K/+e/E9xs99BwNHUlsT7Tyx8AW/e3eFVoo0uUjR
od06qO4zlxm4xVFGlty6Kn4dz8ZMmdMtbex+tZr/lgMGEuDxUPwVcum19tx+1XmF
8hXAelV6F6jyl+ifIKv+Lu4+nvBHSEhT6YDyiYxNVAhaHLZJ52EKW46iAXyCidxj
ivrXanXi42ttqXh8JPxRjDvWw0AGCag4+5L/lCAOTO2xWzhzVfpHA/ui4t9XuYBa
H8xOLBRKgi9xX7WXD1ENfRluVN2/uHAxvvZwUMRRdXHgfZN4EQ0ga6xgcOX00hQb
MWC2lHwzGuhBUr90SMHptodTx9v8zOqsJzA7mzz82jMerQNxi5p1y9BqkLuc74om
6ilCxkji+8EDdciPLI7LTSFRafhpkGVvGyDUxJ7Ys7vKJ9BuPC+l/2/RU6HA3aMw
1syrfrgzOvDRhTHPGc5/voF+StJ/f5OTCBTJMR8Yt/vK7dSWgcqfZBeZy9cuj/6X
36ut9ZZIa+tkB3TFUurCvSOMrA9hadFKcxwGobcuCawGU/zAOOj/Iq4xcIfpRlss
mJcNnQKSHqDkk/n+yW16DH1ZrLjC9bKWUldoKEWUvcIV9dXiVDMn2bkRnZO0HPoQ
wDENo5Kt2kVUJEEhdyVM4PXK6fjilZezvS3oeBM3l/ovMbFViFU3sMl3hADKbcCl
SE9NntjQbp59K8DXnikGyggF1/O9eYsAlH+MSPHvtkWIV2G+cYTe2WX5Mnq7IhuG
xWkY5tjZpjAj6CCHXbCPErCqpNfdYiOqK81xwJr5XZhFignF/TG3Bop8fkDM6D7L
uM75OSpXNJYCKUu/zXEh6Odk4OG+5+mIqM1bHVnJ3DQAfn2N1FOHJFQMBWjuexce
wOe8AOkvTxnMfCgW9dU5w3TNbu7mdlkZ1pwGzw1SagwrswWtxYEslDnQX3jqad6k
aejMBHzjEGbj23iL2hVxU/pqe+Zs4TQQo8vFkc39OM/PQT+xvz81DO0TwtQD9kYg
w3pYDir0vq2YMSDrio9uUqLKfXVLs0xgDuNdc5nsAMdHGTA0HyLhe5GLtUr77cFf
xuNzCmkGt02jnziu2MFvB41KT59c/0GYLtRop40mI4nzIgWFVv+XN85rV+DqdGFu
6Ia5J8RhPIQpjjs9ZL3SMs0NOtfRMaQtjzqf8m3jptn8YMO63jdqDZEksoGDDIzV
RA6pjNl+59XOww+Mou+ZWTkAt4jNj93lvKi3wGW7bRGGYt5oytkhUlI2782465u7
R3YfFtWN7iDTGj9l02Cxiyg1tGDfXF8D+V/aWWFXzfx95ii+/oWAGeuKMy3HKI31
gOnBEHHh8ph3xIYjuYiPO/hK1RaJ47VrGIw4HsKUQUTm2vyfeqZIcMRkNrSA7Zk4
cwYwhnlHFvGj6keUS5Dy8NJRkSjzL6wnEcvU0zUiVfSANAEDKxgJUzWATsamrPYA
NmF6TMoESTh5lbmZ+MF/rDcwIJO3bVprqOi4qOG4rBSo+JOTSHvfe5zW7p9dz7jV
NJKJn9G3jkfgdBaTJxEUhbzAH3o2fO4JkduktHs/2Qp9Uou8XWagqh1Gl/3wg4Jh
fs7AUcuLMgKz5Jxm16szHQfDv76DzQDU7dbo4fP+W1oV2PdQapn+rrgS7m2OV4Vz
tRrfoN8Zv2XaDJFjVSBsRyxmH2V1v0Go5ogDAVDcX6eBDdytDDSUXYEky7QI4682
tLDxgeCSRzXJ0zvukGVRFslCJMGi/pvXD4QQoiXwgj73fEdQLnY1cGOv/4xgRyrw
x/Sx0c5ZyUVO2fSSjoFPHiH6U4955k5tFm9CWAH9tSnqhTfxQYbpcVfoYAHYkGwq
fONOWZES9fYAaNxMmxd5thrDb82nqUPHGaRZ6HqYY8UBAVyl6wJMoNMrSpXpXwZw
jd32QcgaR8agoTFxczt9pW2rJ1W3v/aige6ea7u/0L9q6gAuAOPUP989mfa5YiGS
ahzu+BtiSFebKkBMtkNN0s881f4xkvEOSdlFe9NbB7YMcFPFBdB9sYewZLgQLQ4C
GJJSs+faFadEbxbhkGyH5TqO7qsQC4r/uvxG/Ssk9nokrRf3C1MeAznNVa+4R6Hf
0eyPC98hZ7sfBwKTJDn2lleWwGCZ64TzHn4iS06iKvbU5TSKMsgGr3vO4m/ZVPqV
PbotQbClBKE6yBXu30CdaXAP1wfu6jsCjU0qlouPRqTaNp+ywPtgeWUwkLif0YUs
bBVR16FTdxbHKAdsjHOdHQGAr2HnpaIWOnke0FnhoxNud+LGT4CvlbXHEFOJR17Y
La/+T5e+RrIIWaH2xVZLNRGLYeBoPObwADrtF9iYKpMRbllKidXF5Z5LxgoUhGsQ
57Lti0b46h6XhneMecuzWoWxYkaTu6XA80gkwyEFQNCclaoCgA791TXKwJe+w168
90LBT0OqiOlon9/O4CuJQ3vUuCFpM75rcH/5e01nA+KQxGFRJXQ2H4BEnvOyHrGZ
3waTFNYJ/o+zv7WIPZOxHigOQ9qsZrMfUlOYEcLa0XSdgstSnEspq6n2mbxyATHQ
Eigr8v1dD87IbofoVZj4ODKf9E/vlRcdrvG+J0BdY6fKXvWXVuzdTUk+n1jgw8sh
OxM9DoT267c+hdHA1TxKDB+yLdPjY0ZU/wN4ETwuLdRALdqlIz8ap1s46SfuDgg8
NDVDKhT+6B4IPxRrxOekD8/20a+h2zWckYFq8J5w9pOBhgnUuSv8ZhyAxZnW/Irh
+imbyxTaDrS0H72Vdnqw3cySlAzyWKiDDHmxo0gnoF0biIsS3wThoC255/8T+rOG
2mEXPyotc2/9PbUyQLEDt+FD7sFFcHxLaUSMW2GJaRDa0pSFRRaJ9d/JN45kJ6VW
8/RjSkRRxD7WSMK7fAr0DK8fIBjNJpItaq8jPNGwEvxInLlJ13IArOSga9R2oxzm
nz7cQ/eMJTpke5N3YxEkHee6RS0yjkQsXgfKCjK/T3Zd1jLIF78nYiWH3+9VkEyy
Pef9mJc0NiyNADBCbPMGZof+oCEUJBMxAC2Lo6fQeygxT6dgDNg76GaCxtBj9Lv5
u2lnEs7XO96TCSGpzU5zKjinpdVQ86tSq6+iIsHGesZdGLj/MzPLZbUQnTx6N8nr
4vi11mj8JA92jTAGbaxeTRD24zY8hOxIi6QZf1jWXsO4QYThO6bBjOWZX8g6qZha
/x6MRu2NeXVtwsFodSFKIMQnhzItg+17JTiw2rWGslUwXRlfP3zy7uFdzFMB/Ltu
RLqntFZJ5IJVmw/ysAKY68C7emUtwbAp966ynkD+HFLJqs7OnetJFYgEO6nZGhHm
3TdqWy+UqtQghG4rFv0Y5Z2dki/sipe6DO7HhknNogF9NCSl9yZukfonZ3ALRe4V
N1nZgafNWCag7bEgRM9Z7tRIBF5uWLs21+hXmDeKYjii7iTATyhlByUEx1Vb8CPG
MiTOgUkvu2z67vbEQJ5wCwicg5p/mRen5WJ0hrz1Qx/MrLjHxZUlyTulz2rZvNRY
bd2ZBR1dI49zdYVimfVS5h13LX4lddxViFdoQnX/AVqkBT9Z4XgmKyi8irLpgnUV
pjcLrhsQIcpaYNKFdnWknqw+Oxm5BoNNvVMmyUoFNXr1iCx0hj6TqCjaNEErXuS0
gtMzLuTTaaHqisRsID058kghwqSvMrSBUCG6FsOl8qEx6Zx4A61UsLJX/gP9cXLc
NwOm8qfxoHtKTK34x1NhfhQ6q1czPzmot6Bk6KXl6JFBydisoiA9yoAIOCEyWXd0
Ijb2cIiwiQvEDeQHFnCvAHfM4uyTcuN0ReT+utt+63ghFMQsQRsY0XJSbG8GmToq
JKNltG3tTPqgd8y4bvjSwzcWTlBkNqHrkaKYw00XPL531cOFgvjR7/gUfBbQJPat
c3ug6HeSJwgO+Pi2+7afDZEFEYm9r2RxG32p4sAL4U7QWsmewjY4m4EJHnoWGmNM
R2HcQ9vSRLWV+yNkVRXAvNoE1ob6BuIrzgpTFvzt3cBdcQ9r/UCFTIKbrPrT7/0q
75ugtvVaRh+PgkaqsxFFE1Bm+AchS+M0f+PzSt9xRozDniwtxAYuGDmpAxRdS1oh
OZdL8zgfHY/kHC5DUt41rpPBMTIgUOMkkkyJqV4EpJy35U57QKViqhMKTakbjYt1
ZuR7ihIG3RDrbqZec7RI7wBpyn0Ze8AfshhLFjFp+GNn1BSMVZ5lSqWG2I5VgTSG
pRMwiltKPHdYXX6o4mw1s7V3xi7RXbnqSLOqEXyXlEdmfV19kiDN+ysG5f0hZPYf
IjjaehrCk7qxMbm5pO49ZHENkt03lPLU0s536ekiRGd43q1D1qCltAbI2jU/giCQ
Fo6JW/Syu+MIvdzApW0Dxg3U7ggcjfXcOMwKWC1jSWhpegjzEzQQZKCctnyB6F7b
Sau9z5FEdIfo50aYQ0E+DWldLnkIbZbui4thxCGi/Fv8GvAP1NVeDpxpDA3aTtrO
twB+Ys0KiqIRMm/gJ5c8ogE3Tgt9y6JIkYpGeugTHVg2gI2m9La/WxP74NZWd5GD
OIqAUsxk9IILDZZZ1igaKo+HetYNXtNnQPTD41yNsi05PZ3bO4Y31u2Dh8fTYD4F
bmY20fhK1ysKSIfOEZdNL9GLfHaBBV2AWnKmiKEDeO7LSUF4zmbXZpi/HBCNrTSC
VdcoUCCB4VRiNmf690iArAs971rdRLkpyHdd6eT9N+zBSpPiRhE7x70+eb6vlu81
ilMuCVlv4J+LN9GrZBg6gkPFgN1VUpc4FzgKxVS4TpEdpgP+0XrjSiuRSpikA4MK
tkDT5MgDdWhiB9w0f3maRi0AVH4I/OpBzd/SHhmj4Q+2F1msPVkKrCod/BRi0Aa4
lUC4USanygzZ/omFYDtZwVi+QutdSfIYTqcarOHM6gEyOs3gub5pLzpMDh9luY1p
8EuHFl2G+507fqs/uE9eamw5aqz1EiksvN6Ijr5Z+e4OfakO7koOo1lgqlsUU9FE
WNvAq4CbAmW/6yDdgC0J3y1lPbSsiriK72fVP7I7JDjN8zX6FKCSFY2nxYexy3n8
ipn5vVp1qo/cZ3H0VB1xEIxD+C3usrZqcvlkilywPtgoI3zv82ZrsMv/E6Q2v4mc
H6Mxw08dc852XXLUaGuybbSxGIg4+fdszAIEgRcd5+ZfhgWhQecQrc5poxbgrPeb
jPa21T89Zqu71PXY2AAKj1wT7eTsAvUXXR+XVlMKPSoUzNSqAkFATcImECV8QKsc
iXw2c6koB/ScKxii73pDGnO9jfSyNDFMDsy7FjSXA+693/SS3IopwwfZcI/WV8nM
7jMXFvI5EhN7MX2urKPXwLZRfWEgvZifzGqnhXTMPA/9LBH0pIJwHHcOcG376h+H
onL7Cz9yOkN6MzWOsxFrA/z/tuS3BjUh8CE6YzAwKadZXYmk07Ey9wfsZeTeXQLC
z88TYztkCDl2mQiwC0uEpVNlyvO9xiI5rd0p/uDSIV5AYtdLBQm0vMEjdp+doiDC
feSwBNIri4fph5JbojM3MF8Ndc3cllqDAblTgEQObbyO2Z1nJ6XYi21LQyJq0rMd
vSq02yMig2rDNDq7UJO4PvTEJNPXAo46rvSGp3s7hARrkQx3oyBRN1oSleDGZAT2
FdKMOHQvfhjdxLBTP5IomPabc2/qtBM7+ASwr83CHQvKFr+z7UowCLCZVK9tRFVh
dTp2eQ4SH8JP50SB/4Rb1lXBNz7f2qKVuvx2I1+n/I/Vx82joalbf0DbGl4DLtI+
OwcLu1eYCwdIe6nvI7CQouSfjRPpb0v7s0ErY1erTbHUciG8kBSMauIO9R4zdu4t
PkragyDpNiolTnFyJbJtD5sLYspJ/Dziv1V03aHaMbtliGn+bHnAv+YE/xxGGgn3
B5dJhmWk1sgUrn5wSPToZ9yf0fwZmBRl5mjHGVno47eaHpsjM34og6MuDnP8PsYh
QcAdIT4qByd609JFr6BB2i3xT2YtzOVLQ0SV2/ZM6iaLRdBmS84Cfv/iow5o92Ci
/nLwvA8/pN/vIHqSHe0wXwo0/BfJefZnn2xIoOSE3DUeJxCpnKxoPbwOd+t/98gI
QzACZ+bCo0qpsaXqXG6fFjQQO9DtxpKZrsn3eNT1LbDKEw69nZcNSfUWyqCQXuAc
A03O7IcHCPS/iepxJUzN4QGomnm2C30SHZ8mQvmNicDhiFucVDdllWH8mtTZBN6I
avNqpNp58YNnVKEM6DYfHjJCCwtaMtJ44eFK+A//IL46+nf6KQDe3ANYBturtfaP
F8XnW5GSmS5K/SweUDLkaTRZLDsfAtmEkZBfvLEQVP7Z8ABzXeMc9x7+A/CX7POw
dDGe8w8HEqb562TuyNo8APKFpWxS95mGebhbH9k3XHcjxKvNrUgHJQBjH4Tj0F9r
SH+N+nmB+imHTDS6ifOQ97UyG4HRI1pxhlNZmFw1QdHna6htlQazC2FYW+19YQtb
58PJpNGozhFZMU1go9b3BuWaybsuwzyS3ZqBTsbTM0keX1/e/BqoLiOIlsfFnJuw
reRXdgs5zMhKwhkBIF0LI5vIrVxYdPJ23KXl9YOw7XKsn4BOCowzhgSKScplrCXv
GbKWYJ69HIc/+skl+pBjNKfj7uyKlYdJA16xzDXssJbH8GTsCdnF1Llj1tqg09Md
I7fS4hIdNqd8xz+c4VgNCabyRGU8LqIY1sDVJFhOI9iPO9bf6UqPc+Ix618tcuMt
Q1iLr4zD6Q7hT/NtF1Q3UOBpBTsDmj54K0rPw0KxbLelvAG/k8md+lx+Zz1PFJuh
LcKfwBKItctTcSdaDmzp/XRUtK6Ik5vqccZOJs64jSVriFQwvP8tpdgAMzmbKqL1
qP9Ufuq8Emr3az6HcWIUOJZruJICcHoNOHCNc2EKiw4R07UyhBm4zwiC++M4zAM0
KDT+btL8t97SUiBYqpHqNrs9s5Q+JVVjb3tK1bPF7XU9I7F8o6CMUB3+ytw8hygM
JQQzbb2XU0l1wl8CkAR6hV34C1o7YQ1is8cnBJGAFR9vV65SRoNOYPdPHPq5sZx2
GrzzfqjPuvMlVms/iSHeLOQljjfjlVjy7qNjMPgX9GK2jP/lFkeJLf02QATTeS2/
JMfYdM3rEWq+OXA6spneycF3CK61if+YsUEZp6v3e7ecoW+ig/QasnDHzB72YSp/
kFeAIEC6QCO5R3HKopj2oDKR6qT3Efr0RyeWDllyd71EgV0A5QAeekK9xl1VVvg/
+8reg+6zccPSlMuwZHlx4VsvGNPtDpX0ARy3NanHPs+LUa99fuKFLbrJrty3BJjR
Hvx5A/bI/Z3KIoUltUun3KOX80WIpQPFDvP0KqY4orrjRenjo5xLiRDOokmOEtbX
B3poOhpdIOB6H3cvl3VYCHcfK1ysD17kJBf1qIKzIf81HRhH9wSpbYdvtNZmJQ8y
+G87AEey0JWY7i0JAnJnNaoGyZNTUSCusbgHdvem1qDPdWFveg/trxEzd6T8fuQ7
4amKyT1kR2tfZFPnJdN5/ae1yd5OCjdvI0T59glleRPU/yrBSqmSZRD8SNkN8+oj
xPMzcqQDvfZLix+LTf9dnyfvwrW8yx/N7iz0MLu4Jply3zE6u5HKZGf8iL4KRNJY
t35C9zDPHcmvnAlRpvqOhl1WL9c16l2h5vHrX2M8+F1eL2DcK0fl5zcTTusHY5c2
y+JVp1ryDyIUY7hXtt//WHD3jmR4PEBWeZnd9fmo3pu/IbXe8+7oLYvNBWzcd/3M
kUI7/3/47nb/+iJ5VYs7Tgj7KShYqtplukD4tVxbf4QXfNqrKwtqaUp5EOo6MSMJ
XXTJjGrf1ZHg6qs8/AXzmlingz7k5pqIVBOT0XdUhToUYaF8mVweqCGFXNvKKTY3
v5/IYftzGdq1ccdmybw94nm+uNya3tm2B1mt135xkDH7YhvOxI4sw1/U22mMo0me
P4XH27rH7mpnEWN2yCGxEAVFu1DXKVPtWw49CbNHy6KWivZdXAwekJgi5olZQIQD
Q1N6czXiiZrGyJEz0CWDTQJ/fcvJ45f0Bl4cZzmcR2TLCIzt4IyoA1Arb8p3DB1s
l5SqE2mLz7KeVTiTGSFulBwvPxRcHjFxQf13zyXQum0yJei5HFxUhrdRsqWnJctc
fmuFqTRIMspXvDyl75Mp48A4urGv1H2QsEXqvQ2v7zoogafRJOf2rdbBqmio3FXb
Td1t1Z+j5NO4h0ieKISmaAIbat9FRGZ/n5qVufGNHRFFItrY+ShT+j0zQgwKtmgu
xW3m7NN3cLyNmA9mhgXq629Q4XsEzERU7x1tbYUd5p0/q7wcKb0Z5Utn/o03nwHc
GgvH67ZdP0lAcMn2O+K3uLkO0FaH1TDf31PQDa1Mj6RGSO/9GY9ycbLaarfe5nwf
A/Aqy6JdzW2LmIKFTsIBruBdXNmSuQ0tkwqeCczVD2oG6FmffOuzK+IyyKPLzoWE
8Z8rVfzmsp+SbMvecCXXKhpqDejm37/VbRWPWP5t4EbxaD2k+hCeDuEniK6S5w1i
Sw5zy01QQPWw0eevoH7hXgAkKSCH6I6ABik37iLYQ/8MWs+qXVpdhvqSp+fhgJey
Yul4WZmqNTNLsu1XskMvNnrj96FKxUX+9GrkCZ/tsoNKOgrSRKqgxzibjX9CX+CX
BirKdODUSpp+lem+cg/VMREyh0YxABtN3FyJMg8EXAeJUUVCb0LtR4Kzy5nl6Kdb
9H0kHRnHQDDMObzA/USZHQxQYzN9RKWX009kbh3oQx5FbDwGiMyTir4LYPtEnh3t
mJr6DaNhziHdsKo3MRrDwcQqdz5yLkKB5936xoH+Ah+oOElkWpdNzTKDlwbz5osO
FCn4Xg78UfgKvdho7bNn+dvvoi7fdyI5S3sQkq1lOJ9UrUqgNsRPbny8tUDRYwSv
Xqh/CICy9+yU9BhR31z5Xx1R+dHWApMnNjxCJcRmm7A8LPi/ROU0FESS/wuwhPby
+GSc0qc95cvr7hyE3XgbF7QBrj67s7MTbYyNylhcUN4jd1fpYzJvk4G+isc0ehCd
fThgBv8kNq6BkG2nBmSTOQZ8B35RjM3CgkV5JWXLi2nN483plBcluM5LQZenSDgq
DgDb0U/GkP3UC/uunPoS/JKtypt0DErFVT5f5L/grSUi4m9ELUm6LUyl3f5z/WAS
xgUQ54/w3qTm2s8RfN00LlCSotxrXXFXjuzQj6SbBZhIHEp4Pxy8PZg1rwaKsfcW
a2fVBbOFG8gkoboZy8BfrsApW+Vgpwhps1i9nf145pGRbmhiQ/tWzU0TjigcCEEH
yOkEldKQQOgJWJuqaqJnQJF88Sz181JNrTjWRLKIQUtOungp5fQAh8D0AiGsuQtG
5p6AWjiXgHjENNluOvYt7vuGsIMNWBme0DzwTRgO3OqRavX8nTcO0xvl7DgCVgUc
SZBIRqBCOcYmP0qbYFrbyNo0ot+zGoZ1szCf3GqMCgf3JrMEcHJmcGkioydvJX/v
wDwSnwTolW9MIWkjsfSxnQprCYlxFv8H6Pdygoc1TuTUz8RyXzmPy+I8nEfpsOSR
shb1WAqqtkfXht1MSIlid2A9W89Zdk/yswXz6S5dEZbrq3vgTYT2d4am3w5yId7x
kXuCnZP2ZURh2iqMhixt0AkWXB0fVaGDF38E8yXQ+X5Oi8DAMzfqW+mP+yRq8oec
2EDbsM31Q96AEDxS2qkm5GDBWg+rGHtV1s4JQouO5fJXAeFBHowZgllCeIsCfhqX
Iql+XZodLKYZeR1jWISO0BBsesjHg8DQqIBCxcAyw8LrPclerB788+dPMtImdr3J
yldX9hQPqtv+opXUIAoFXIBY9GRbnE4DHKfBDQ+Ks7B+WH1WGLxOuCP2nhPfrH9f
pjlIAjux5QXsV0wd1wHtqyUkxj24NBXLpLyUSrcm2FVKpbqzgGXGZbotMNrartzJ
/tYsxtKxJ7laeyXkci+yanGaovHPiTWlUoiaxVu5l/xujHCxEpFQMCeNxy6rOFRf
UM52ammBSaKG5BbGpxCbDlXA2J067mv6jNu776l+UAvdkIm/BtwX+6BEvoY6Z7P5
S6AaAo7rsPjuqP5efEsv1XEQv5YKxdvPzr5CovvfyhAEnlJYjyMJD8Wy+WJOS55a
0RwJvpRNx2vq3FRp6euCZI+EVrTGjyiWDufnEffFbT9vUkYaPCX8kEu3OIIwRYyg
Gc54rZMcAQzkwTaD78WcZGuzscfbFoHVtxQt9ecFqfEoRX8TZjBktdMp/Bm6+d7u
Ma33FjcNzQRAClMKO2TOCqTFjMF7IzBZ+9Igjw9QAECbNtb1sog/+9lKsywplLrX
w87yE1I2JRn7RM2qTCL4AwAQxy+vZxxDKQoMW8skAWreLDlAfsABTtUY6CCp60//
1EMRjjkNAYxPgHP/YkoFIHzTBgxMULoCrNRp4CEWUMHRcVQ7ZmAb72kg5Irr8Dp4
ZbIdtmAuZFAixfHlfJ+DKJhy91VmpXRrV/2w74b5T1+pD8sMfUhac+Qze+6NShhL
UAliAXPjqDdhk+Wn49o3VEWlZM6flQ+AflOTjVwsFUDEaebH2wGlhDZvhuXHgKS0
bSUND9SCmyCbvBtbsg61AOAJBhf+OLqrDAKXrxvm5LZbnV0QxdIDO+IsX9S6m3ul
39RX2lgdy+7hXOTjTgeV89NauT1haM0P9EoUUHI99CBTy3kmFhvAvGRBf35Lzz8m
0fVODUjQ5YTLwMMoQ625Nqmy6gIKhrIfV76J9xcUtOK97Tu7IGVvOD5thO2oOpPh
8r6XAgNjGSdjZYG2tHz+3Z+KxMfTNf6qeWl9mcp8MPyX+AKHQzFi85KTXfDjcxLA
numJJv/1ndBW+uAYcNkvycF6FsbILymHwaCDQKZaNfq7MH02eGygpiuTDIYKPnoO
JOR4hrpwFs/m7fJVcbHDSwCbtkVNFzk6IyaUOY7SHvU/LYTqFin9zoTp16mTrxq2
jRDGWaK4yEviInwUuxeVqorM/IoyS7LqrFvyt+vweu0qDyOJz1qQ4FtUyhAqQCnp
Z5XFDinQc++grA1zVY9+6wfRyUL1Ginx7Fzwbcb52OLD49iw6+ltCAbr9Okk21dL
SG8uY5DjqFWRvNpzR7vovwYeAyL5dRH4szXRRu7SykrMjEIaC4E6b81hHg05O6C4
7z71R59e4ERJFw4wHQBU5eNmq/633w+8oDeR/JG9MBPPGl5vhCSO+yI7RNgNHxXD
k+eWq1yLSQBQ2+eBAJ2ewz7K2rvci5+kv7AcN8fAfEm9RBeJCw4fK9phiFr3uDTL
Fv90NeSWy9898BisHEFK2wQhxUa3UtOMTCtehdGJCivP+A/D8oXpefdKozbh/vPW
V1lih9fWPT16WA6huOXvLzRtYDTpl4VWm3Hs1wN9M179DP6WrFSFx40J+YX7Vh7L
OWgXIUmiC+00PqGsCJEYzW2bMDVFifm7Y3T39idmukzOoNJq0R9rxwlXZvLm9Ep/
I9LGE7AB++ofyRMJc5rH8OF7SNvVWjKrDPLgICu28d4KZtkLo9VcCgtKoBlXi+9z
9YBeH4b0uqJKN+99MQdC9cx4HdLhBfN9FH/ngzw4hS13xhxazDp11iM1AGLZmff0
ebeZi+TaYNQANThT0S7puogyWM5M7cPE5L+uceBjOB7JstB9/5/NlAFHjM0Vbeok
kibcGNsANTc7M7q5Tc79BnEDRgEAJHeYCo7tbg2SXRZhu94cOKApuNIghgUmLYSw
tFc/SjTLMZoFZ7FJVSAVIr65JCY+A2fg8rtfYWXVFM4fjQlFCfbWR08DSEUNg5Fe
uF5jaih5O2ZBiHia92NXDQKBlcZtDiSXOQscyzDApyWyUJE/ehMUzvZUti4N/QrK
0LhfmOHLLBXhnhaU6oQPVIAwXKwZkFFlVpGcFHUwjiy6XVRnIRAWx7vzij5hN77i
Biag9lDZuoCztPoCYUSyKJIgfi4VoIFbn8wpZynEsoVqPTFvkABcxSz09B2ah88n
2hMUhauxApXQMNLwFCmKsn1olBc1KtjIuueYvLqUtm0+K1/OBBg9oBfzc9hAV2Nw
CpJCbUTgdT9VyiHsi/QuJX8zq+QMr+f+LDs/wW9eDwhzD0r6mI02ADP4T+9QD+7Y
upPEomoWHcoTSXUfTEcNF+9AW1PgpXZnVIRBerxRpPxDwWFjtgatyZ3iv18a8iDr
s8d9PzXMvUBxvBiIrclICJ88qeM4muxN3xn6gaTJnyJL8BiTGHUpYoDqCUDT9+D5
zNKJ+QqAonavQbi/x1b5W7lqtfgnbVnx4ElkogJkb00y9bVD438IVhXiQyoFhQ+5
A1qMF6DRd9u0Jc5kRudMv2plVNZ9WdMtcUtzfPPlJCMqvn9FNxGXetv/Bz0y5Ov4
lAvegSvri4mEAJ6HvhsSoCAka2yNTnH3NauyBpSDNYCZPFZsGZMM4u4TsbYwdMEo
6b1vUVqxABU2TTZz9p/NQyc0StilkMAXQq/QnAMAlMZlWGQhLCLVqnqgQHhFvvCW
MN0mkZYgksO9mLUDOFtMheFSIoGqGsOl2+4CUBwhmJsMsiZy/mZAgBjZUAh53I/4
IDrWwi79SV2vGM0JQaVx9ec5H4Dl7J5DLRwaaUdbKIXZDMVzoqUexAvYNZ+FGkRJ
zasGDgDnOMLjZWjEYnF8/WCTp4nldeEJAEEhb5UGHgehUUvb3Fen61Qj9/DptCKD
jr47URoKEw4hMQfblL0GDy3sW0EPwl1+oGunMoUoeEqekLKsoG44DF0srVq8nqGz
P6gmvv2XQRm2+vyz5wrYZZ09roZuYc+MWCbK/8Tji/6pRFzykB06SBMOJlFUy3nd
taWnno8ov1935Mu5Ba1PmJ14yWXKw01wxtVjRG6csQ4y2mJSGzuLMRiLCSnqv1j3
7iVIUEGT8wQhJ7dJpyFAJz8eabLWPOkqeF6G94Mce3abYs3W1xXiPYJigEcB19I9
YqH98PltfhK1BOQB3SSe+SvEjrzaXprYJN7WTm1pdruJCT5RaIlT/38t6LHHnbSY
l3YTXL4W9Qf5ZXJr6v0uo1SVXFjqcuF7r853pnc8k7au2RFvrp2WXFKv7ugcxWtl
UgUgRxnTvPxBhS2urlm93BbgymZy1hRItfITAViFhJpq2vMN0lCbIBC82e0NJgm9
PvjmkjlLiwO0Z9EZ4lZy0zQrPDjfzqc1+hG3qW7yG417cQf4cyAb9KI5U7HohaLa
E86TxVIvyhibf1ZtZEPj2EoWc2kxIWSTXW4zH4djyLe9ZogaKjrxijsRim6SApEN
Wfuj3yKFGDRO8PhLyRN3XR8ReKhXa23TSSxD4BTLhL2T2T1ftjZ11qCWpLIrK1ln
dAmh1BWThIlui1KDsrONm5dr1fjHVKm5m9ikJqa+FzZIwqRb5hGmk2wZZahdXNSP
fOrnUUIz/wZiG6pvq5KpsEDqXWzIZP8x1NV1625hkpI3HnxLYxXFI5PJ8+QfFcVF
PYmBRZWZFeLhc5MDUehdot/OW7xJQ1/TyMfp4Kd25wxiH+ip2JdbbCrOxKATB6Sc
5040dEufQkSJPsIB2oLEvmn8Yy2YrexA+1joBLitvHJImPUQ1bzy3ZLsI27VvpSg
6ZBCie83oYcNa2vC06u5HAPu8DrHAmELkG/IEGVui5NN70wu+QKfIHaXLyhZx0KP
BveuOK3QpnUhnWI/oS7MO+herupxI4OJ5NCEEeGVzTyt3NJ4izkDTh89GWiPAl0J
h3uLutmEK26I8CqOmXcdMlymkK6ThLKk+EnnFn1oou6/vZjn6H7JmSDOeRoAdmfZ
tdNLiz6SmrJsVPhAB2E+rWrKJUaAXieGb2ug4PlziD0E1TMDHSydLG8tfXIo8o3L
FSwpf03iwuXuqtpoApBaHE2WHyWANTZiP/3uxTFZnb83DORgjhyPMOuqd9QLVioL
1aq1gJI/FVsfBjLVXnt851Ry3zsfMg06n4UUO1IPFRd9OXrEUKOpaYFclOsjSpDP
SGUVb3rjtVenYVj0aop11pXK8YP+N88hqSUT4bqSxj5H2vdqx56sbBkeuC9XuU2I
58BBMPCxVitV7K3JLBQGz7dA1pf7TkM/akwjdKvZToLcDS81OFXULSBp/xe3K4HM
qQkIwrTwKRlkTxRDARJ3tblQSivDuSN2aLI9pLmhL54GvGBPEKKChbGllKYCW1SJ
jiBWRH6p+1f1W4gJGVMUnPvEEl5v6Kdbv6YZqVQcUX6bZjgsEu8RtiwZDsN14EZd
OwYmK0dRavny59zKc8pEqIGw3wpNY3xwy2CrCbUf3ROHFcLt6/USqgeOrkbRsj+u
gMmnsnqEK+CIJDf3O2Veyg3yfYBCeuhxWFG2kH98e5SV0yrCuaBvCNN6UgpMAAas
C2/j/XJiP6Dp+lB6tJwDTKOHMNbclag12kR3KKU++5WbN+/KBpJZ/7kr7v5dJmSu
wiqbZ3cwFiNqLqR51Og1xqFaCfTm7O6WAZwokIA+whwQ+J/SeB2t+J6ZIbi3OwVF
wadG6gBs6B2TkNBMnHpf8RgD3xP2Xzfge6vea7zAlVoFmtuqC4EZbWvYkMGI1SPA
HkP8RzLK+LfAWKgIJ1JWHSuzP9+h+UoKj0C6Ok/gVzCUdamz9DeiwZYupVZxVlsF
PhjrRosiB+rOW0Q7gMKlxTKGBdvs6TPvDq5wZtGxe1JlUuCm0zLQafib4JffGcp/
NjbLkJZAYNqAXMydzG7nS1u0vcI2glW+thLgZEZZw4uoRcEO8SkwGamwOUn2V+Dn
6kct8iNa7/f8RlxJLi7sE1F8wzdNOPkiHZmnCQMj8h5IcnSyerzQ14xOwiUvbzR0
E6CjrBh2bPcSGE28prwz4uHIJ9t4c5b0pqfW39IT643dCNKVdjpkDbQPttIvR8Tg
lHw1/XPKFP2frT3MDWA6M3gSmNgNMmUTLK8bcT2IUL1MnjHKbHokt3YIF7hycZ09
YZ4m2+0Rg4zkmyPT5v7XoY3Yb+kag/kpGsN+spyqkRkJkoE0zNsGM3h7uvvLsUzL
TNtaeXVdcLvK2rcNbdmNkiOfWMR7vGzVAoQqoluIkz6P4044tlFBoH5W0YgnVVac
S4CDhuFR41Z5cAvbCUiYyU9n3rzAAqPmLcgv2tu0z8LR5dQE63QL3CtVkXRX5Fi7
snSjBKTv3i0+8koFpB4ZW+RNr6rpIRmKnLzJxPMekq1GA89GdQ+4Gg8EFwuduOzQ
gUr2lEjJQwF1xelNpL2Yc7SAYMMOZbciZMx0ei/TS9Fs7HMbK+v8kY4m2Y4fcOnf
3DdQKMeiQkp2PZEtEysdPjJ7P2Zzsqn/rvOVgwcyU/GuUN0uWAJhFOkvUfL/Sj/Y
lkeVQCkN16caQnpUL/bTfGlqxRA1j6w6J2rCCzAqfW6BPOFDVYBq39BMuLSMz8x1
jlM/nD1chxuqiyN9piZta4QYVIYxuZvya70MO5LGI2Dy2+WVXuvmNtNs8Yq9cVWW
Tz64EBuqYGuwuuT6jKRLwgDlp0Yd1jasX2gy4rpivRH+AFWnJKM4U3ptmJLsJyRH
wY5qfqfbYfC2ceo+5PJ/lSxnRtGu1oK6r9RABG4yU/HOgUHE9NnRhzGdhxtSUxdo
69L3zF7iEbL4jL0LB3jPgZC6h+xWsYoK95Zrd0Q1oCQ08YbFT1iZlhnahms56DdT
EXSuKCw2QFVyBRZ2F1SuaBYFhPGzSPF0GZbkFcFMM5VVAesU4GRNCv2Z+hgIvKga
vCqPklqLXA3pNqMzqhX3pDhv2Es9JaPz3Tfq1qy24O+SuguawBio0eRl1mqA71d+
MFvVXQWR+XstYWI+5CaZV0C0YaE2U3bdcTZuQHxnJkmGHCexfl9b9fwahwH+NJOR
U8LLRBMIMakXd1IMbbG0eLTWOgqRza9X1fjx9178w846Ag64iM/+pjISlPR/V/zb
Xo5dTiJAE8xpWiyKMGBlYVDBp+3XXs++WhvlSvzndF6cdOs7uUaIDDCw7YQMT+UU
DJkFcdfE8acN8NYoGCSSV6rl3DaZpTfQhyRNC4Szfjnzje/yjx6PwUTpSYv/t82J
geEQNPiUiolkdOWKGZ/TkwAQgZfabWIEq4KRibPwnExxLetTeNH+KEZ2m0EbFzbq
iRYzIiCoyx8lNrB3Lbe8TqLI4284gIG/2pRIcnM8ROHOqrxWSezYq6hw88HtILSU
nWrzdUtsDxhUKcxo10YtO7uABqBkHIu06tKKVde+Al8RvNaHAw4ou6YAxsNXA0i6
z7x9MPOG+2OhFEuDd3cGQ9/Rx2oBTjb+Xl4JfXqfIE/ZudgXdYoV2xL1pQX9mQOl
AuEFGWU/0xjg9xFOYF/EDQlbVpKjqVt2awBYn4ILWMzCjiLLRdD/aWTkf0izMY78
t41hMSldEQaGCgNSLGjzdwIrsFF+4x5T/KLousAgRhsN/eGCfnNtfZ0Wt0FZCLEQ
6HHSSEZcy+mf42c0F53RBcfDEp9T3JiUJIEv/kz98qvd1kBtsDdjU23V7r+xD0Xl
9T/xY0P6lIJQx0Wjs+mdBUFmPktRPr3mVnIo4hg3BTEJWQ19lCYmbqKWUEHwzRPm
wsh7IIbOm1plWwvzeO3GCAhXU6GQeawhyubD9aeYyL5RV9gt+nAQEC0RAs7B6gQ2
i/KvUvQPiYyB7ZER/ii/yK68t7hcg4cBQ/R0omZ5V2Fxpnyj5qlSBSfbCpTJLfZM
zx0Kolv7EWpX1DZdNG4UaJoK90bCklJfFP77rgrNFcNMppzcsvWHWWLxzLFhwKKc
UsdIOr83GZyqgD9sYVvifyftX9l/pNjUHjxHekdS4v0JYLnHc3s2fGcEKEUjg6Nt
YLRs3jQMbqICHgSN/qWVnBLirm61V0fiBUGk2hbDDXQIXZ27SYjg6iOm441yWOMG
+zqgx+ALIVKVFgc0STwR6TNnC/cOXcpPSmgOKj4J5bX0Bkp/TtFUKaaSjXa/R0br
RadCP4orhFQ6AIevTtS93pJ6vdgiezLl2W6MW5WXWHS8ceYqMjcNg6dI/22CQAAo
NX9uMEZLTlFdfXQTfUdUFUajFMeTR8RtIQThh1oqDHUeVJj+0/YVTXHfloA0XS6A
bVvZT+/r/t+Lo/0OldW7AxrYMk3JH4Z0RyMVWFp9+XdqGFlRIx8IlHVvRstjkdBz
QSkE2YMVij82N+CxqdnNaJjMkOkYr4Ju6kCg4pQgnVFB44APtGqiHN6UGXHB3Q/n
aUMmBkayTNbiNHGZHYJnh4jxbfk0iYIg0yLVwtH3bm52ZGW4siJm4Kn7JS5z5EeW
eWfIFFISvgG91g4kWFQ41VGB3cm29olzMDh6odtPiEdVM4sp1PThOnEEm7h5m7+M
BTQeyEDBEksTbjIUSPXaLweEW+cmzk1XIQIWMbzei4Boqn6lArI/fYCfW1vE2rAI
EDXB+2D5BY2b/FB0AUhkJTDSh0H9ubMRmaRzlAmNdeyZdcpvnCzhvOEPmCTjsUmQ
VeriKubyLzB6NEFQ6iX+5dSn/GQEd1wWBHg4uVZhaPHD80OvIiw8Z6Rn9Cubbc3U
GIqLE5Nrau6sIcTC5IBbXHW/P6GqNFBa74pzGenKqdedXyW1DKVwH4+JzmmIwjWV
cV2qzAPD/7mCi9lxNrhCB6dWK5wiJAXnWGieZtjeCQ6eCKWqAD04ki8ENj5khvaW
FR3oQmfziVN4sbm49+e91EkRjmoXuy+dOwYxCnq7RPt1yNvOrlCERfs7ICZgGcyV
SmUhzInx9PujqMVGTa86exn3wklLnjifQx8INpIFhHk9JWut0Gxsinn7sTQHZSnx
iQOviDLGNHt8VjtglcfXJ46jIKnopcBYFadNKk2jH/L8CTjN383reQL51dbHITUb
z93BUhNnjLUYbtet7x1xw0ycxS3C5k2/iiBHZ8Pf+tAQT/DhS2WQPR6dqiwxQcO+
cXexrB5OsDHqP4d+NQ8O6Bf09rXbATOIFYTh6CwGs+SbMy6Y5cqYGwnBDRpWK3oP
KnnJvpYJubW7g6FAi+dErhAr7WdIL1K1f4LCxIHM+oD6/gWRIhAkwCdr15KOAEFH
UEL6hjh5xfWCTAt+Fb/NjuBozZ5rmHLiW/CjNGt3IdpgdnAbL3FlpVqDf3upLDv0
z1V9UYc5w+vcS4iQaEvbC78kembMId7mZ0uVtDA0SPZoP4XAq7ekl+l2BFYSSN5W
kcVDpu27etPWYC3Fj+sp7dIeYFb/4Tg4Sfc2lzh0MuRCM7LplplzNKwA/y9eyRXF
mHJ74II4ju3t8c71MN0qhe+/LhkpBmmk0qR1mkx4yY9/FCit4ockEZkwxRm74JF3
huUqMRHwJWUJYy/rkGPzwJorU3eU/ezpiHUyxk+irenEmjq7cZ97z123eoLzZrS/
7m2EjWkt7jNoVqwX0UIhtUbdv1JxxB6mHcB1auOVgfjxNDZlhkCTD3wNV5+VBRSz
7wl98yvuWy2wLxSME8L4VqVG4iAxhP92BX/12CIhAThtzv/BVgiJh+dfseczi2rL
JSuzKKOFnEO6mZsDtluYr+1cDah8+6KgyF1WKD05BW4iA25pAeo2joyBESAlBT8i
v3Cb3lZwRPloQIc9dYWx45Lo4DuAB23iGIugLsp0MwkfsFdDrbd3kX0xBXVh/a02
yx3aFUbSsAYXQ823iGSWgXbnuZPtNgVotjH33hPCzXmiy9AeJSOmxlspUyjeJpl5
71LXWLiMeUuXSpEcsLbjl26VQGTUQ5DOPYixYqQoWb578aKJKVkMdeZ2Xd+s7J8D
QMhQdMKT4AE4zBwE/VDBCcj7nQPtsonIkD2Zm47oehP0C4fKhhT3wmZz9kMy37Xa
DzN4o8njyhXUje3n16QJztqNw8MIuCZDPifxoEIvK08z/StmJCdOChQk1pvpN9lT
lR8gKq7NEziqVlux4UBTVL/hvEE+Tgw4ITXSQmGezNFdKazGu/DBkde/dLw3e9cm
XZaeYmGJZb5Uj3Re98/aZTgrzSYpHicB+/Nt3itU4u8TOicEfdvR0jEHWD2Ni5T8
Y8/vk9MUE2JUx9Y3VCQ8rGrJ6eOhVwEWlCrNDXBeq5mahd78RC+ywcE/jMck++uI
/lpZuMmuy0q15MrSL6GxrBRIA/RU6wETcgww5g86FDdQ6hUwPo0Xf9n6v8a/0RdD
k/SyHYKW8+GNNJ1u+DLGnay+t6Xvnv0Xjc0+HaJ+101hQGdmDEBTMk95/m30eoXi
EN0FOZT+7sdRZVKxo3vPbwePko8KxrFbSzE+4eUwZduVKxwETwrDAw0klsQ4IIbf
ZZNtGpuXh+gyOGO6MnOqJbAJa4hodMmHNSPOOT5ySYN7pGTzDaY4C6R3OhF/GwEa
mW7wZAyNzh0m36XJTwutulZpdxzZiEW4mZgmwacnCy6ANlh7UpYdsI8Kx38RXvFp
aeS3TiLFOMSzmVWorT4/A34LBJbuYeeloUMBFHStdhthIkfmA8OcJmZhcOXy+spe
t2+7MLgRQlxD3Am3icxu5FLHgfLr0F/JOpEZKYmZez6dVkClfzyiUH2Palx5VbIn
KmaqrL7TlLQ8rmLXDclBWQYrUJvsqL8H4F0wKeYdz67PVtdw+fWCE/7tK163+MeO
6aYKcEdDijAfKneZRsURcgMGEMSAC+lIknI2wjyD7FaSkrmUmYN7Y44vSN5LiGHR
7LYsz25bT68+S4p64OpqxYS30XL27l2xmcYxXMpt56q3cZjogzkK9unGhlHRyqDA
d7cbye9egorqBg6AsaM8y/bPaZspYeIa1Nxee+FbDItlky2MtEKsuDwguogv2HUM
3LhXnwsc/+5QuX1P2xrvxbhmhbXhI59n6fLuWyr6snsdZejJr/fhVbvRx31jtjBO
W7KVmgUx3pwNfdvQWmlT2nWZPCNNasD4RV9Zy7T4w+HuoMqf8wi7Ywb4h+hSXgXL
+7hYgsF130zcpm6ISIuKUSyVmjjhTZyqP7k9dPL5EENr+LlxCH/YShYDpyJi3j7L
BvdXXEVole+4YKxcB4hDiKMf5XKWaqukx4SNe+nIwQGUeyGLp/NCptAjqRk5XvKq
AI0ldGzUe04V+fkG2d07J5gHgti4i+QOuCU3vm8swgdm7hl98oEG+oaIXUvNhyJz
7sOy7j4C5whNUOK0xdcehJ22rp9w7OEmjl1JRExd2tJr/9fDNGHICnLGTJeDcgqm
6ccOjWx6SWCWK55FQmm5yCojKwwTJE6HzMEhoCrY6gQZQtUhQr1Ed1bZQGp+RwyC
2HKAr4l9vXybUnVUofh5h3ImeGEO8aWECzH7WvW7VG2s2CbLFzip5Q6u20EGF7Pm
Ar6Cr+vPF5iSlOqWEnarZqMDzFfCHe1fUg6C5NIxEKWwMejoUDcYrSzbujBC2gMJ
Dc1FPjdW4HRVA+RrDBxVbidCdj3NlOgSHjjS/LnOWgxieltWHYhbmgNDIuTxvzTp
jnItaN7fVK4V+eKFvrnQKYgicsJUSENrfjENFCtZ+LoD9POrx1Qovh6Fs0TZ+ZUH
gGL2bdZwUZnrGJ9GVpYqoZaGdNx5qshCBrvCbbhUuWHyp17hj4iiBOvKdxLduMC/
ysNMii3dAUZlQIo0rNvIi57IQ0cevEG9yrNdKDLOBTN7fIPwuCufv7DlRPk51kX6
KBGwWHfQgOMFL1GQl8F0PTpgmK0emRPgqMqQkLbRFEjLfxK6IrqSVGY9/jSSZ35m
U47ejQLbVC0eCcz0K2pgntwslDstYQ0T4Xrxj9nl7qjuwHckvGE5RX2dEI4XrBo8
CHMX4ydxItNjFux9EVi04dZ8ec85s2YV4hXlUy9bxPRXL72/+9R4DJkA0ejtIHxy
GXTHsfCOlj89Jp6U507l/F9kWA9SFs7YpctQnL73FpduiJQmfLlF0pvFbLlpgAiX
9TeMesfK9megKsoLBlIH+7rGFe0wD+iUJvYT1rLaA7CDoC2Ak7jm5WIdsTkPpV4I
3JHZe5h5ybv1Ty9Ny+QC2fnoZMA6jThPpap1cFvoqKaQULLZP/X6wloHmPwsRsev
Ze2C125mipeM8lRSF023Oq35g9+9e8wtedHWpHr3m1ekL1n1MrVxweAjVuQEMzCB
7DZHyxQ2ltAmejqWA53lypQN1PTmW3gKwwZgf7jTvwsVA/3JPnlmOGLSowbf3jb2
7yrOvAa7xp/48pa3zhHoBddDQy7IW0j5SQRuv/RdAoAbQWpHxJYdpkcFFGmCcP/r
z7s4xzTIsamxjgfXgT1r2o7Kj5wZe4UmJCccsExU3wxJ36x9cgDohk0hZKvltX9b
ePhDFusZc+YB8aYzMfo+yADa3cG+v+DYBtvfwRiJmfnJBeYI4R2xEa0qIghHDyXr
qe7yJxNmLlp/hOu5Lak0DzSTKsIkPBI06+uPe71CBdbbHsxqe2Sg4xByDq89iK0E
qBxPJoZUgCw5DffmhT8anGMDMSy2zfZ1oDtpJt2f0rLqcSdkMs86/YcQnAtcm4eB
1VK8W95HJLBQ4u8frWSSYGKgv21ITBdMvR/5uflB2qJSEan/2YuENB0O3WA08R9N
fAJr13MUY+bclpEXKr/hw1CwRfcFJNEBNQ9p4VZEOzMAcOFVGWwZy71201ay+9bZ
Sg0yFgWQwlF9sgHLV4UrbtKjDs9eznOQiKwr3OqRlr4RhB8gvGu4nCPGtQTV97It
xAnXnCpbpq+n9kxfJFMroGciM65od3HTKJEwJvHluOJSHnBBl358XXDebmoMagbS
51Zj2J4lc3kg/5ux89H69lL4WREscpS7qZcGqPSznoID/azn1B0nGM2af7Nyp8JA
ia3Qc+nm2ho4fMeyU8ehIo3idkNNjkWrWH4wFKVkWb9Q4oUQ6B3cRiQvq1c2YXb6
FabqwSa6+DVzT480zXIeLrJ53j7LPl1i8yGiRVmf2YZKemu71t2xpC35+J5xpqxz
csO82ry9MyvCzbp/NWD7Z+c27oud+Ldl6Zti+BCQiRW6A/YXiL9FPvR18YJltTEY
QFrzsPBcSgppS5TrSK4SakHuGa3R9yyGnb2nnBhABJ+d2LZH/v9U4HMRdVCWI6bM
DX+1m+vzpwX2K3coNSLgG0uJBewuowagvke0x27RaA26fNVxU+aCd7q9T4JFgkCo
AIbhc90Hnie1yRX1IqWbbV2HRgszgVPB9qsroknBubYJcwyj1IPQUidEEGgHMoZx
MUA703tN97WcMXZh5Xq50nkAvRE14qCPF58dizv/EwnMIfLOnU9a2EQQgC1IbeYI
QyJwQQgSaXk8HbYYPnx4LMh8r1A2IoXWEhyRWND9D/+ySBrb2TCM9NLtImW1p2E9
U2xkiOEkYNhB4sw1RF+NYGWqggKDu7QdFiLkXYgKirxlYZT7JWCBCCZTIPIaowL7
puj4F0165iL8EjnHrN0Q7/gBzYGadnGp8dsobkvH/IzrlaSc0pQt7l3OXIgfIzxj
OBX03A6svzJytmz8Et0+K7H47soJZmIM+3SHTZfWqpsTeEdd2vl+R99ZCJVo0oR3
XdrnIUg76qQfVY3N2EwZUYgu8b1tGjhzUfLcvW9AJgv3tEiJ8gvEDBGv1wA7LmrM
ezYfWOUFItGFDn39MpBYM668dl9Y6YCOHz/V6b363+h5Fp/2rxnq2VjxXkfFbapT
MrRYMzGyeAnfbuqQ+RCAuE2iBqaeJty9UohuesRJr4Jm8foRNTbFIBgltXRzubSc
gnL48tUCXQ0OgBXmo00MvFJ8pml6KYpo46Z1tmRHntNCMh2z3yo7RFoAmBlXY0AA
ub/DZA0FVBaFrb2XeWgAEbcjZ/rKWjUFG1cosZEMckeZVlyijksKxw9oS/Zn/tmT
hZK4UA1qrT8eR5SFUXhgNM14hGvH39DYc+AeUxlzP3vbFW/lOsDsF8WnXQ4QdyGF
4yrY/pXF6yGL0SKm6q7q9NJ5GnkTTV9/XWln8cclqEHL4gCipUw/hkmUExK422tx
VcvwUCzu5hxL41DL38eExR723Qa+HsVvd0hcKM0u1s/H/c5fJrxOAikXeX6MYDj7
riZeKMGygKf8YomUDfXhDhHqcFNMrkrHo3AONdIX3Gzjw4J3Z4RxiEeVcJgzTctH
AOk2jZ2ChWKXIaIOkGE7C7xiSh5pNenQ3GoYOew2T/xcirrHotNxs0MA9e6PdBXb
9aqJlBIYgJWvLzyjEM5zQbRLZ4wu7vAPMtfc7PDrc9C+5eleAL6lwywNaItWCx11
U/Z7T6XxA+rhSt2tYyZXSUl1yfCbq1sGTuI4R6mR2Kf+3P5r/axmQmfeiK1ap4fl
UkgqYOhpvaRxU+eHeiIss4l5vCVvrNgqlttBknxKTtHfQdYoitZEAfoL4eQc46UF
K/a+ish9/PGULJJ69NaHnehXEtaKY9/HTsA3Wofs5MXJMYUkfW4D8CLykzQpliM2
AAYF/Pl1kgtWoVBpBrv08qWnSRlIhdqM5jBrvFIlNuQ9WOpP1W7lc6o8vqjczYZ0
gAQkrOyfeiO5c3t5aDQlTal25ktzVgrHiG/ofvVK/js4wbWbW8/Vk1MpckX+TV5R
Cq+TAB8BXjsTn1CmVqNBxVGeokSNVMG/8J0Eyz0OCq1qMfKINvV7a469lkqOL9ef
T1Ysz5xdUa/lhuY2dUk0vnw87PDEsSSVmtro6YL8XQUexP6UBEAXPw5J/KXaDelF
e1pCYBLZRNwDUrxXIAAQQXC6S0mGQbzPOpaei+orPrb7wRNZmh0E8VnscaoQvdKL
mEGNV92OGhobi6YZZUn3wIwyIgtDKWplfPnRn9KsMqunNqRnWjCBAoU2i5P5s7Ct
btNlgU/z4+BBuArO00uokDzY0YEPtmFIDSvDpCUnCtCk70gWMHAHFq37zvlvCUNy
lurVP2xDjRjrnW2AHXa9oPsONpd+fpb8QPpLFy7uCq5ksgy/d+hVHoPwFGcKAHZK
x1KQ1SnPx1BRrYt8mUxqlTByi+1d/hFRRgKisCtmMDM1fa8SIvpZokdFS0S9V/jX
Bo4v9gEHSlVVoZ8UbE2AYWzjY9XfrofK3lpNh4qWbEzT1zFMQUhFw4xXA4Cdxio6
MeLf5u1Oyh0rcI98bfscw074Qr1XRBWsjl+DEvuSuPWmqNa8GXlO8KcKmCTTFp9x
p4s6MiDt5ObqMWU4/Iuqm0/mH0uGTYs5TVV8w6Jf8X/00tSEpSfqdxrIWMiQzaT5
w33Hly78+q3DE99qJhTIIdpTG2kC/ZIvKkQrO3IZMJOqEjWTgv1sbTy0HGQnYne4
iC8KEv0XhzMMkbdoLe5SPPxmM4rncv5eTbR9vK+WLa7o6cC7b0HGm6uuM5heeLUs
v9mpYM/6jMcl6wXrZEmghiZW/aJ+R0Bp6ju629AkuU65ODPd3Cp3WAMzWa0n396f
Sd9HTnYMdnrWyn0roaEqTCnh1g9y1VV+VWuxdP5E45gXVKYtoJrYFhXy+Anrgsuw
kYPRGbDgC8SENIn/pDnVJdXEIL4P3pJ4icG2tUVEfrgAHuaXgT6ri+4uFM4t0xpS
jOUmtzkiD1qclK+OkfZA1CDlX+bj4178pQ1EAqeS4OJnT/kw8qw51WeqQ+a1MsY3
9RzBjCmfm1QR5rRkVIB7A8GSom+S4Gc2YlN82xiOooPBzFWXFWqoReG/q0iMEF7o
c1ScU72wLc/KW0+qkRtJbhgbo9lfrJ8IPDFFdZNZCFkgB8C4Z9GmHw6jRyZ871sQ
gcrwzL0bCBsXirSxSK05WFu/IL1ZW/rK2bLecvuG+eGB1ic+KmPQ0CALW1BOF8ki
bw9yjcruVH1IpE6xypL/jRJW8T9Wp9tZvYvu/Kju3Lvmpsh1HalURfM3sQDu8dMa
plBbp1zqT+zYpwKOnGKgdVf6wbX1HQpSSX5/E6EJ5Df1HZKqgDRcSu/KsdC3vvZq
EdviLgwsHTMD9lml9fH/ULz/z2abx2XuymcJyhNjjEYgkdbSbtbx2XNQFt4Csu2/
+4wCAc2bnLLx/2RTTjZ7tlCFgoFpRjO+UMlayZaNX8toWFEhQTor/G8p/aSTyPL7
w4n2SwMUzGxv665MC1FI3j40ZYfw1MXJzPitCFrzL5nsbfOvQlYgrO3IoSUna2lR
lztIcchzvnZNDvxa11Hiivo3Kl3HNqVbZ8uIWQ+P/xL6CvsD5nhgTvBz2qyWUyUz
czNgZQCcYMA7pL3bqoTB3o5KZrLwExLvEh+hXqENF5OoSX+SSCR49yecUKxRGvd+
qEl3l4/eXCMKaAeVOz9wbd/73VTs/cKVL5sXtohXxnuP1PkdcfD4F9lPUDinHbZm
ssSbreGlOjWVWOkeHSiuyVUnrIHZc5ZajeIKeJ+UT12ezGZHLk4p9ZTa9Ofy1iMw
x61YBiYdUMgGU1k2Ye5qnEYujpBeJVq5kzaB7rqMCGKeL62cAfZICF5GSnZ1QtVt
V6K1ESMU8LCaVz1RBW3WplReYPsOv3N2z0p0Qg26NJj7tdcU7Ek8FJ5yq+jMbUve
7zmQO/nvnzBAtBl0ef9ikhJ9TU9ytMGsK9IvxF+ZeOy8Yz2hCrIom9i5OsO+HXVu
5/P7crFCbzd/fR775EpeqUEEOrZelRqyfzgtLYh9VJQN5vee5oWPCP1j1ySAgu5J
sHwLleTxz4g7pOKa9nWbu6HUQLIzsAtWcaJd3uGNFotrEWuK8VolMHjE0lX3X1PF
gCsijxw63BSKPsKhsTHlOmN7DoIbQFH1u+CctMSJ84Cc70tJDMp1DVdq8y8FapSK
LHW2gMf1VeVaIyoVkvbn1djK8/3Z0fRvTKzW+i5+aQOsUXzgPdQyX9UAAFOe1jB1
1d/PRr4FtR94sJSY8J8fBf3vnZ/p8kPJsHkIchQHsWWf7PFgiHgiyOjf73sWhpsz
MSqgx7fx39V9NcmstUjQTcC02KAjIaHbdpYV+mxZ1gpmdRUyhNJsrTL6vjihLIPd
mvnHovRb8ze97XNx64u0W7q+q5X5poboJFW0ez165H3mi0MwiEFRrqvdkjhK/hU6
ne8SmZXk9aLSPRg+oEi47QXo16EmgL/4q+E0aKSIvJftCI1TSEFsxvnvY785KP0F
RZohS3A5MnhU+ShZtl7Os0+goKqU/+H3502gqLZCiRyLE2QLhfQ3LmQnx6nsvVFo
c0p+28l/IISywLPtpq4V4iny43XBunUmDRwISi3byWv2QmoV8xU1UzL9mIVwSftS
A9cwSW6OZ62v1D/YWWQEa/CJsiHbBBQrYj7UwLuG5B4waCjGmuZduap7aQFbq/uu
gmfjRPils9rRC2qZWG6YCzzW8brnZpRjnxz4ViKLUqpZmmJT/LytyR36TjOz3ZRL
kPFubjl8F1Umcg8K6M9x4iBkt7fYyuabJy01LuJNKUgr69Hxe1CQqA2O2H5w2+40
kUUB572Fn7nCevInTN4UQyNmLpT0fxnL4+VFZWd5FeAzAbgwsS93VGPZRrWHbC4i
NvSUam3zt4sWCbg4PJ8D+/6e0gRFXpe+fjTj9oeh++t4C5tdVSxZar0bkWMFn9a4
2JUu1fNSvNp24E5GRFnvWocDLSCuGA/OlmIGwVrMvTeIyAoyfEDznPf1AURhBAMj
mppoty1sP07G7f4gOtQ1ti9jW5wTmImIPLU2E8pZ8ftFqNCqOFc+eXMq8HceUFzJ
cAglV9UJK6eE6kz0BeceJyXSX0RV8v2poH43DMz69twNiDUhWLPeQBmgo9d2qf2A
RTruHcY+96M1pXzUl1sKJuJ4ncgz/VIE0BYrOrEFv2p2NpV18NPmGtydm8cn1Uky
1mr4b6fL6NahEsft38zYNy79/p/oeRkofoWb/O+hXTt+Ler7eTEl8CUyXXcB/IIo
PiIfxfTKUCxHhBUtBsonXEMa7amDOeX0S+sZ7A5LCVv5kHwhTXbyzVZeryk+J+Ej
zx1z0Zteec/dPzPaMGR9AbtzxT7hwJfFg9hQWEL5duBIpoW8ndcKZ0D/1Tv+qXon
pbhnOT2K3a+4oqfDU5wExYyF7qqTNxVzd/2wIu9brDh0cDwZHXSGH+cglbebjrzK
3d2LMZSIsZlWZi1QY8taAYKEC2Pc+TVpau6odW7rEi1dJer2CpNNn4VKlnx3aGU8
WhbbioSTvu1/Jy7534JqJFajD/xzq4bGXcKp/6pbAMluo/RcWxCJrrO3qj9zJ9vj
RKFltXreAgseI5UIjS8cdtFvTZKoNJfDmzlunREgGxQIGjDNzHer0yW3ZeApXMni
fyTBUVyUBLVKasXxyZoqJCm2ms6Q/ZC4WeAc07ZqNiSP+x9qVaKNk7CnHxYoVZ5G
DJdCozxjGghWJP1UlWoe4lrwlzUcS+P3daRSC1uSBt4jLJyJX4YlaniRmXW641Kv
k3lblMHfQjBn1Kr7v4SvONK7pf+2fwwyOo0MCYNQsNup5KAa1rFNoW4ohwZ8c3wM
bHBkLOhzgRH77v+MeCkK081I5Ur2qC6Kbg/T3nDDWdPltk0KXk0JjJLoowZX0tGf
cMIbqxmUQN917Rzdc2tvXjw//iVI0o53QRJ2DtE2SuRwLZrtT6BczuA1Lz23BZOb
SNqKP1Zn6tAKc56Tfgh1Wj1S5NUNH+DadylBKhPhEqj2qrocDpGo7ZJGqVoyHCIN
C9svk5THLJahLzE+naXhr650yv3SdKMpSPtEdnuGgTTzgZcXyfg0j3y94bSzTvn4
aQ7r+TPTInrNNhoxXSJeZNNDIcs6NW1Oz8OcL7O9nZra60vHS2jS+XQKtlexGuYs
0lQrPio7D5atpJr1UPZWrgnNs/p6ONN5SQl8U8gNvitJRJFSBJtJOZTnny3ksxsl
KhDKaY3+wkZXiWTD+EdGL8FVRBEoXWSajJwfyBaf9pLS79QVRDf+1teAialC2QQ9
3zGYt3mT4qn/9x3nvY10Tc2w33pnAtEPu6xJ6IJ4p81jY5DML+1ScFmBEoaW45b4
pwh2FN5hM/h6jEECOc/+vgNzwIdNOHZMlkgMChxD4XLJ/jPL7xn762uWhD1aSTzN
k8mTbJ3CTGSM+MqDwVsa1oe4nb/9JquUyHjTzWaG2hdJlyxQIrsX0IrPyCChwQMF
HlGvcRY9/vv8TfiaqFgOHEwsj8NDoaoLS0tLEs9XMfoA/Hiy7eIkjekxeuHnWBLM
hMmkbDMQ8CSekWMTVhvrxlvWqlu20D7nIGfOID8KZtLpsCOSAPPJIGi8yPP2WoeH
O2HOsNHNpHhrmlIwoeU858ov01CDfNYLSGmytNc+2iFgNuNUlp3rfDWsbDbzOOYG
maf9HZZ2BaS/WG4Y3GcSALo3pDMxGqtYGjz0O0dlGWqDy/cB2cLsNaC4QOw0ywIk
t5F/C+JPosCaqJaaJmYHjW0tKdrEIzv0FpuajmkzOlBbPEnsttC1lZ5QKdBJjj4T
Y2wOA7E8DJp9amTUNGWBvSEHiJvRxJ1SpLewVVjOgrXOijegwQPS1gii5hsPH3VP
EdUwBgO3Zb2D4IaIOLQ590Zh5E4FR6drWT8t/s3qU1sbqIOGWyzczNRcOZAuuihH
6+za4RX+j9cuWNSTcGlJ4z7gAqSB4xOlido2qaOMU/jfk0qhBsZjvqJIJFvmZrLL
PfeRBqQDxHxxNJkDC4Ocj2DujVWQVhMfqIHvSBv19Vn6OBNRY8rxhFjQbVGPCkDC
3MyK6JILeSnqXxlfhcLh8Xg63ksssHAOSsuBtCjzthQs/JPfG80xPWaOY7rXTmf+
rbxoMW7E3d9sbPNGmLaaSJXeTi2wLr8a3r3rqxM+3HXlL7mX++OwDWEcugiO699S
ja56HzjBPxOCZTX8sYzfo8DN4fR0w7mfR+A+MvR/2RpvO5w2g8HBebv4q2sK1uJr
dAopn1RQr8VXz5Pux0FxnLdWZsK5OMdc18xfqZKHxKgEEe+1s8IR35TKSuNONv7b
Y0CbOpBpCXmkk9Ze9JMpHKb+7CG8G2If/z0eGI6SfhXs9ohaFu8QQkqAPEUjEc2x
l4lIWTWqdfIIojNANmFyVtV9AD1soSR3QOHBXTydTJrUyj0RahMRJan5L+LjZMDw
iKvSoGoMANBZjWHRs7XmstbSZS127hMPVE2AF/48hr5zTHxRCVjmrL4Wd7fIbCeg
g2DXWkidqYhOYzMKPjPdzhZBlX7amvBhRoBv38oMDadWynvLmlrlzjGDiWCuX8hY
56OMS/Y5LscWW5p81rgb5rR3MHBG+SMLkKr3kWsH9qDqcsj2jOPxwIiPYW40WXkA
MK61zubEiCvSjh8EC3LucYRo39Dx/KQa31BXwz9hCu33QR7n73bohkswExaIiisJ
Am86l3BLGoS/j9MEdzvwn5KaA0852J1026ykzt77R0m2OmOm8+hMTdQ9tNUvkNQ5
w11znMRSEFTaUi0KL6rxWfBTjl5P4uZMS2K/QP22uT5OT9FnANwNvXLU9yyNHwEh
XVHY8MkkHhdgaKSKSDt9KnC0/gvqIlt9Q9zIPcmzp1bqjjTGcce3bjxi0QCv4MA3
5c3R+gUaMpPbCUNvAX+xCDx2pUS/yRS6kpJ5JzW8yMpTIzcoG2jSM0tzwdzYQ4KK
3Qra0EhHAB3jLwQYETaqvMU2FyYwby4qlq4X5shcKysZsbptVzHPqPe2CwEjJMDG
ZLVY//tjh/tNpmAM3+YSatBzWqtMAbg690n/J5WQyH+5n5p5bWAvqw8hJBptu+62
w8OEwBldFIbeF0BgXehjjN2PccJNRRYpCKKJbCUnKmRdpvRZtux5VDK9h6RQNnDI
19ngqSoDcQUdyLU42GlDBcGR4FwaNFSM4z8UU9+Yex1LP4JoiaV9uUWu3ZHAsrZS
+c0wJhjmWlkxqIIV0Jq6iJmrw7bG4CYjhdZDE+RBMk7EuesCi+1ilW/TnNL0gBMp
N21dQs2UzxUjWbx57HMCtaA88hYJOla3ueDInCA8XwqIs31VEDUg3F1lLHX8jylK
A6MJbofFYYQx6B1668AKE7T0x6mAJnYrmmY0p0lESryBd3Wj8PG6SpRCZUOpUcM1
ksUs2XJ5c1qsHEeF5J3GA8U278D53G4DfUutoUFbKYSgYw9DYjpobOju4dmTcZ2r
M1K6/Oty8eJXQ7IxbyQwKbkrTnZh7X/w3wiPriabgDdElrssPNf3uOydjD/suYUO
qMAMQpqXjH97nVw4W8RfBvDdbFH9m5/bndiLQ42T3QSSj2Muowrf6Z4gQFMyLy3x
vcVbYZR8r0DCLSAYiCQqUtKdviyRiwjLngUQjujntwuocWwTc7PaYlgvv15OzwTm
qgCEDYS1t20GvWUfXRRmfjcOEypxYPqvYiFIo1Kkubp+I9DLZZDN8O68fif6pRSu
6WLSp8EbZKS1VbXpbUSJk3DYLbzuxOuRkHyOkPlzuolekcz0Io8+2oA+DL5ANUjk
hQ4pkGkBAfLldr53jYPY7ENwngwymV5YL86/wyuWjiYznIz5K5gklAHk7IF7RDYH
mxd4N2Bqm1Vc3VjP2xXw6Zh6bs5uPX6zmdmKllPnQOe3x8THXMamS4I+9p7WIFhs
KiPWxkMHbfhza+owlMaFIYY+Th3Kk1XWThJaw+b5QA9R4jDFkqmXcX55mcYTZ1dT
SSg1ZxugXyqKPQFWzowupb1+0JCzaNOWcICla7RGNsjmT+0llHG+F6SNcBX2K2Hx
P+rpn4a7C+MF423/K9Uyy2TU8jwbIj6V60BtjmU0Pmz2aUt132CDmjALiDX78qx9
jRgE4apXchdWf7Aolr2f5wgvqfgopRx2lieMXiWEHXqzF6P3fvo37fdSvWDb5pB/
u0d87ehLiqMrSk5goKFnl7qac69FPsBdaRSkgFzhGta9oom5ucZgxAU/GfjtRmqc
U01O9Id3noyuFJ0OUQ5XIq8TM9sa/P4Hu5EEDQNXWYRMpXsJ8xO93Aa69cB4i4JN
lwJu9zAhS2bg6/vM7eRGw/KLuiJPUSHrUOsVmd5SN5xj/qnPTSylPxxfoOBVkeoU
OnS8SPCFa20dqOfe6nRknhBciuOYazE4MFzO4ilvN1TCR4K9ZJwRtwBLAACeZrvH
vN8pMOFn8ckNTu7FVgsDnfW+i9eCVKmVk6jpJvPDFyohQ4KygnyxPYMv1OOVV+Nv
Kslrj8B+EHhon89rf2MvIPZISms+AXaojHYvo12Cx8wIDuXJ2Cx5el1y/+kesXYn
UcaLWTgPHbszb780YPVX3EluEet4DPbpHCGHqoB83TftOuOAcYc8QLUbFZaQ22bU
z30E0h3kb7SAMRsOs/e/AuArHgFnQmy6oFDJMe1BVns4BYlNcHFF2cTnB9K+xZi9
asZsFnsG4P6jb7U83OP+Mzx+0sDoj6e1S2fHekYp80wVkaN+bQd4KSzb3G3pC2A5
9UmxonQQ8a+VqW2tgVm+UZ9x8SVw86pd+9yQp1ci5E1zheJ1kzMNUKY0E1XplQUa
xTKGORxdEw1l3SM5ogKskP3PEEbq0Rs+fRt1mKcOEIVgR6ZVbSqT4vwEFSc9KomM
M1ZIy35iZys55Zx73OxBUP9mNyT8TYiN1lFSCpmCu/6eCGnihlYStfn1rsCrhaHa
jpECd8ybs5cCipiq9D+ny1A5f9VZFoaNpJGohb1IxydTW9XP3y0XGFFXkMGhcWce
mj/SEl0Y/s+QhrZOlO+huzw6yxP7AbHonaYuY8lRaeASqMtSGlbuKKzjamfA8y2M
OVx4ChDPzB4JRozVLaR2eqzY1j/uXwCrX0bsr0cqTHKVxsQAd78Lz3yBa++FbM35
RysfJIkB0ETUVHKnMf8ImJymU3sU3ObTtEeCt5snvbdl9r8CU01SIRETqneO2KbB
VP5TGwrB+UM4MGK1ho5mtWFPargoVqPC1fgLxDqASNZ1dg7n0HC2RFeUHGGpXV2/
wIkqrddV6JpSupJc9L+NA8TR43BRMWGtrodwhEV0uZc+APPitM3Nv+DYieCYcxHp
VPtkb9ai0/Jftalt7peuuoeCreJjibppL4CATRNSetWZiQ6R+R26triIFUMvdFQu
/St6SoulPYw23nM95ku31qiQMJjKrsa1GgXlhAATrG1xyn1qtfyVwLKBSnbwJMFm
S2ta4bc5DmE3CxK2qOdMnsgTasoeKIkDv3l6pjs2DWXIcBbSpshUhbaD9pudfQl0
egLV9nDflnonC/6rzm59hal2P6xVRMcIOiiRP5WKjp6TxVMDhJA6HcwdCqs1EOKi
uegRX6J40elVJov+g6z119ZvZ0aIZh9NHetM5MFS8bWRYKkT3zAuqQykzIyVxSMc
jh8scvpX+rpuhKueyJbAizLY4ZM8OT76p9Pw/57VGLWHfatDoZsvwPjjYEc0qyn4
ov2w24gaCsNqmvhwa+E5tVqxv7TqrrJBVoZh+j47kkNPJHAqKYk/luXbxcGbOzy1
JrU9oLd9FvVmzhS2Rh+b4VEiEp8UO5C3rv1YMAH9PyVqas2WLsFvzg15zhrBzHKk
gIBoJcEygIdC1TuHjREbqNJfgZI1rvAh/foUPXZ6U+jUqftKeGi1KFymPfgSTKwV
SNN0WAZcA78GIZ+E5e2UklrI7zS1sq04h+ghBfU43xLiUsFNgc615krawWeoNmCU
i/cnF318h7Eylf3u5eZmzl2b1liG52LIibXCPM3/og6eJjnOs97WC6+W2X/DE/AK
zEdkwDOWbG2MTBkdwgikurghLOFRKYiCtgN6svZj6lFrZ8kyB9X3ZJIseglBsdbT
9G1CVlOnQbqkTa6fjqktkDNzyxT9kPA9UeTEFedpXnvGqlZTtHY1HYiHSJjC/Hom
DEt/fCvCA7BG5CLJCEGR+jLdg1mFmrL/mMWInJ2IJGbEk4LX5oIShm+DcBnMitLv
Afn8BC0foUiaMhSosi2XhPopYlvJ/ua3jHVjoZqM/7LJcP3eOJp/ZP3ClDp7niQA
mP5B8RkV1YHJ8cK1rwdRsaL6Ql2m7u8yZMqjFWjSZmbq3KQFvBNUf39/4XMBllyz
Oyg5aeACuYhK29A9jUKrcHAFyRQjbZ94YlEbRArvahrihn7/HqIUV+m5SSQa8n/3
3F7yIkzX+8ru0KNgVKcI4T8Ib27Ry/Acm9lB3ld3JqsAlmXIKTNs/LxP+dPGtLxn
Bd4SwcVvHk/MPnRpAb/yBm6tr1f3fcV/igWR/8hI749gB4NZjN3aTwqW6M+4WnCm
uOU5EtpT5a48oIgClm7HsZeQ+6YhntCsG4JE32vNsLgXjQVlQ+tQn3m6riEP/Vjt
QSK13XEoEVZS8IXJ92rT/0+nlYu0AqxIbfWVMjX5RapRuxObsxj7gbgVltGcAvTY
J6MoNfjHMjbpWXc/q5jw1rbITsnGxSdkPYC0cCD7Sv9Tzepv0RRtNXxdGf+TvAxW
rd7aslln/5ZQANp3BIaz2fHZ/HAyxjWzhiG7+c9tBHuIkyqBhsaV3wVtkyaPgQkh
Ya6HJXDdwbh1wJ6uMhio8O1d7KjHSSemmq3mTq2677BuQK8RZt1sEY6qjYfKo10X
vHXbw+Qvqqswrw9oUxN50U3Pkmc2NDuJJL8lv5fzdaGE5iMLt52fn/0bQM5j0UgB
Y0WusciqZAHuikSMEDaF+HVVmUdlRPG8v9V0Jt3DuAkslMbW8MpAFKnqUxBcNXXS
OURJOmRbHp4UZZjrkvKXjkL5ZEnYRR97JcEuy/3cgg2Bpqc6Q2J2gNxsWCoiUDub
EoCgnrPct65hRqVZsauaIaDx8tiGYM7yFEKqKLHJH5HnSjKxWXVgZa9FLReeRvq6
NdZFJTs2/aO0KTVj1mhru4017urfkbc9r/US3eiVP3NcrBM/h2Q5ShUpp+2wnaYN
fJg340yAPurt1EacTSAimbN/mD9jGNr7P3nGUUYx0DOdjMixnwG7i563WXcSwjll
cJSH9x5luTt8bxH+StyB5JPxb/Du+QPvT/04ypKdAShLNfvOBJAZRHJL2Yq/jjCQ
kOVU48ZGzCMFbqW6EXtdjifKpB7f++1gs5WTZgEghLehH5sIuHoIENoMYNYD9oEl
/+iDphwTP6v4CQGvLRabODJDtJHpH3OeKH1YSpEc/yMS47gqFfjOiV2QbOz2t8rX
8KCxx+OfJjK9pJU0tZUtmldkfVt/mrWC+5VvFB+9TmfdVMPJf/MF0BET1TVlPX6R
QKbIZvGhpglHnPpQ6sUdNpTKFlC6/MArBW2Ls7cqO2sG3vTaXV0n7m63BnOV8qdD
JtBHiDYPWXqr24Fup7M1SNmSJ7umddmNLKfGtcUT88Hqq+j0tz4qdNA1xv7J2hQk
pg7SLBKiTY3KGj0W/mar4Ko4SkR0g0dT8lBUGJdrsRUBF/4BMw5JyC/sRHho9LIY
hIZOu6eMFD8MM4xG/4vx9Cn1IxXoF1Pi3w92ItOmT4rBGEQEd/UPoATk3qaAh9MI
eqBqlb2FkKSYCYuE0oIxsOcE2cBOs3nU6QRO63uWoIKuzVX/EoisArCIF+eekgQX
gGcXLGMsXZGY5cOXR0yKAJwYoP0+pevyejs0G9KXpy254KL7mxyZuiXAwK7bklgl
7ERKK0V9Ye8YpTJm9nc19BEeM0i3dTOiCl3FFHza3SohxHnS1wAhBdSj/UjFTW1i
z6qRU1lq8OE6NXL6degOz3IuZ9S1NXJgzmFWe/m/eftuzQA66jGPe2SvADgpYvtC
0UxK0uW0EoDnDZYi6JTULgu99xDFY7RX+Zc8TxYkQ6Gl0Lt9csheRqfej0lII+5B
mtGofcEBSfcyaSOemqKa5+40my5ZQdKw8RYrd+K6Cev3lOk5DA/XZ111gapkebI7
mlDz4W+efW8qG2IpTsR1mGu18RQUOsuEcicGGSXM00EJKrPP1u74Sut0dDD/59X5
waALvLjLyqgL6e8ym1bEM9dm9GWjxdA8mly9OjIJssrJ7bwEV03uPS59AjkY1+3I
mAjGb0XxpFqiKpggBOW8uh8UhMzpNn6AS83XKoZF33xy/8zgD/BPtvdmcs6vB+O8
EvY/FzDSfu7qdAqcqYpEjHO61yAwEmdez/jMDYy/pDgA3MPi8Bmicge408q75E8X
6xPOpudfZlsL75Q/MyxaP4Z5Q5m1N+aNpOGxXmp9hecmvm5lS/k9ToqxevS8ESBQ
PBgV9ORupoFboF+WOj8ov57avU4XbQVr5BvE3QSdoWbQmydTqM5W4vSAXuGHwUbI
A4oH1WYu+Q3+ZYD/1Qkdziw4ITgpiT9xj4Khxv/OoSwrq21N3BrDDRdtpZEEvDrt
jzGID/D+CIHs8zVWht3vLZNXOuN/fnI+7Li4wzv2U6KibAZlyxmb4C3eCJzMmx22
2kBDqjyRqWHIpSiL/nUZBXbg3MYzP0GG/WVCHChToJHTZuxEyBAiwhgKdWNI+2ze
cs5zoZ6Y1CuTYw6GSFsyWF2oBKekXrKlRIQkHf3sqAkbOAuUAlUhlN0brAvT6Pv8
zpDddmBetpTiTIzl9GT6WWXEUnYFtz2cVa5Spb1+KFgmmxiaRgsgQu3t7p6HBKdj
7CEhWqT+UoYEITXL9n2C1Ax528TYQGSEfroCarxT2S6A9Hrzd1JcOD+hBH2COIy9
9//U0TxrCcsR7F2ExLqrASdVmXRud6cc+oV8MRoHKVH1xxCs+CzYqj+wrfh3vaHa
s6ZJ2sW95/h1BaY0GxsMKldqelNLF0pOn6vp91VZelBRbHLfqaddCyoa5d4lYu+J
b4YUZnkcSCvOwKdYEG2jUD+7iOMczzAo3trmTtSl6fi+q8v59+l3+ppDSF/u5TNb
KMJvHWDXzw4UyV01f2LFKJv/WQW6XVPSTzuJwHdBSi5BIVggZ5YJn4EQD+6fqk40
trAq5zM/Whg5mzyTf+TZz6l51iPVx/h5kk8MmzQ6sFNJ6LhzcrZl9wfCHy6/MOXO
smmoScaH8Zp/zNJ8IOqEkiWS34Hy99Nt4oFuA7GNAgOBasTW0d9xszJ5zb1UY32j
45DBceqqqe0XDK7HWGfmrNBvkpbwtKUNv4AwoLbIhynDsVHr/KkzeatuP4uw/s2D
yGTuy48ytV8/yObVnfE2RrR/DdKtYZTdEdHb4NiFQhmxvHJoDEpTATZWP8AE/uOP
O8LUpGuZsUaPaxr+FBxMats79GB3L7af/1jzi7yeC9FFhRlXxI/A5rb4PZ1FqzvD
VbYuLlPMvje2nb3obmZ9fX2wX0kqz3pYfDKsAxJfQQO47qYU9hm6vuCEAJN9s6X2
Ngi1esnx9qcJG/VT+rCRWS9/IynIphzJHmSw/xw91CgHMXilnBWU27gpHsKZdcSe
7WNEOEyFI3eLGPsybHsCYqAIPzQmMRXDX4I9t/0uB60KdyOgoZF08DVMn6NX5Pcd
LxJs4owFC0vJ/1A42pMSMKlp4W0c0ep2nvZxvtjLqBJfy4GlZPgnBIJIaiftwDnf
AcyYcTu+cJpKTilbzb4rwBpOuGlRg0vQmNsxh/+JvlwqgrLwszFy/wFC9Gdck4bD
9pB5wpRnjOmfJKrNvC6Qxw4t1XTP5jjSZ9dU3KpvVWunUPAePKHwTHgYyHnKsoVq
6X+ewRibuh5ojSrTtO8zBG1aXznk0IsTrex77gPzivV7hHem/uxF6oRlwMEvOPnw
WHEr6/42q07n05tJHEL8of1Mh5ZgY3BBu9HuRE6cOJ+7HOfPSM0gfEevt8uu0w9u
YFmKfFsH+Ck/ZwCpZ2xHCbE2gDDFn4ErjmxABM3DbBdbAHC9Wkd3SyJw21AAxrTO
7AWVU6XVA1bqoOu1dgZZT6PtI7zOMV/Xm2Iap3IDGjXNKkrIkZVHcATejQ/SCOWZ
hz9AgF6xMoXx+24KgXgvD9DCzyHmEVpQibqVTq9XNMnVp9YVqGd/jJuAeFNVC+H+
xwfCnYYB5K3flKbYaBJ3SJKf1h6Et4cIkhJJRvBAKR9hlZ3ODzrK43QPtiaRp2o0
jcaHGfunADG3R/wfIplzxEcUlYMSb0MukNSD5U52YO2BwR5u5j6OTJbGDrbsf0PR
zAat/b6jLJcBnW6wr1VCqWS5OtKNCodpLS4hDxObnBcEBosZw6K1ohQ66BTG3dT1
FAp2t/n1l9/ZF7IvzU39PY8h/uUgaKAn1J4D/6kr3XRbdz/X6nG91guAwdJqHJaL
EDaiSj5UKaV4mzSlHtBHQEpdeV3RrW/Urb9Th4os6MuKnmH8Q/Z3Hw5PLeUjNb+y
juCRK98RNYY7fMRG5MPaedluQ5J6U+/ryDmmZJmPv+tmBAwBOZhdPJ9L79rtlCUA
Rg1KZ6kU+WNTITEy2+v9rZd87JIt+aF+ng2GkEzQDDHaHMK9OvXP0V1eGLIHTof0
6JMpqc0rK8MoxRhSmw0BP3svcvGBJg0nD91a6U0IKDQnwNrSHnUZ2M7C1FB+k+sd
EEEX9/c60WNk5scFJqZAernWumnmJGM0dpnoL6Z7U3hBWiAJ8dNfEUQHDtH1fXFS
tUj0n+m1ctmh39VSRoh6iG7mBVsFgAIJas8tXN1O6KqX2wDj8HbGACGjX/X3OMHi
qe5BdTQ3OQ/5gHejcJbn7yYwEyF/osmWSQ0IPvqEos4YG+cj9m2uxXmKuOAB5jFE
09BaOAutqXLiYmq+H3d/d8UjTlSCzylLVeaID+bDR2YPpxtIUqkJUoZZE5tC9bd4
b0OtBDvxWShPs0U1ezkmIf3h1OuD5c7AeSYJQxJNLq+qmTZC7juvmZ2keVsPNVkt
xXt2+qS2ugZxEmM5HOa1jbkXLQVhzVFZySsJpwZSf8Q7X59mqx/3psz/xAOSn+u6
lrMnEpIyMnnYnPdfyzncC86uFSvP5Rxlx18liAB5Tkoe7jet0d/f/OyYV5kEEkaR
Ga+QicZh8tWX6zlqgrDClEeuJXY9cVUC12M9Bek2rqkK5Vru/MoKGTsDy0+9gvJM
TzGDwb1OlV21AUkpBOWgsiXj8c+eM4POPFECcYDh3xX2FFeovzrClRznDl4RAao9
1OyehPSKGn6N3Ov8NO0x3xGVpFDBpQG/y+ONb5f/HcvXyZhMd71d6gzPeWmf1bMc
P5B25PrnJ5BYbNxCzEBZ89BDMaL91NMac7NaDzJzleX0GqZIKsKlNK237KY61Ecg
h7FxLTi+Xm04w7FN+mnKlKe2NC1LLgwUIwFknAtAIWzJdHmfiu/UZK9zVONvYNBw
H+6ZmlgBT4B/4P0ED/w/6r7uy5EDOB9O/d720xI4y3q6qTQWVJvJIGVmZlzLo6VW
ytU4Cwmg973mYUew/z8tbbnIeM7JOM2fk3SQ3LZ581pJ9Jw2eGXd/ozymwcMdMS6
YrFZODc5G85wP6ow4En7cxIp/yw0ErHsaVq6e2H2SFivgfNiDCgnz1dEdgBAZa+I
f3G9WsKKOjE2Iy+613QrD1i2pEJ4Tn0rfUKJgyy1MIROA4LuaPDi3TTM1vPnMXn5
DihViIhCPK7oeh/aZW5G6vxvYmOCUp6Azv+s5rKPVq31PxxfFhqzN54+yVvHBz8I
BbDj8vR6xE9e0GH1zhUKeRMXe30JXfP16TS42pwOtmLJ3kZhj3WFIVy3FaPESoV9
mQtJreusNFiYQxq1OLsXLiDLTJeywCZ7l8uP7IU3lLDWrxL2V7HPeBpNGExnDndl
tbNHOH1dznmNNx8AulGzqCBUgvM94QFnsqtUgKAo+uO3dbcJTJKmuwPSYUaMAaCE
cZ5PE3xdUMr2oTihEjo9IZGvSU76Pd/kM+5Ar8Bi1noTg4JFJrNEWSxjM3aBHyzJ
oEMC7h2B9LVDPPdtaN6vzrqpXWFZdwQNGRltgx0/C7vOmlKYhYdp/E2axZ50eB7E
vFf4fXzdt3DCIqwDwJVZN0sHq6OGKXCfcGivOxLjV3JhkaJEjPzhvRzBtD/nMEWO
z9d0Wf+tF3dM/VVq7uaJ7j4H/oOhVPda151jAngYHGQNQGjhyRNACmu5G8ShN3SI
/GzVWGpCzyf8g8QxPW5aLIMpbbNBnSjaOaRv6yWeP+KCV0ZWjTZDnCmp3AaCpxqy
T3Uc7OAbO4tlI3MO/xDL3wVw/Pi3BtSfA2zHVbkqiLwXdbyQ3t0zjbykOcanrZOf
lJAjCN+T42bFPWi4No0fDy1fLxu8wKz2mdXW/Xv9qb1pnflGXwgZ5tPIxQByVlix
9CJ6chNntTuj3561Uoqjszqi1oixiEUGS4lpSxSOTuPrreYfgoEbqC5Y0IJAfkSz
jsg/TnZyJghPTZSodaTPSZSM5hGykS7ghxcH8WtiLQQRkdHKqwzf3xHuuqJd6faC
c+zUqh41SCeosrOBKgaIYLu/dPYiwxvl9/H+PRGw98819hini006CMMiF18Q/htt
ThULWvoND0Ub1R1YisyXjn0M4wU2G1dXojO6PbaGSWK4UQuer99vY2A260A1BJYJ
I2pYcKoWmXxDXfM0Ny7YuOL0wgtHpup4u+/ZBNcDETSQ6cvYxOcT/wneiPg7Qpbm
01St3JosJIfNiVT8dxyCjrmmOaVNrFdm7dacqcvIPyiWv6JCpyB5R5QPiAMwm+J9
n8hhAc4POxaM0M3SCqjjXiY7PhS/+rIe/aqnapm0ApjZru7D5u2rl3UKqTYW9YT5
+/HeUmkbjcLOZq92vOik/mqocdkbfS4QMySsdmEWs5q+KAmx5zS5VGcQ8rSAPwEH
a7APKvlAzvSAEnmrOWev0QaX6skNje5HLUcHvRTj7o3SznBL46YdivUkj+bSUDGh
0R436u85Mvbt10nJgbcjwuMR0QB6j3OZDHyx2gzqSq+F5sQ9wI8VjzgpEj94NeuE
Rzta/Gavo7vjbOwaMY9ijgITYC+qctSddY7/Bd6cWXPphKoa272rrigR4fbP911s
8xaEebkNiZ31YY8cN2eVwAeKQcYT6EKZyEO1N4giU60eE5PwyY/9vPE19Y1mbeCg
pG1wCjUO4RfN2oMwvAeupyGFHWFByUrua/llWivZc+pKUoxLTxfWy2JSx55cOQzN
hiN1dRtNPqVKWj4kIdf/T9MWNaIqAANjrO6aG27dLPYBbCSoPMg9GA9+PgfqAdQt
zsrFagSgjI6GnG+bQuxgvL3Zyc5j3j/njy9AAMam4zCaeYU4pu/PCjM8Wwn8HCE7
envl78fcfeRqRppNEgU1bKJEa0T7+ENcfMybYrFKob5gAjjiAqD2o25wwLg4S+mG
SBEJ6s1iC+s3Yoo+arO8qRHxFCeyG7A7oWml5XkB+YZmhyHcw5aqkhGhX9ZUeE9+
3kykvFHwsedXBxt4ENkJ3oIeOYWXx3uohJfuVVkY3/rqELw212XV1AzhzAfz6Ql8
x5yqzVzNKxAhrZCXQbeAZiN3X84jr9hLydvrlekCcNRRFvq2rIg6U7HxvVlHYLMh
yqgmbUWLwM3FyS0s31YVPCuAF/HAXQlhwCCkkrTf43gFte7wbpBSBtjVeHdmA7f5
2x27wFQ0y6z2Y1jqxG6KjURL+oUkrxi4hEJ0srxvvLFdZ7saFwwsqzPkhQmtGm/P
+KdObshU32axlreqL3OPzBi3YLGDi7HEoE4tvEpYnPTbVtdlScvX2Yild92vgyNL
kkVfXTliMjT5Zbzje8glqfjGWfTuDaXhokz0NEqWNYnwY9Sc6tQd6ITRRoq8sRw8
u/cw3doHpjz1qsetI3LacbtlgRWC3Ks0kdRHhJzwDc1e44TQsQn4KIGoyUzgPyeE
Gq8cPKpr7pQQRnj6lBmVFEGUyF7s7Yl+hnLjTfyiWHnI2RdGQB1nUWBEv3Fj8EVi
XtZzLvD/4Qo4BuB72x6OMqXZhZ67o1mv55jI0Zr6pRTL3NosyqN5Z0mEe+ETSZ9f
/WhANSJLfn4hpYJi/FGsmQiomlsNjyWPSMeOhYvmMj9Wm0xRFMhm4STfWxQJfzw2
2qz8+28Z7rLpFcd6aGCJOF+BMLyUgzA4ZUwhCoZooy9rmubVofZ+Fnqy9IoLYPTE
JClKU9M+Eg7c86GlTCkdnXJfNePq/BX7Rh5uSk14SKGZcnpjWoi83bV0zqIiWQcs
31XcTCT02fmF2fjiw22yRbwmAuJyDbm4ZWYL51pU7HMmOzVJwHCfP/3cuXBLVIde
NASm5NsI+YJSvFZO99OtfuKWbf9+kAWlkHnGam/mEUw58y1sZLnodlMZw0BtnMmF
+trR/N5hYzwgawfSuFfJL8RfJ0PIOd+DAcmJzC23rsURK2Vn3TcRQ8Wfg0850hke
hT395QvG7oyMLGuLJd9DEJeJTufFi2G1Hr3TehFOjPz3D1PAujsqy0zeq8oj4Xx0
Qh/ddsgnUx+HyL9GgzICUOprm6X+XeY/HhxSPYh/yJJJgypM9MTaZLDGTt9eb9MV
RMpXTg1RGZdUPtdO6WjBc+mcfN6LG8Gw8Rs9s09CQ/ib03UYMS2R9X2Ip2/nVitB
NAoFqzRbcp9rzj6TYfHa7+gP7rk+ULisNTE3sOZL81AsoNkqSvikoNjOxfrzYYJM
ywhUtmS4DD5/23TggqBX6HMYi0V0AfQbbdnJazM4sjLKQpZOsoj8Qcin1+uLOCqh
8ukg/xKnnjQAUtyDAyRoNrZulqiCNxUEbVAcELxEnU5fcg7XcVL7cHcKcyMcyIhP
1sGo4Lf+0wa4GZ9lT4gn35KyGizO8oXVn6oXEpl1QPNDZGVYG3oymlEkifU83Zjd
NxiP5BkU8vqKaoR2egH7WbBu/tLq3iH40Z+Q5nTTmKh7OB1v/6i6ILKphmGspdgv
64Y+41p3ZErasxMnr3L7I0bU88vjDwibL1utwtrb6Msf27e1hcrHQvzF0K4ME/dc
aoXm/si+UE//q1UjRPdy4SybkUB9PnIquckSXEyKux0Q63xuJfTbGdCd+fvQqSx8
ltDoD8kMJbOuNbr4y9UJRGTqxdbmeIVUodcSk9YaoiHAvruarqjgD7jxIK8F+HC+
36robbLjuykVnZ44nS3MhBy3n4OLsAbpS2Lk1cVoQIWLvm9ShR67IVcmEqJkk24k
ygZQDHUeBlb5VtioMkaxVoZyHsMDodaLx0bKnNINfq6LWghFgZiL+LEVJPMc+fv8
06H4trTlXC6oHcbBW6mX/Lel7JyyuK9Xn5eAJ5vyleN4htBTwjTg00b4sBxfytrV
9WSC5gwS6xsbqz8MuPV7NLAFYMd67IH4iLA7Hea8p+puPhc6KEeAQxrCw8+4Va67
5JJtF3WHTTL/dLjEYwBQ5UULsINRQIr7F7mW7q28ZKCP7w2efa01TaM5G2gGrev6
9dyb08JCfCfRI7/46BRoGe4RVjZ+m3mV1t4SWE736113nsjg76KfuodqIyESgMYS
8hs8/Z9QVy3uUsb6JBX/KSXGtGwFBqphcppkZeoFA+6vjHlQnc6RSYN6lfRVUSkP
l0Sh3U0WS2IQ4ArBZhgmdYRctmWgxIz6d7pdznNO5epqZqJdMmSUDq6cQRURvoQL
UzxAkdkouPpqc1eIdDetIWCD13hoRzzFOVQr/mTQRjrsnpdx82BOh7scbnSYq1u+
oQKX8Cs5/hr5WXX1So+LGNN85OFZin7xffG0gn+8lC50/jINjK6j0gFlgvKJ9zOo
3y7okHYABIc1Rsb136mtaXPMlTJD7A7BJoNWa4iglicTvi7FN1ocrC8Hq0J4R/lD
+43AViyGBD2lORkRX+ix8PBbvI7W9mDvGp0IDHw5GNIJpnVvRvl1qxxeh8Wkdyxb
lhhwM+Ks7nrh5pYa20dTTDr90wMggJiNPCfKWP8dOplQIg1h9Re30yuHfIijRlow
t4M5id18rUZvnkNypYGE2FLRTtQUOw9FhwZapguZdSeP0C8TKfLLcaVz6F5nwguj
JZgBipHvTxESqgxJ2IY7rxWFuCGTWHKKxsXubk4lJSE1e+hSRTETScssVu1vZyPw
oZsvy+8ERswCY7f39Y2AAlFnVow31WSyMSxHbzMNxsrRjaYNi5q7bzX592BMFcRf
sanCOUeW0p8Tr/t+dFUCo5Jlng5b/8SRyj5ffumi95rH20LxUch2lUGEE0OTTsAh
Ks8P0h9pgmbxsQlsolVVQl0AAsTYY1aMkBDav81Jj5o7qigaIQXr0NKhkJSemzpD
vx6mRkiIiw4Os7cOKDIYxg4FpQOsw85ubd1FbOpcnrcM2DkRHAslCMaGeE2BtTdi
KyfbMBxjIWwpwFbkAHINrughwdcZJ49YBmj0z82Khx6ScJ/bb7ezKeHB7u18moNP
nb/kE0L7lBRf03pEeuMQdhMJG10VlsVLs0eV0EM+OZnreQwSp2xSfcWNXDRUc2c3
TtOrfWiy40Xs9ETWPAi/w9hW8AFAqjguraJaJ7YJdxAK6hyRCyokXoP5QPEqPQW7
OZ3A6B6C7AHkrCGe39bx4DcFqSVZZ2aSBYuX1zcMw98/VmRCJXyHjECuGBJvVERe
nenGPkfq3jl7/XnCnXkn0hf8f6wa82kMn4kiOYAOGp+q5xlX2Phi5/ACEGlAKz4g
a31AWvUHV3nsCq9EpygJWOyzKbN30crLVV6pb4K2JZjJW3m/TDsVUrrZsYAYgAza
AdseW5JUIHenmQruWK6C24ISBn9wW6/uHNgQkwdqOK4BotZL3r6YtMMZi+ANYLXA
UOQphWoWsV6viRjlCXdyreSdqzpcehC1A5IqkUyPi9pEs1SBD974NFanIlkyPsrZ
/Je3Facnn01v9VqnYbtTnBaAlxKH7BKRlO/m5Nr0jPa387fOjsR2Ul/Hhznk761O
u+v/rw3VLLBsmUg/bBucipSEDTVedB5j8wenwvUS92EaT61sQzaQZZKA/8XutPOF
+RH9+xRCTBZ4OXXWIeyKby+em8xthYfMcH8+cAVctbfBZDCGeebh4OtHqPB2jISb
YfrQD3Z0o7/ZEUHR8tM376nxNT8Kw9i4AoE039jnYG8SJ4O50E9crRL/9XEa8a2d
g+Iaf2OoRbLn8CV25heOfrNELSmk6TB730p5Gjvb1rAuPyJL8PsZZpYlMUX7veal
q1iobkzAyPjV5/yf3is/f3KGk42TjyMLXWVnrV8eQrFBYE8XMTnbwx7eg+ZrOkNz
AW+qo5b4n+kmMtDTJy5CX8kdVL8hG8o8LPNyucY+zwpzrMV+GdXKF1c5pv7OPRL0
VcPt5AUlY7ONl53PqofYiuQF8snRkqj22NKsqwuUpjnXE+xTHvbwy/PlOF1Bh5pA
+l8zbFHhCJrQPNAwqTnbukCBT4ZWWpTcJPkjAg0ySD7+fMHHHo2MdGqSv+keH40c
5jbYJmXD+EaYNiqPrdXtW9Aw0iy6bEmrWG+rTUrVtp3HGpCjcvyRaZTYk1uUnXqO
1xQtrbT2Okgwmg6Iowbm1U8OzFNVp93KK6ifLwRgUSh2aNYMJp80VtuJQXlJqN0q
nQ99kdZzG1t9hgQr7VhDKUGC9Wwct44BTNya+mT0R/gKARFQCRznZJEaFWxi8Njg
JhpxBWNTrs7V8kp5kZwLaOoKFK+Baf62i+XyP0f8WuohGH/pgYl7HgnCOf9mzbAR
mn913KB/3bJBpPxePyiKlSyT6ErSm6ZYR/wXr4ffK3w4nkekpuMySRy2nlEQZ5eV
BBIwgKkRJeM3RT/9k/REJlRFhzpeamd61WLufSF+CKkG9h7B7AnidwFk/FHP81vu
RTXWBuxlb97Lx/qarzckibafF5Vhi1DqpebNr74oC4xbHKAcVb3lf21DWEf3sxk1
Y4fUxuUcV7yC344IWgHlZm6ptfMNEXrFW1Ttn+W+ts2uPYAPXjUr/oYE5E77mUe4
V/QFrwV2VS5vdd8GBATNj9ZQt/VjqdWuOkkebHlxmHlCjccWimZU6VQR4y1kXlJy
RyC50Gn7mHvQaexRYuj4gVxRQHS4E1ZYG6EAnWffvJOS7rHlPmU+v2C3p7foddlT
Nw5iQ3ZCq7taNx8OAuaT0zHJMaVVGj87j4nLKMxQZicl+uySP4IvAPXPByH0mmU2
nBQC+2wzRr3a7mosgbCFICdMvF6iswaLnaC2+7aanV/AgjN+JuBJcPfaGKcLTzJg
Y3ttHiimpdJO4QDpucFmWYsyeBSue6mtS7G6c5GDeRM9EKibdgovo7bAllrW+jAK
Lz1dAf7NsxQR+D30dNFaL+M+jQ5MLzSowe1Tho9XDkprB36C8Dbgtu4iQY7yZdok
cCcEmDr/5doHbIkhN+ZXhD5vUfeE77xNmM5hlOJ1q0fLLdF8GwzLa6VJ6O6KkI5s
SnggjBD6fmV9KGIZ4LK3XPyckgaU3GR41XWGYDeRICdKKVrXn2fN5lE5dR8rTP9N
HinRnZZOR1nLM4mcNDAEi0g4lp1vDPAqqiOm5M1VuQfuSoBC3MymmJUZzWeb4WPz
67F3hZ0OJ0STYiFMqWor37Oey8RfMolHz61Ct9i18zLCiS/2sdBCbE2E4g9ZIhCt
hq5/MTYH6OJKAhxlDaKUBEcwXaU7CyV4rSqtMUcGog4AnZrKyBT3y6ewjSwi03Er
o4uVV5GzZrq/YJRnNdc3yr3ygPAs/SKZonfvXEpMjdPuuygLYnPR2g+RVU32QJ6G
b3lg/cyIgEJ6uDsIxS4DfScb2oO0iMMxSDkJkmPm6bbizIGL0Tq8bZhlkHekJ0sW
f0uevouF68tICN9kfWf/VTJazjnrx6sF+OOjkdSeO23XaTDC0qDiclRhiS6bAUGb
SMwb7gth9tTYVz/JilIG51OQ1vjf+UxygnvMod/Bku6bXBaN0S2NlRwvCJ2eK6Mo
0BhO10CZxDq7i9HDYgKZuNwnAavrLyJ0ZH60uvt519PelP9OPL8/PFG0gxqBQyGB
zuUtzz0qlxk6wLSazH/vHiSCltfKT8tY+VHG12SiWMgNPG8AsNjfUtvIAwPsku4x
t0q3Id5WVoCrtvWPeuiBx9D6rNvPviIyJ/F5B2BIb+c3o8c3JlAqgTGRmGROPmR0
HKIEC6j/vMKkb1YzBD/MENZC3EsTlU/rQHhqSB6jOBhZSNgo059jxjaspWGtXYcG
YPEZclKjuK8UFHR5eJDQ52EVdgUYVXOXt8m+p4jbcuMKbRM41CAVncvPV95nOyOd
xmKSLiIgAxTGtUDxL2heQJ44vNI0ZfMNkczbNoBDPFtqV3KgpDiFHe1kHa6JVMmx
UOmI+XEMhP994qMnOZWjmWNcv5HfI7h/cWfYPNA5gAKsHLx//vyzalKMlbhVNYaP
aTRrjrm3q3wFMj4lVxRF6xecrG0DiseQRLjOAedGuvBSzokmkRY7mQRTWZq2XS0D
A/3shp8R4Fb8/+l+VoC1BQUKd8nkzjCE/xIzzU4vxsLDzdJ/pW9gnrYONgcFK5Mm
vLrZtXQjqoie8dJfeP5RBw8qnktssrDlMtfTA1umofBU/wFy/9jbhHPyPpOvDjny
yQdjSk5jCgrflQPLfX3L8qBIdnS0hRpDvoXX3xzHW9Q0+p0zu8aOFUIXmtrBDyMw
E90W+abUQczQvPwJ7dX/H8OunXeuJjl3NLBKQiZCb1tb6IfzAGIPWMyXIr6XpVly
NSjqIWAgyd+dTHwVGmJffSkzRgcd4NJt0wwZX78XBKniNuWQ1qNITTdMLDsKxXkd
gT/NZzHoxxfTmRAHVUsP3rEc6ORgdSinek9WsDFicmqeoup2oahE5KRO9X/ySm0a
Kxst1AY/7c1vLOIlA4e/zvggKj9vl0DFs3vpM42oPTqHXQuYAZ+nN4/GJcKYRkz9
dmezi4foEkZg6zCzyeOSc3gixTs7dLKsRSuxTi31w9AN4pB1Ec5RoVwrlZ5NqEgY
9+LdQ3gIz826utzqKEagtd4VfJUuIFvSgIH8bJYHCPgb/bVkl8+Bs9yJc2d1qB35
y2YnTp640diS7oNo5fdrWCnav8eGsIXd+bv3WX5/1/MLDjjUkDwPSHTZP5NXgkoI
sDDKZyxv0C0h+EV0rBXtIuxFDxr77gM4eq8pNivsgG9ScWiCzu7+ry5NjEJTGiJP
7lFl/z3F7gTTp84Mr8zttGy0jkoJuG4XYJb/XUSAWz6V4ZyltAsdWMmtq+PBqcjQ
ilJby84EIpJn3tpPKcclp/UL9Yb6jOVJOJh1RhmSUVBE2j/6j2naniTPHxtND7/W
Cel/zBh5v0aTHjBnDLKWIyeSQiA553vhgTBXYu8y/lfk8TUCIhdpvYUwcNmqfE9X
kKQ0XCFZ7CIo3Qul5cJtYOaxU+m/Pe/8S3IlvTRomHfhFluhHReeHIfSDg7FSV6e
TmpIY6fMkNRJ+0Z0FX4gNedRgb6ehCMXdgZaJuw8yGYOrrP0pGK1zK1F+GPZSV54
EqCQ8LY2z1arw5F7g4ve4XggkIUdcrJlDu2Jmg1qqwUrOKIX0AIRNavUru3gz5As
91OZEakMm5kzUZVc/IL6T70r91dDa9II0OwhwEqLAnDr88Sa7EgliKR7yhzwBlVk
T/t55pwK0xIbsnHy3X00pebsRg4ewVb7/Fju1uYZTZuF+yOU7fIXFwCM+z14njvU
IoWT090zElY70Spv8s0ajSYCdT5Ha05ULEm3eRXY/MTpbgQDqz11+3ISg4SPqEig
ccP+hA6hcX/sAAU33ORFSoJLEruAvAWWqbKgeQi4wzNVbA3OQnh76wbuQrzDnQ63
tLG9NiudoYOITYgH3I9lW+iY27MvPrne7Gmm5IldP1vVvzl3bLjR9J6m8pm4R1ZQ
fmQmep4C22H6ac0K0y3RFxlYFP8sibVgqMGiCyDVANxJy6PtSa0/9Epgy1dICv5l
WJ05Sb0O6J2fCIVxgN1y1VMHjkwO/kIUHGYJ0D1gQY3y1W+ujaga8F2VLwv1ExbQ
NgeJQxKIjKOXBnSXqD8WOsFF3T46ZiA0aOTLLgMaX1xjODpBUjPqlHdvUNdvPjPg
yP3BgH/qpG41Bhw1+v8KjJNE67GAOkIciVQc54oPBJZbK617VlbTJsuagRjk8oIK
L/dkENzTv7nMutS+rfpytaMSLVdg+oQJ6ii1ZdW8zhvvw8TcAdV958K59nmEE4r+
rEGK9e4GwAbxZttIdQPPM5tHhp6XFGhGB9cvZUKunSFyJ/Xs15/M9TTx4tM1pczf
sRl1R9VmUtqKvu/29tcefnWBJqDzfUVdWH22P0lewJaCPnWswDgqEO3R0eoy+V/7
4UCoL/xV4Rz/syUBk5ebYaH9+32G82bUDD/jC1f/6q6kak5bp9LPBTrwahX2Yc4h
KJgIeuKVaKhqUS6tX63M2CIyxKuC1qdMs4KWhORMJCiBgggQdYxBIX2LB+v8WyQV
K5LHaid3mBAD+WyHfgKahTRm+nIGTr26Lgr10GyGQU4Fhhp7yfpDLzH1TOYXzJvp
P7f05O2mFBbsOq8/lunwCjhI2akmP1Vsyy5YUM8VVzz4PWGuxVqoSGmyEw9Eve88
8/pMtjjDtcAqdVyGTNVwhDz1E8RN/LwEyA78hJ9WDRAIWGEmm9bs0xE7giT84IsZ
t5gDh2+2QbXww8+FWt1qYxL3+jFl2J9cU3ch0v9vfQxQwBdp2LckDsQnogfl9zUB
T7SQnGDbs+aVZ1qA7JI9MyruojyJfJGxvvFoWgz0OV8maMURKz5aLqwoINy+JU2f
fk/SO9ossZfbabz+XQrCdaUdE3SWj5qgvyGKue1ZPp+QePuGxRvKy8eY36sCpKxk
8lKoCmyyNTKiDRdA8KobPa/D/hIBYW4vQZIsX0kGbPHw7mIOs8zU96Hh5DR1VZd8
LoX+VhjKlNeCHLz8lsq+4NF1DDg/C7pSYzwT5gruv09ZxIKHoCFDFj+0RJMF3ai6
EEMeAv1jnyLrQ2O2ftyq7UdMeLV2gkX4Db7FV3JdLUjpiooOR7yjfcgljWCb3cvb
NBl64NmjwTLOGMbjNl2DT/GYH1hCZ4EXi19ADFyQyhGE1d9ghwj+YKCQdgYp0vXD
MwZhfsIG1BNaKHSYOkfeXwiP4HePDc5RwfiQTl4MyUDVetHl7h79sWwcnIoy6Rlo
UYeahlivQlmGfRz9G1WdVIBS+pb1krEoUVFop/2cQH0BwgPIy5N9AZeIyecNLbpk
OCBlbR3RLwr1B3bkgLOjLxeMAD81cxNv02qKGUcE+bzh8/SZUcFEFqfwFSQCEkKQ
UE49BGMd5m2ZgV/Y+dQwYdE3okyNMeh1jlID9GiKGK/0KwfpYMzG0lMgIOjGvrjI
QiDu5pRzWs9y/G600LV7zWRoT4VBoYzZXeSwmNPB1PLj6FW2v3UO65RRqL5eX4Gf
dbDomhHg1zn7XY/atqMC/UyQwECuzFXvydgv/CXlZZVjVJsIuznyzY3NRqUBkxh2
jjeLocLUd1HynEe3af47VRVJogDdJ/PD/lrkjsN7fbwxvc7u5uoCaDCPagZR1eVY
q/t1mm21pkJMCcnrd/9Ok9VBNkVqun9hfrmM75RLwzTkOFmyhzwVuycI3RIAG/2O
T3MpCuTfHLSvq6mHmG9nyNZVnvN8z629tAv4P7uNLuDsoY7AXxEpYEU1ijBDb14s
QcIZ9QjQb/1MptCnc32rFK6WwQpVk4TFGMQAIhYZhjkIntCBK5YcTOBqYKfCH+su
WREek7r/gGWgKNROa2l4cc2JaVW/aRD7zone47pOSi0vfVQNW7YontQeZWAw1xIx
AdcRSc4H77GzuCgjMubVzLtjCyUgvtjbk3XQ8duXaheO2mJe36ScUuHcKghpIJWu
SblNyYi6TqP3zmibs7Dyi7gll2DhRWF7LD3w/Ff6sa7kEKvmmbpTXRfNvU02SYYI
umYIbMEjDWdns2wpN0JQR6FUeORHxoQ7oy6jo/1+ruWaQfJDVcVAhNaVFlSlQ52f
ModSdsYaM/yVXWlS2iFWXnqBjGtxZDIoSDqFf0QTmlsEVVyCbxLbZdxEMwz9tlyL
LWRJOFyOVOrfZID3QC0MSxwGgJYm6b9AaHHLsl9fbrkJWtriij6yzQeLvrteSSP4
/40E0jMi9qTUPW+YDagRLHd+xLdVGijyfXMRC5uNWsGs+uyN84alTCH5hwJnwAws
rGG6EA9BycvbgdGBTL3PecWGLR79ayRG+cNT2nVEBWOn7KAR2p9kmBvKMsh1EEaW
NXJPstXQYuAsisXx+2bPco5Mr5Nk5cdy6lC0bEP8CE+nr+9nqYcvEr4qqqTnerrM
pw84XamluznRuQLUti3+mrD2bwPukP12l/UinEe9k7bwlf/o4HLI3sPuPk+k3SYg
9XTkksOU4eGLY2YYaJUkaG1pIHvrc7oH6EVWJUl1oinqn3ul9lbkx7Dm2Gj2W2wT
v89jYuKva2DBJOt18EZ6dpnHLqUmiuUtkg5iXDFcTJmQ7a/32vEvzLrvtJotjQUI
R3E4fw6U9d9wlzTLm9lnNW0/w7u3P1K2PArfnRk5luHSv3MivHE6h1h1rzFdI7av
e43iEvouNVWc3xSIv6kfkrm/ACLHrx/RgjAvQwGl+4z65WjJyPl92ksEwm1Eb+q1
dZ9UJnJ2UQO7Lez1PaGDWGaoUtXIG5+OG37+dJHsztGzJkIvc5QjBQKTG+heJPxL
f/pW3z7VGf1feDFS4XZITZEvHENsjdzlX0B/ztw48KXMSsD5C8E9e1qNKZlStCfv
wTO8GQxtOqeUzSp0sW/91REdOMAlQ9TDQ4iWqvJrkNxcC9mE8PrQCWwWuMPp5suR
6HQnxTo32VpX3QOqj8SErBzF+RnaYKi4f9OBw0iO9pFR4pIMt8zLMHZglCNwcTyq
m2CreiVIZ1MeR3zTXxypHuaiWPwoB8yxzl7MOIaxdwTimIWMySQ/xXndmv1ViozZ
9r+Ae6owDD++U1vz8mcrwJMK7aDsNcfcLnU+JL9IKLI1fxMIMWM8aMHbEvBGeMW9
v4d/Yqi4On0CEWwEld6dzNVlHtsYBlJAlIxCVKUfNDy/Zuj7P5jjXnYeJU/eNypG
P+XZhKDvHJ3c+S38F+V/QiAo+JUmwHLZn3ouOF3G+DFrIM5Zq+tHVvjpPJBLqybX
dALrQ7AzrwdKECSgrPThcCIYqigK1WADJtiZuED0ngFcom0y0d0PXIT9mOETEvdU
b3OvRE0B032q1z1FXz3RsROxzIommORf9hMt7Gq89Nwh+AzF06mp/2s7hQglp+QO
/w2Uq3bwefFLgoTeI1EJOAQzfHu9GN8H6pxXWIGRlpkFhCoFujcvi8UIFAyjeC1Q
4vRcivMIcJykpqw9oWdwNsRQnZ77uJx5lq3ojvafmKdln33jdIc4E4EvInGJXwQ1
rzufnH9oR3ObVojfad0g9yQLmiYT5+mJQ/cnbReVOwgLGvFk+0ElOIkdr5ZGfzjw
sRQjGw+TheyXnDxXt10fK5vVuvRoZa5PkxNDhv5bwt8Lhz5wZ8v5KnDbTmNvm6vD
BRBbfosbz3GfSdZ7NB2tdB0dyf2BesNT5Uj3mCleGzOLDhqW2qbJun4PUiXs5kvG
AZW2D9WDBZIR+GDtZQivFEsgh91F1Jl9MpukFAvlroPbg7O8Pg+MJ1pOqGpTLx69
TxjqLryJoaBhqTCrhX1mxhbIP9tUVlC1PGN1p+e145ecdYFfKA3yz3/g0unTJ8y8
sBHtuPDJkf/0xETeKM84Pk5GHjFJY1tf1L9RDlcC19zy3dIL758BTO31Og+J0QXQ
8GBxj8TI/aCH4oKa6NyRX7ToTVzIEXyhnk+WYPjwRT3jg+VY3yDS+K14WwCbOdlI
mbTcMgCgr8cq8iz5yCBA0T/Hyp6CjuVkjZ3z73XPrOK2wS/lJf8ft4brIraJfBR2
MVq60cSt43ZrP5SN0so2ouRMPRm+IRMjHwvfLfa1UTZ0gNi5jokZ2knkHCUK0Fo/
o9/HiKG+gwoSHJIj5cNF7ATC5LP0ief2XoDcFoHPPZUDawd7+4QUbywrJwslSMb2
pRZl2/eiJz14v9LmRtFqA0EBoHiGdlQUTYNrkVhR2UWhYce1D8enEoY4bavccpjZ
EnnlOXMMEDVghMjH67KZnHq1r4yZQClxmZvVSsAvakJ6Q0yKFq4u4R/OFxW6+2fv
f8Qc/CCzlyJ/AryRouh0ftlHoyIjQtjWJOwasF+uxS494e5UFXPnXTZN06tv8OGZ
dzk102RzYY6Vbn9VnzyueemhVtD08t2LU3wS3HoQhGqzsdQi73w/Jz+f0LGPgqE3
6E18R8N62VmOeqlml1uqp4bN2Bgev22oNLgpQgS5GpGxcDPhSQBhDxcxVoCOb8gf
orlJeLwnZI4Uc0Sk7QsJr1sGQqOjiEdDIp1/J46IrlUB8V2MeS3pVpJD+pChzRUD
zzGnw9IO0EZglfuB9IJlJfzWawwQksQbEkLXw9gU5KXlIR9aQ6cS2kN963nAUUNb
1rA66xwcCTWli7C9zteMeO6IDmxcQC09wRbPw5Wder2bEHD0tsiUEqIu4Ou3CQUl
QLVNEcokeYxm697HLVIOFFWmeZay1sbzMxvJA1JIWGJTUtBERnrDXRks92+msjxO
eZlVyAosmT6ucPusI8O7Ozd9vaC4e0nj0+IVkvnZkdZx+OczG5L3JlMzLzJe8JKD
E4LAUTyfckxmbplPP+z7icXVNEp75oL8Zm89FuZ9B8DuzmhKI8rt7LoW8dVIL9Yw
0gkNB3plc23Ks4gg+B2CIqxfpNGQNZsZ7yoVbOEJmxwiEKjFOEZfhCyaBS+O09xs
vfSkc2UEMIQhvnFP1Bi0SqsXTpmOMN6QGQEY/XN9+73Rqs+/zE8UuDZ1QISXnG/5
MII8g6bplIyyw+9yZ9ld70oBzopqETc9dcMERPWJPCDQNxaiuhcKXQwSCO9KpVAi
Jd8qPz4456R6b78IEzDTjLUuVGy2qvVDC2Xg+8F/4M03xdmBk0Mcu6ACJXdIlPO+
P++8e/Wl/xp/is3VCQUnIM04VZ/0mMxVAt6tR+unTRZ0NAWjHRWZ7q9bwRqQuLrU
igoVaHMzgo3HlCX5/KvcWEy10H+EteeCC7cL4hrku9q1jjBElWeNv0bH6H6qTqMY
oWByBVjBIu5M42bYiWeDAcdIO2PRPG+ydij3G9rAZn9wgs4cDgI/u3sDroUQc5pN
O3AKVqr9hxSxkJVulefYs0m2oIuQw7ur4UqoVO5WmNVZWoXdW4/1JRRqBOMxAirw
eIA0bxQpuCHor1L/Te6Fbv8Wo34xKQdZxN2R9t3et0ZlxOc7+JNhpIWnqQj5u3Zo
G4jjgGRgd2GZWBYeTwmnCu/j3cYTKHgolgTFsD21WWIzkat7cr0voBeXXPoydWk6
jpcEsin3wZtKsphnA1v/T/xvM+J5xUZv/D3ms8zQKM12WSkZ2yhsINBCReB+gP9A
zT50cZjaL7Vlo7AyxOGOkbp1/mAOsn8mM01Ts3MMMlfvgUEmMJFy67VKeM8VhVve
0XQeVJdbvRSdl0GoR0vY1ySOG9e19/yhb+do+dybljA9shgFxFYbKuL9cD1kCygv
+XOIqFcd3jdmAPPse7yCMwnyCyWHHh5l9UkWA5Fj3qQEk8jFdSOb5gfNGA6reTom
yFsmo2X4cXuIxBViGVqzSbeCkSUIfKnKyIMFraNNaHekAlT830U7buYHRlQDRl/Y
QChFD2k1ciy7l5XVxIDL6ac2ddT9eLlovEbrLtFnApao4RhRSlmdpG2B2HbswvjD
gopUYhpGDWpApYfIIRjt/WWmxQ9A9yKBXmVAYCd3OKcYpWtQZc72Je3sJhFTVaav
LrHo+XtkMx2ER4O3Mtmdlkca8Z7Y7tIo2pYC0nh+GbG3NWu3eYdh56lAKfq5nF5n
RU0yTqyNeNKi0fYDjSP1wWXpT+clWfPdZl01vDOKQMqRI0JD3hIzygaZNizLroFy
WLESlpaDyvuR4cSOPPPlJL/3U1rTV27c0BfiBubZx3F+LwNRi0nFDT1RmOgHf3bk
J/EBUv2OkIsmsX/LDs0Whr2auddgoFIWCej+1qMRSzyGbgHNT5hPq0QHHpD7GHi2
/d5vGUUNd7XdxPc2cJy0R10XxcbU66TnXtmNpPrkZLp1qmycHr96GUgufXg2YlO2
rkbppgnHmEnsZLcidqXQwiCGYLbcFt0jSfmiavNQJbzmN2kE/yO/RPxyU31buvOW
l8+9Q/q1Wne1ODSpV97/gYHRVYYuor6UySeezMjj2PmYW9nEIjBh6TFWgRcL3pHm
/HFeAhulg8kd4RAU8GOFSIw/874mgKWpGJC7TRP2SCxN23OjPiWe+ei8yB/7j1mA
SXnrylDsLR4e6ySji/39oEJOjgm15YlbqWOEbUqL5RzD4TJQ/g1EVdJAvG1IIvZh
XKjHk/TtrkCF/BICoYJxgrZResHHl+4ykOp84X7aYWm9aDDGE+uy4nxvNYrPSuV1
wC5vR05UL9KDhc9kLfOv+kB2tD6tJdomLCwuOs3aSI3o6t3uK2sR5RnNqwQW082Y
cBm7zJHmmHUfwr9VLwpCOUcF5wiblpciaQFqZ8bxMgxGdUqWcChfyMuCF5XewvzK
AK1wN32u/NvzbSK3p2t3oCj08T+3b81cA0nYXUgHI4gqZA7PzrN5zYcDnoErnzKG
khLLuVBN+GFwEzNn1/97sNNCKv6TEtGmhJ+VWNnF+lhnPhpPeq+JAdKw193vZlnr
m224LUQXJ3XPq2wEQYZ2kNfmqnJ5NH8MnaQYkdGVv4kbkZi28rt8Hez0IMVWr7j3
To2QOM8cpmo5xARXV0pp1LH21xBc3oGR67Roos5j61so0HVKRsbksMGNGku7JjJh
E/TLr9Br+bYGWZ3e4K4yO2f2cS2WTJrA9FL16xfm92iXj1fbPFSZswHQ5rSArBK1
SwBBUrZrgzFsmDimxHpR60NPbiKeEur7kQ/hWO4Uc4MUmxNHV289q03xmdzFOHOn
ZP3lnw+oQsqS0cqyH7XUQ8ElEkIDzJr1A8Rif/93Ki4v3QbZ7RF1crRXfTajt12+
lvRn5MIQzMyzAeomKuK3lebZjF9Pc3GxkFziCWDYSJF+nf7eLA3+KqdUx5ofY/+w
gU2IjJuZ9DdwfJrSTo9n6AWYdPeJP0FJ/4wXruw9GBvixnRIaPoAbHJA1hV8JHAw
72/jO+IPHnKCk9pMtqFxi5RRU+WiHCuNv/in4F6sYne9TC3Kt7Mom31Y46IcnQh0
PyccAcip67Oj/sSkC52F3F7RHk24fftrFLvu31W1MTv2R9T1Y9x2IW+zHfCZHnY5
wj4sKZjkTX9ukUMeKB0/9C2bHxMOw2C5OI4TC6h33mmQvCUKpuM1GdXgl4StOYRB
kkDWcXcfH9Grp8Dgq7SkOcqRR4mcub0rx45ZlwKWXOBQMVMJuQ/lwf3tcyyiyP8K
FcUyx5JWpJU22GgHKtghI3zeV0tsZYFSmoTiX4w5ukaY1frvUHAk5Q9Kjn2uiUWo
u7mt0/ghD6ok4/bafhpxXFmphr765PLB5/a2yvpoiYv61b4btMD2fLMWU043elVr
Qyq/6pD0WBRyPk5MoyYQuFQ3jGNJ2h9IIJVYXd+U6uyVqgnQa89xaRzFUd7j3Mpq
ZcUHCBllytJEwFHf019v16gebt/gBwvzVwDMotRHyXu6Ynz1gYvn8CwSt0vqFdl+
1kt6X7mB1n3yjR1zNKeT9kw+fzfvDhNp029C5uwIbOqPNChvprdy69LDl2tQQod6
EiBdeuNsr8D0dQF9Ssmio2Yf4HZ2egyZrSOQshelbOx5uJLxRk2+6ZPnzUhUGzyn
DCp2u4/IFVVzmd81+KJjzLBvA6/fF7rTJc0zyZpJy5PecQbcCYA1VXQFikb+VPG9
NcxA0JwKyX5IBkEwmI56Y7d0XauRvdNcnRGv+tpdNXww2i7BpymQz6zk3csfI3ve
BLDniDkoJ8/6AvHyhdFUxb3b7Ul3xWe+6mKPZgKTIsFUp0cb+RL7slngkt6/cDTx
EanQlNOx0jFePVSz2sY1DfDprKRvEaeGke4OaiGCuVBlqW1jIO7KKLeLMFg+CkCm
rj5R6s0DPy5BQsWSL6MIMgsXHB0LTHEhSEs0Dr3ZsFjoUFQ3yjpvQh2xVdhqv2CL
gaso0caNqBoXFZPWGgeGcZk4miyo5ziOUy2QeOI3FoXWhG6MbRocT+zJ0yGNj8cF
In77WQX4A/tBioi44mzLhc/r5Ew2sKE4Dj4tSyH4NmgmcPYB6/TnRPKJ3VZBzVQ2
wKU3hycxbJuFzB2IMp+Y4Dm95GlJUomj48s/TIBR9KjbXqEg7HZpkLFIq03B2Jrx
tP1AVGGk5lYQriLNItjf2GvbQDPcRqV0ZGtPBt8tMLSL1rjdWVqR8TKBn6BrVN4S
U3XbXEEUvFyJ7uh8rE4pz5oy4Uq0NNYJzR3snrfiu+OXkpDsJnQnjOEDsIAj5q2r
U1sBUg8Ut+PCMbI7R5tMyNArsVKm2nRZPuy33qKwxQ/FfpBvC+edZXw1uzXLxfUF
cnKhESvS0zqG9PRGKE7dLJv5F60Utzbn1jLrMtsgKhyMMZW6CI3UhwQeeFkgrt3P
klnitZuY5ZTim5Ia9Yc1mZ42/K5fo1XYmS50B3ndYl8S3b6eW6lmkrFl22VsqOND
oj1SIjKCSmnK6Q6IqqVGC+ZvgJYnuejXdyhhQjxHkgQWQiX/ro+ZOcFspGYJDxMd
ztene/qmK1virwlpy/EsXWqZqL0o6PF14p3mPoa7T5QYUtqqj9rHSyMT4sTcyacX
OOAV8lzZST+bTDbaLzMsMV9k4hSmvKi/JVQ1jJ+HtrOWT45oxwg35K+3BOaodbzJ
wC8WMYjVPB5GsrB4Tbrqrc+yfvyzsiK+hYBJBJ6oCkh/HAhZ2vFMGuBBzF3rx+A5
Cx9DH6PtOecfj9MuNFXa2QqzauY31/ZAMrqWPaNmCIE1e4DkwOCiAuuLcg9CUcj9
2sJi2uc8/41c+rJ4ZCx4+eU5PWiZbu9KEaTi0lbUT9ditMXXuhKLDE9Mkf9ojdrn
GHudQ2ZWiMPrwh1+WwZrFIk7aIgEGvUtr6t3S+GangPcQSSie2+CrH4WaKBusUZv
OCnjGUViDixXb23k6ITOX+/rjWM/+6K3Yj5Il+hNt3c2nkH9d2pB7Z3EIdZBJ3QA
+ryFiYGHzRgA4Oynr5PhQHGDKA7khDVckL2ytlFHF/qAdusQhyWm+bsYwWQWsf6N
nQZ8mm2Euy0WNOvbuLsnQrO4f36xGY8YzJ7f5dHi7uiX6pVxyb32WiH+YL7l0RvL
6CiKybvmhTPB/ILm5mV9QSaDf/mYt7/hcva6937pe3/1Zxs8q+UunEZTlHB4LRvH
OW8EocmhtY88m4ntpD7IH8Wy7C6SWWyIkl4I7vCjphejrYdo60XJOzy8uicCJchs
9LtsnL2kdSOcF4/eIDXifafjY5rcf6U4X1QTUHCvmJljZp42PP/bQg2wyYw8CDng
ljO8rUZh1qEOa43B6x8LwcwzUxl7u2E5UuRIJ1XB8VQpHtRUYiIE2vKk4LUAvdPS
98bCxdjq7BkFCAmsOXJmv98bPD7laGX4whzrcoJSmdAgJklqJ/jbffM+K5FKnAwW
MzTht85WcmTP2rs+9kHPfAPPLh0QYCM1+w6+jClmNz44G/zW7KPKCQ4wusOxk7gM
tHCBAWM6ebc5rDjtjwnJYTtFKjDjwzu0gj+WTyRXi5ANbybtEgPo0uYos0BJdUjK
0TRvsKyiTHNJ+u9E5ZOXdQhDAHfNBR7XbJ9g/yHM7vUX8SxQMKkttSz7RDq+CaTH
WN6aVTTaMOSZU5Bhq4VBFjz6QJMiNSNx1UIHUbNN2u3LH1mbM/wa3yV4Oufdvgiz
BJ50425rS7t4MaRsuNS7ALmDwf6NoY+nFyKPb344I2lyYZuBZNIEhC0nm1FMxe0u
7sovpi56wQp9pfjrmH7153dAorAQE5x3xfQ6jJaOIwcFV3o+Vhw6cKZzH0Ozr3N5
rkzQ9YmXboWmp3wZtM528oeD+Lfcs0mytcT9N2w5+dlpI+14udIvB8k3FSk8XN3f
uObFN2X5ihWwacI6wwyNIKaLs4KH42ii7bWQNgCpZE1Km2XJMQQZIdXQ2Emr+jow
AH/cyow8QxqQ7SNpNf2MAAQEp+ZLLvBuN5SRfVBcO5YiuubfK/lmshssZUeT3qyF
VWg1bPA4HUlSXt2Ft5Ngv9QKIGeGZF2poQHxWeQwvK1282u7bayYJbUEU5Sv7Ziq
VfuXj9+KCHJC71uRVTcfDVsxmLyXoiWlg5NexqbX5F7DbadTCDMj/x7kNbYFttOl
TCq4u0diHmlMBJut+V9h9IJoeYF/poCXtp/ZH0C88ri+bdXnbyy1RXF5tkHUOj+V
3je+ACp8ibbcBu7Ig2vT1NUBtz4Ep4gLVFp55RqOsRZ4VaWYwSjCutkg69p+Q3ds
9g0GRRUwnErWgy6rRaUuBI9SEosvZOFDwGnR/3F/gyTssS1dti7+4U8i1BWiSv3k
YmFVxbFjDloukhIstaOCkw2pSi4bVMqn0SXQeNjIKdCXeIt9KEd2AZwbtmF+Kjnp
/ObtUqMrcCLvuB1n2z18NDnrpWHAI026M0OlRQAWexrmtLny+ielnAo11iV1K9DY
i/T8ZJEBUg+p7lZ9P1moQNsIuLNQgnHeAeFikywH713LMbRK+628zke8Mt3FCET5
PVI0lu+c6pTw7CVDS3hEwcI3Sobia/PpN8nLC0vGnVmzUG7LzTlh3RXx5vn65KgN
SwiUhfEuH9HANwBb6AgFcPYaJ3Xcprer3CglY7+vFkrKf0H0k4yGbOjcPKITHIXk
rgkT6gdbaTcoNZEPgOKbjjEKvk4G2cxHZy+nuoNFRQAPyIXlAfZfcKqhwawWzeUW
tajLal+v/3fbPHHwP5vkJ+MiYjAsv636JyOH27J11HrUilLXJWlilS+0ZfuQHEH1
gyLFvZCOZq4wIyBdoPuxKzz9ktzdFjdcpWRhgODc6U7o0gJx4KXzL+OCKjOISkEC
d0n8KQe19NtJv22WO4TimlEaG39NxUDHe4CdylumDJ6ZwD4QSSTxJ3Ng2c0tPuPO
0xC6g7KxlmfbN3QfSpbzOL2F2sMvbq1iKFX32/jKUDsItDPWYoxw50HOajBo4LEM
j63JhoifmGmcNxW9P5eBzwx10PUcQlZxvUtE+61HhXZJClaXNqmr4D7g9OGz0DJs
RvRRXBKhdD6B+YLpjuC/S5cjn11vbLvOtv8g2o0gD7W137AeOAigkQHPsLLwQy4x
wZb1rqS6rb7MK25tDe6pd4OQXtf1Pq+0WxtaKBJ42Z73Ily5We/ldxtl0UZbRYmM
0ipr4ffNcsaUaXcQ0ZO00GVcf3lINZ+qIUCQJpd73NtnwIXjpjXE4MTpawSnz4kq
fvptZpuzywDeOsTzr+CX+tat7v8yD2xYsriTnX2QaDqezCY4NmxTzAzKgI58Z8Dr
hpvsCMHfLpXRdVcNS8JPqhJ2YuVR3y9PTlHYj7MS5s8YGoR6vOZcRl/XxJt06WGh
pHvImqhy8ftNw5WY4SY58adXyOwtqP2PiERY6poIU9XJxd+j/edqD8qJ+px0XsmG
UNJYvSsIsCbqeOs5flp+zHcFnMLX/KOpj8Ml3lzBsHPbVcK680JT1LU3lKQhFYZw
xnLgCIZJr4FXmRMuhEbGIbt/zoC1zBluADWp3in1c6Vt5GAbFUXWv3ZUWp0eKHBp
mdHNZV5+6Ptdaq7t0suZqh/PMMf5cuF1qyZ2qP11DJpyJf7TvqkTlgLE6mDeNV0s
gqml3ucyDxSwQ6Fr5eKne8XRXGo0s5gYoLtCHFSQah8BYXVsL5ohcceTYTz/rgM9
X8O7EOyMOTbCKigpB694WV18EVLYdgfSdOwlBknoCoMnX8SAaE8xoK52FuDjQehL
hGIED6kfsHkR8XUipB8Aserq2bNx1qWafqXNmfogcTiP1tCrPGrimi5XTqZAYZua
zMtwgGP1bi7+M9/9ilTfjvdCK4+wqK2awQhulSuXFptyqL5BsgUQagOI/khnFjF4
kyEG0E1pctku9D7gpHD9GXagwKDlPh4ZU4xlFv6bGvBZstvus6daXSefHcLDx3Fv
GyTfuwIve21hzbu1sTlnAJhJ39XnESuBvexxwFrcX+4uC+E50Po58jCFKWSjNpq+
RbbpEKN/MyWUGBr5IgWlRt4MoHJwMvWWJz5KklebcpW6gTxfAisMgN0IKuS4sWvU
xUm5yvwOSsfJWxGKBsCvwviGr9k65HudXRWskxGCoz+qr/7D+Yw0yH3qTtpE6l4g
HBw+44aVCdNYiEErx8FPRjMUgtfqmVmeqkTjqqWPToWQ0myAgjf1xiKS2htYAjV6
Xj1Y+Fyhsl6pPVWylM2VifZlr7CCoFgXKM0fUKLmPoMG00peKl+utIvrMsfQeJzZ
T7dRQQGgA3wAivKtoqBFImKNepgivhzo/J+RE752AZWXjpqjaHyWFDaP0jFYJUh5
XLpohqZIe7LIlwpyQvumV7zZLVxtWK+/sV4Kmhke+1D8YCsuhNh1mjT1E4tu+9xv
jD+o1vb7XxTQ5sTtOXPnUo9DBij+lL8ZjE+ZJm//JzUKEAMn9bqopzKSebAyyMSn
GdoD4G6LIR/nI3/q2vLSPbXwjgyHhZqQSAKcioxFP5IUJCAaCzQBKsyAX12F0in3
DrXfWSYNDUBrgteJbg0dJGWTWRgm87AEZ0jxLKHyqn1QFQyag6wVbMAkT3nV+W+n
hcuVXZgyIZXIXgIuXgyLksGJDPdQFgXEDIZr5neM2ttBpx16kn+ENxn5ZHpSpy+I
9wa1D1PyTezK3I0FFL3yR4WW3oKRoULGYnHENtMzrFsGdVfAjuvcFd4QNFDuPNhH
NsV5dPc0SHSUc0R7+P/unK8Eby/yjLRrFVjhBKtawhXRTb8Q529FuVvCcG6Cg4Dn
4swGNJGB7jjjtz9TXvixHfq7ym3f5ffN5g472Tejje6TODZ++4NZyJDdcCFBlp6B
PpeRfwX92x8f8n542xoIfqF5fLIuJxVXZZfwtcXgnLNNeyESfYCMKoBKjROXdXRi
RD83W7Udt1lMg9WLTfjpIrnck6WInpzFA0/v6wGx/5qt8t6qDhQA/a+OdqnSFanz
CZ45y7bQnSqJi5725DlVc6b/EygK3jkDgQZQowFI7gseoQUTk5+Hw09UdM3tq1FL
0ofPvq2QzRJhZfgWxYndJQILDSSH5A/1IEdK5Q0aiLCrs9wgK31Vdl5XhNz5dmRX
gBeoYDhoKBCu4k5PxMPCZnMUK38aYkqSAIZkZRV28tFgtxhvDgao0UH64COKVi/9
ehEMDjkv9DOQz9X9xOwaIqTmqp/YMg8dYNNnuofCBJaWnfaVvlJKmVqmlrdk0oCy
9VD5Rpn9to5b9y6bmmGKXipgU+Bia6Ay6/ulVx9YUnVV7FuTp84Y4NI9Kz1MV/0T
Zc0nDxAFwr63Wnq9rkpePzOcRZoUScbQ/l9YZ8Z1p3KXVgbnHu4NQbMg9W0RWn6V
HDgDZc/+zaGSa8lOFU8aiZA/tOh3bbRcLlP/pYsMnAfK4AnE5UF1LPVF0AFmqm3V
takAvYjbXgyxa+3YVi6v4LVLqQyT7St5iN8MgMV1K/MY4yFlba8klM2ZyM0QDJeN
V0RnHDZYnSvH+9SH3JqU/9OCkeoRUzEe0VkjGJG6Y5WkgibOlxN+l9BVOYj8cEd7
SXd6dnUJNObQdnMs/jnNgx9JNLaoaZPn+kaGfx0367wHgrZrdpHRu5tNrA68zrSg
Kgg0wuXDQct+18x/CJFJZ7YiC4epTwtjKQv64mtqdzxSQ5IAHjY6sSz2E0xKGxir
hRAJsl7LEyLruIsFveauuoGC/ykldXD86Jl5L2ZluoQRkgbu37t2TJAM3GT+8KsM
AceNmvq5eOM5mnmZ1HxSnM6Uga9TPDHVvD+p+DMuWcwRWYq7LQzmXXYHjxVf8U+W
r+AqwyFnOjJyPDI4ldkvDXhuStyWXCIwPiXjGLkoL3Qxq087it3Mw1906VStNyW4
W70plleNpuXLL8VA6SG243qSwTOfyjOANQC1HvCZWAeHqiUWJuH9PzGZcc/UYrNN
rdievyE1uabLMUin0nWDF1AwfyFJbe9WRujBRpLGHKMlcsLfyNsZm4zGN/Tz+b2+
QmPPmbHY5taif530m7wJ8/1VwMh6iM6N3JZcItKNGnwIHHSYDUa/ZArBQVPtg++G
21Z9ZoWklsh3nnlGbmgwZPcr+vkc5kPjCbH5qFuBj7PY2G9UZWGq/eO68xHRSYMB
Tt7HbcJ1fwZfzGAD2fIqxLc6/9HenwglzfgR4z4v/xq8NAogtMnjGr6cRlaP65AB
gSvXwNURqlyehbYtdqZZrjdAkbY0w7m1FGg9792MUQKooRUV7CcgsUOUo0JG8B69
TvRaYfjYrZNODYF2bP/nK5m65nvkewCFr8zIEhqziQ4rnRhKB47Mf0W/8YPUIG8E
jxnwgucbZRf+DRKHi3wWkDFPZEjJVTePAMWUveBxR+1jQHjEexZmFLMyYpa2K2Iv
WsF9sSwZyvEX0OObxvlycsU3OnhkWJ+IDFC3cot7Hy2DIaDaR1nof9skIcMagCWc
2m1FAmwy2+tzQgHKf7Rtd8qHz2mcQrQDMUIRK5+KAlmE85X1zEsPSo/T2jmiUAlK
sK3OsnPBBLv+E2kiINaCkrjl4PBjGeC8J1Z5K3O9NIp6R8D4vH0VUSvtJiYZ1S4z
HJYLWMjCVpL79AX1BN1Trz/Nup5afhg0HQZ1RTP/1kgo4erD6YF8huDn3xXBSOS1
de3qVE+r0DbkmyUOyiTE6316S9xGz7/jqKSyniskQfNUIFH8kGgtcldC8qs8nwUe
t8fRwThrReZCsVed2oevdXcPvEykO/5rRfNgZdCP3zTtrWMMhhlZrkvc7zZtQMbb
eISFWpJxJc/P9rXzGlM366pgf/mWVEJPLJz8RwOT0Bu3s5Xf73qEIpDXFyla/tFR
E4gXwmjPddRwKzZ3HeMWHYDsT4+b9xEsjn06CYVLvUI498nPS3993G4K6SFOO0oV
GdMk5uP9mFJ/pb5bsfrSrha0KngUS+zOOo5UHE8FNed5c5omTg/hX5C030uDY+A7
bRrbeNWIcdSea8O3/0VYB59u49vP4OuH65fD2e8++ax4EDWC+a/KrFRjqnzzw/xm
jMGzcJfJrT6zpRVGBu70KbOvqOEpoEo3qZhf4DzgNFxybFaeWxh6GXE/Uk20IBNL
b5NvyHZ0atXV2HnABFNI9eynBpXrRrDDECfSdTRICIb6twgxs1zYPPXBI/dmCzO9
TTHw9M4b7RnGAdw9X3v2zCcqtpNcPuW+j4DSWcAVTB/aDZZw9P55E7byKq6PqsjO
xYMWucR4V8xC6UFJk9WoEEX4+PSJ65nYHcscuscp5qoU6Qjkdd3wD1/ycrvTsVSp
sfCujaItXPlyUBfNTLJQU2ZlbQ3kcS67XZFxJ1122J2ZplC7dRnvJInKvikE3F2o
YSF9jq2WjDjlNBkBPAhhT9WwLawgZJGC8XxlWenAUaMNS5B9CRG+PmfVslfD5QG1
w53jb+t16OKnSVYaI4DddpBsRB3m8UVdvHwvSM495ZR63lxu/0SM1hkmQ/7d8g1P
3H6KSyFu/xdl5QH+piXdDITXl7fYHcl0glnqasXCp2/SLy5dLFZs2kBtT/cD1Ms9
5j99kHCF241qmDxn4psBqR1BYUsLPqXAiRJKn2tktOriZ7c/y9DLWeeFoyPnLdM6
oniHbwmGTUGv+wXdFxfHt7k/l7PPkG/xGzB9g39iAS6N3YQINMnG7KqeV60O2D4s
3cca23Np+aeXxHqJZaPlKMr4+s804fpciIW6swKUTtjt+NpOH0PR7oKKZ7HV55EC
DdytNcBv47PNr6oo5lEIxt2A48u9uwnaG9nyZkWOM2M72sOL+GaOsj7oSyLVd/JJ
q6oUZ79hNv2Xe7ZzCXCgZDH+Ron/hf3yzDF1k2snjxg5CVsN9qul6kBOBrUNAEeT
XKr/6mXMd7CXjz5IYpFgJ15Xr6M/2V02nCDg+IsDWIR/yeocal5rgvsy1ZbIjoLb
m1LbSm607cScv1Z/aL07eHD1z21IlT5LwkP7hwHjG2DziFWopXpAjaMcGWD6l+Ck
zPluVZ73gs51okozFxkrWqEzmYVPvJ2ayZVGBDxfoOkpVNcYXcJlF2jLdw328RYQ
VG7SWhzc+oZ+F1x3u7aSYVjPB3aYG6oMvYsNxrRUBv8uv/BYA13RKUC+QkzSccGS
DutH/Bf2TCXLL6jgqU1wqMEl2zpmuNR/y9sH7rTRK5ORg9JzAez2dVooIpbzhcDh
bJaRLbjmSs2LZS67Mn0JEJuestZ0RNeMe3VK59HG0v6i0+eexdfggUbOahkD7US+
zMnnNCqo2CUYcoFW8rDg1dA3WX2Dw+HOeOMwwCOhT9H6dNOt4vLz8EICcJ8DYdZ9
TmcyhoUycdctlAGicljY7mCrKcsyz2jTX7gGiYr0jGda4rEwo8g33x/zvoRe9yAh
QtIhHvprR4E9hRa3UoPt0pId6UCESnk4kd0R9j1932+FRigp1g72So7XaX1lXWM3
UNc04oMX3a4NxsT+iLzVklx8gTPSp9WRJU3t8EHJ4StCHBIhaeckrst50hUPUsfT
Dx3f87f/SsrHnBXwTPLfx5vo2bohRa+mpRT//5EZLJkt6//xAybMwuXWXpLsW/Ip
dVKLrZH5BB/yMTuSLCuEemqqXwPBTb+Lts7Lr6tlG7Oo+Cr31k0wKMRBTWsuahmu
1hrJsKFqF6jC85PtKqrnVPIr9VZtd6mp8SV0fmbY13fcU9kbOB5XW6ire+AaOyWX
RnGv7hzo+6dw9vVWNT6P/oYmXCokXvN+TvQQsAAdG/m8x2aA0ScTR3gCdnNeFiSG
nrv453rQV0FEolR6SBdSHZPvanayx3psNlgDRSU5YuYwWDYV/kFMkw3Jtx3mAOWz
Dkb6MeCh6TqfoX8/lde+W+7ZWZXRqWr2I9MvbNmrgV/fe5nvOIPW+vDoCL+oAVA7
s/qz2UnA+Y7oxUVXxuBBn9RHIVMrH4N6/MY2UcdHAdgFXx6KTkpt5ahu1gTaVWlK
tSETFEbRWjtIncRdPJoKMWjfM4s6JUpV4mHKJbc1qtQQjgsH7RGPnvXGVZxn58lR
bLPyEWpW7g3PcO/H9aeyXTI01hdO8UhKUH1+4QePp5A/2gRfVbsRRuff+F0JKIhO
fwt00GueDuGnmYfnmfDMXFreqoC8mAhTMxJ2uSpw7VFXUOR3d7RVAwCLvVoDrhWN
c+KbhhjDXe6LcBBOo+xyi9G7mBU4D7nIxyQz07FaAtrlfnQkh1eWZI1rnEcs2Upj
fxkNYaLQK6Eq7IJLgPLULK+6gVMFHAf4hiMK2W3+gnbZNU+t36TQRTlYnM089U0P
XuEJkk2aqPEoqpZ4wUP80vKv7U5BPXkPNa+OTUYcaP6IvLf803GvegJNX+rWSPmR
B2B3lH/S3CVAJSNKNb3s5qSUa+HAEbpGfJpS97Eb4ijufjTO/umywm3BiiWT58F+
+UPyHtVSt4pXZ1EkcvY+aXQ3fxFXkg7VVTycISCWxikvfczTNmKawbVPWy+WIO9y
y7FY1Dp45UF52SbSDvhD9J/RXY0VRt7fyuxUfMClNpGVPdUorvTPc635TDJ/pGu0
7VkzeOZe3xg3gy7D4jYkwMLk0CaGR7vK5uNiBXqSjuqoG7Jb7ZYuBBTXi443cZ+7
e1zAVrqFaBjTk5LTxyJdK2Vsc+lV2T8GKrDWWXELv9njLMy+Vah/VQ+ae49LxAMr
lCJ5oZ38kOqnFdaTIyKTExuI2sIWFsOsI7Vsi3WuTo+9fdjoLhvhdoniWr7+hx53
RGrp0HoPmhLsd6DPUn/KjACxDH5loaRknZbn2any3Nl2vvFPCTqG2wQAqI0obb1E
TXmJoX+pJXkGt7w77G1mqIfkN8ElqRnDe/3lcXg2ad9g/QN0jvmZjgS9RuRvi2Jj
3tu/zqlqxGXATysLeb1G+8Je9O9KROpQwlfbq+Avlx+8zan1oQqqKOrsl4da2kvX
15N9NjLFsb4YTX0NWWbk4ORaEDfsTxEgyDZrg8NLaiTmWrtXLvmOmWEiv7ywXRcx
3qhze8oIZwF52z0zpIVLSHNgERRMhQ8VEf4NEo4+o0pgk0pW4PxJOJXog1F6OwEo
HGmoQVfSee98VMDfy9Z6G7f74m7hJmkRSrCz+yY+k9j88FyWnI60i0oOgOekaIVR
CcZHrxi27nHT6tVFWpC6jvQUF1L89+i1Rg/L6Ek2GnTOJmY65SHIFIJ9wnGAUTbc
VCSmjRtuJUpNg+9PKFqzEGXWFvnIqmKvemHdzzXkZ2kY+FIaQminz3DOrnN0Riej
2bPqflnaHJhBTAF+YSNEq/qi+nMLt1sN6KSZfeJ1a/N8nwEd2qgSA3M95YF4ICUk
aXcF5vFxN/odHMiPzbzpa6GuNoXs/txWfN+9jcYDsM87QNyzwWK/iLW+bO+WleUp
e4gW2k3FETg7BUmJKvXeluK+gHdA723PKyQZxh82s+XslDcbxGL4iROidaiq0itz
ZskfqPK6u90JGyfgJqEhrXMPRmoEPiLINHn0DcJdBLgMfRB9mW0P42/MxEuYp8zY
0WgclbpxdE8io0jEXxsobPyPobiHlXJVM+BxfXsojJm2pRpqUvqna0LP2I5WEq04
4uu3E0ivNngA3T/wiEUfbovtoGG7F1QHwk0mJZnKBGl1pZkC2ALesNvV25ovbPkO
ZdBbzknjoa0uKkQBFWSy4jTSOg0MJ/qBwkxAEb+5fKN2pmd4FjW3v2uGK5xsYwIo
OeL/AeAn/dE8i4o0zgsXHbbHmF091ebB35TuHA8neZq3r3H8w4AMly8P+eeZJRHY
axLh8HFwnYq+JS8pmrg+ZVy9QUyPQ3A0jWylqvRdQTn2pEWFRFL/X6Pjx6438xRv
emB726o6+iRXbNbvnS9LdR4dsqFagbCdK8bXgYlgtGzy7dbkyK2jOcsKHXU/JhkS
yEIdOsCph/bv5xiKMifD5izJGaBHACqhKV44ezd85NXGRpF80YMDwO5+9wXhDcz5
3HJIZjlMVXuONDF+/n/9UcR3pTJ74fAPgmAnYinpjOMjSUxJCHOd9MGFL2LUSf7H
Q85p57ZpiePD/FvAgHX5QCbXFgbryBbVPaYcz4PIoSouxnDjMmA2V9OUNKETaavj
g0MHIs6hFQ2nNfLmyNEcq+ONBglmLvl/WwkbepyTObeweMCtP/HHy+8IFTV9v2KQ
y6iiGO2LQRwXhJd7wl4NOWCOUJ/Vt1pUaFkH7Fh0aGsLtfBPRUCDdri31QaFbwkm
n+1qMDZSpVO3/sPUv0Cpd7I6DkSSd4+0rZMv0GjV2hnfRq3FEQt73h72+eBGMRUB
xXftqgAR53cQwh992EULOXFFIjzpdfSn3tm41ZxYObdIjaGxcaLgbC3nkwW9HZG3
d63c8llteT+gBdcmumacKszGJrXtWPYWEpBguUHCeUwwml1ehiUTAyy9GlUzzXtm
jKhO3HGyYDciPd0jw/GLR5RYpQrEp56v1O19V4UZ7kyfVYGMDuM+xJ1HWPbtN26J
4ZsjQr3I5tPNNvX4ORsKdGWzhF/riXk/S2K/4L/YkD0MJ4pp3ETTC9UlSK7aGbc1
JizNeH0l8IOnALwQ39veCX0lPcxIAsZVSD2fs4RqaTgm+LxYHYD79sGBIjdZ+Qcx
+4sr0L0Y9Ott2Oet/wL+xRqmxQ+ylBF1/K9FDOQTPIYgi6GR1/kx1Mpsn1pigABW
jvxE6f/p15aup5g/Ii3Xra8QR09QaeBQMledsCPx33Ukqxie+T2KDCWG30FAlnJ5
++uRxCiOcMuBdRh6DEMiv8KvaIBaPcIYVsF6jhndE2U4KFQjuxKdkcN6lRWoj9Pr
V5sAS3rfMPOL1OeSFnZuToLj/oPc6cx2pIyRDTuTN9v24DfCvfSxPOCzWNTwPA3z
2kcdJTMiD5QA+L+/KeEBk5Zdrk8BCYn0eQgS/gtmrMan/q+329w+OC1rsRAKW8Pq
BRbQNLzCNNohOLHoMClzuQr1uKvqY+8tr6NcTXqvgNeV9I7Cbla55gNbXxSRAcH5
UHdfXnOXcffNNL7d5Rgngs+lmNgapy2YyWrXcdZgRIwvQBw0maPO2bY/Vpi9tXAR
bbmNApKzorUNQXmfehxZU+bd0m/FD9iIsr/twYtI6CEvtr0qtmEQZ65ictXNcFgM
gaKXyv0qQ0pPoJbkJezqYNbk0oK9YOhXrKMEk31Uhm3mrSi6fDQZ+Xdz+PPDZAgs
Q6Jj/qXYUqchwCqunPcQ25Nwhb1q1CQa4JKvJOs5xIP9gzcXyrEidXXlu96Es/s3
0GK4k3/yhkvsLH7zTjoznK/u6AI6IvcLy3snOL757/27Oa1MyipWnHIoFJOEbJLN
7AXLbCR8f8yNadjMY4BNoFA75yi6E2RKf0+CnUkIvFfV3TNvJvjnFevxztdr+PRK
udaOgR0GZACH0EYwV/QYlLHkkNqIlPbv7l30fgslr5SVPAnDB9qj0En7gclKXUXH
5jSoZRlHfc5WjF9J1w1Ay2gCpONpg71wymEbSkCFRl+vTie7P1S6wzb9jyvdihEq
tY88DJZ2cI6BwbYPjx6DFGCxD1MyPROAcWNdJq3+rAfJzE4LpDykJYYCWAgQuaD2
jizYXCHdLfmYi4E55b6FuuSlHhSlh9SPpXlK5nurv02F45LTwQdYHgIBQFLcjkMq
VoXh5dO5e3nUcG4IdeefwX4PDXjX/e5TKk1jmM53PS12zimeob8I172tf2d4jZZj
3lBg1iRFJ9O+R67DhIRN7GNHunpdMtGUr1YGoYyQeZcOw6y/WFyfPLybcmxNdLVa
0y9l3Sd8lxUs4AaIi3rScC0D1YnC04AahhpAfmu3L38rSW7xy/tAWHqYE7uJ9CJ6
fH4FlW1sfrg/upBxoLewaKRGZrUEblY9l4bzF7oWcgKNFnyzj1SqYUZQxB3igD24
g/Le1r8c9HWENb/dyq0CznbRp9HvNhPdm5G02aHUHnHkLdH3dyNpiTYVFSMk0gnF
DJ1+VVM90JelWHEjA+49vCr6ThVVA3i0Vl3e3T1DlbbyiLmVsVMyTig/H+92uvFA
j8I+xkhDA+m3FSYGIZyztMnXcxSEb0T8sclwC1d650DeTnwaDCEC9QQ0pIBHAD3U
cbrkFR1csyzU6RnJNd4bkuabEfuQICQ9xjkjIiZUCcxSLsxfjjsXzPr06d0xWwJ4
Ivoz86/d6T7P+YiqXHKCo1SjL8oBWFFeEwIybByAoH8JSeF5wQRkKVaIUDzDnFGE
PfDSBaEHWwlTG7OP0byD/sYF0+YCVKDDtGUazHwOZOhJcWTOnnilU7+ooqBAs61V
F5h2GZ3F1v0Zydbm5/BgZuVQqYw7ryhTiR/UGmNitLMy+rnjeULus7zAWX55AaEh
8jK85avU9/49itNa1LLWMiAgCX4f1LVx472J861hJ/ilyo3F8uWW8zD3luqRHoPH
hahbT9UN3RDw+eVihBBHYU3Rj4OHi4i3xaX4CPakm+Qk5QoA7S7IgvsR2jfv50Xr
hMR4bFSSAq+OfRaqwzlUEqJpSng7sATdHgpTYXOvjE4cmQ1rUc95Xg+7PEAg2I3l
tRwNHWClTg56pveFLfICJV39eHTtpgMca94+Ql2tmdnPTJkmBSCMRXHTSrO+Bu9Z
kZ6SQA8Gr8ZbvUomLxO1h7qt24rlLJb88PR3IGjFBm0cQFn4FQt+X2hFiJNssFzS
VkZBlofPLfJOnz/0vYaDPuI2xFRdJ5e5XOgL7gm/jG82q+0DVQqzC+TSKVhHqXAN
LOp6h41u0RCKBlPvc5gb7bIEhY9iTlB+UnARZoKdnf9Xk256hIXR/uPm2o2Z/xLG
JJTIsz8XTBM5wThbJdcqO8vpY089bQvM4REpiZk/oDn9eEhsjQNka/k73x+IRO1g
3X3JuTkZyaaAU5MHLeCXj/MyrQueU304cztE6fENBxlofWL7dYJhz4iyzt5r3apL
MNAvBx2Frdta+lZJq51YpvYBJvOXqCRwqoYeF8oEwxsJVyYQJ6yb5gP0eENX4gGF
yIyavdiIOIJKsPTRfg64x1SoYlPyT6k/8KPGltIJ8evS3gq3OwQLOkyBP++li1CX
Zi4RNYqS1FNbFMShbGyptVrHT9b0g7HhauOTxA9+F15lgukzv4KMyclC8fJg8xLq
j++LmDMMOcC51D795/fZV2Kr2/b68HYWfTaPbtqnJTTOt46NdbLv0UdRd19CyAba
qiX6QNrqwJ3oFRnSA/0XPIbcgQiQgugFG756+GN44a5/WFBYBxaE1c3N6AzBxjSc
GoG7vHGZG+iiuHPm+TUhuBa7p/xtNe4WuPqw9th/TOiwjZU6QgWzM5b3J1Veb3uy
6Jx+M+OsX4fpObX8tBFca/RsRi9gtKdADtlohBaoOkBVqYAurxbAMTbQSUelntB+
S6aJ3HHLIUyqhn5ku+X0PZYxFh00XkQQPPQPLyh4zysEAtZx5vHhzXSaS2uJ4BOb
Pggu5Bpc4IO9eewicyT+V+5QaSWE3diKp5FzP9KVQL3aJ8NFeGyZ8Mz+v/KpeMgk
wrK7q/oDp6e2GTFnZ9rSJbLJ+qNJi8KQKNNxd18dFimc5RKeGMHMQkplQragDlGf
GsU7X1ZoISNcG328BAOG9RyyqjqJNoy20j41JcozKWXUYiQy3acktdDWc8iujYTJ
hPopKhmniDTMhUJWtOyZpTCNRsARd8PyLcnhA8Fu8TSdushu0/tfJpcL3C6dSUb/
lsUTLk0fkloo644My5e/zUuATfFeXMKzAWwojQrq7+Yt+b9OQ4xZDEMc14VJK3nP
qPlTrF8H0gVwU46uh6nlCJ+EZPEwONJ6D6dFhd+Blz2EF3g//i6RFY9d4FqmY6pT
/QzMoxAG6c+LEJ23YphTFhjmlWNJwTZf6xc1jC1uiRJGeIz4OoU24pdmQcuK5SgT
Ul+GJdlLliwETtW0rGhNCB/H1W3q2oNojSlFrRnzKWB/caJQWOneagSpSrhFOwVM
pbX1IemJtklyCkuoVa9mouw9nCpjAOqNs4dDYhWRyXJj6wwiWWf76UfuKNva4p/m
NwE03EANmL4QlBIaexQVo0UygAxEMa/uJ9mRs7Dk/mSIovvJItOwwot0KNGft5XC
O0GNlknoEOvy5rFFBsfvU7b/wGsA6H6SvCiFXlzf7xujsbRu99nuSFN8saFMz8q/
NZu/wuKVGSPkxb+e/0pp0430YiKVwH50nPpofBHEavUJemzYd9GEgFkioWvENHRt
kTDy5qV5hDmkOJd1QM/9GMfd8WXwkA6VZ65Zy1fYyMMl8FOgMGQLTmMNJ/1RA+HF
Fm6dVRjGEQ3lWg1xZ6bCCOZrn2mIbOAM4rIZj2V2nmyHngV5MWrvvEwFuuPgUUcI
GZsRrPl8vdhfXzw6OC+h1kj8YQSx5n6S35qfdVYFhS/XygqhU+ucW/WReNKJy7bM
xwjrZC2pMVzKHdceZCOfreDL+osmbzjGN8BL49rVA9WQwxZKx1Ue8KRQCIFBeahO
osCX/g55f+AKczr8fnMb5WT/lsyBqYlXMR+dBAs0vaSvr4OvZ0bYdB0Dg3rmMMK6
95r6l41jug3nSl/XUhTBwWY+UpLKAZs3MvZlgCifj8piRR4AbjqaxNQtcZ6pZNNQ
K7BbaU5GRRCz8Cdg1nvDYqATRvOOhEaLqGfHnLZY0GXYqcla0LUqoCAxjkYcI6Xd
iFG/3oxDvHW1uNwrZnCypXJMhcH4/KpBJ8gVB7vbAgfFdglgKSqX4UfxM/+/Kalf
ffRAZJgH06Ibto9PH+EGP/OuzUxisUGnTNgNap785LSworMvbN+sQPYyv/r8+kVM
TU4HDR4SL5WG3QeA44qJrlbZ0E89qhsxx5sq05T1tLWoqvJGKP5k6zfEemaXpgeC
Onv0kgk2/9yvuv6Pyldy9y3zyV4BstB57s8xzoRmQioZIIuBTfh451j0ASDLFmpb
dRI1CXfmaO9o2Amo7HcAKYXjIZrKN8QxNPsouCTczQ49UvMljUwThiYjrO0cSddO
nYCj2fLkg2PgcTjX7bpg4SBxPf+1plAVhuWPfLoIbHkUD4MazrjoR5q8QBIbWhGN
snRLwMSQ+gAb0rsiFYmOuOuMeCKROTBptXH0LnW0zOjm/RyU8l65SDTQjxQetsmf
UQXr0l9VB2IeXVWcbDf1JVgkaCL7Cc/Rkq5SmTxou56dy9x5AYiplfihk94IoEtW
ALKDP0EdAefi9+DENrqKDE/se5pHL98rE0Avz599zSZjIN+Q+DV1M+oJz+zW91V6
IePHh7OvI6A2WpKjwGY/3nOfUPUI5TH/6PoaOCOrHgbJbQ7pcpXfoKV+V6/Mdnzb
vx33uCMynVPplcmDm19gYnN78TTvg33fd0yEZ22gNmqF9OIeux0uNezZNXuBDy/T
XPoow+rcFC/3GYXxRIX0rieszJsiIxtE/47atcMrulGFGy9Ubf1EBt02VKPpde2p
Kt59pxrpcGBRpOXx9HnMLry8eliLhXak7k36SELJVbJiOTuTf2xwS+99ygTjS4By
T3YdrFq94XX+iZtc0iXeqInrfXX0SrLDsvJw2z+CDXzvssKFeOZvNnOqELOpVNny
AnoEPRUK45CkYTDK5yaUaciZ3d8ryBjmWkDm+sKuyHc5m1O//IIMI0lDbr2WB18x
6vieayLcvVx+CkQcRpFjhg1EWT08LDZyMbm/wGZeFa8CqCD/zFLPr7dnGWI/IgsD
ivYn2y5wt5eS98m2jzVMPWm2T0Qy3nlAbvt0PH1gqcG9aTbsg4Ixa2+Hd1yEbkbB
FR4lZOm3HXGL7WR1mz/5tt969WLS05pMZxLABSQZZsDuilzIHRT6K0Hkk/hsSqQ/
W9sUuRJuAH5hGhHkMHVK3o948QqOU9PedcfTuN6TA1/hlMMEvQpzWgA2ZxWD1Rhw
2NMqtnkHJz2MU/nauXKleIjaPY5lWdoRSOEN9eDZZIAgelW6uaKMP59Rq0n9Vlgn
ZQDltP4sRj2uW4ZkMZvd5Kk0wxPwVy+Y49b63DpDQNMrr9xjKWhj7HC6QGZ0HCZZ
+goKQCNaHPg+b9FZIsSiSo2HTuE2lsVA7c+rxyWx703RqfKsuejoF6RN6JzM36qC
avWDJWXN6MxpX5lUHXpF83RZrL4nYIDVL7LtssT7fvjVacsVxZSYTGy+buPObJOz
8lhd55BclD1kJB8aWI7MG5F9CwdyIYKCE5Byx2sgIMKBJdH59cAGVGMgMMehV9Wb
jzuTWi0aAP4wpMisyj03fBvxhLvrtrUTlxOcOp1YlO7jDU63tyPgFxqi0Hy4ejbk
FysbfEz3dOtlusssZtTxyPcdN/h86avzcr6vQH3xqBEIJ0tLOefU6bG0I5aB1wQR
8h4Hja4J1UTEbOYeifk0pKogRt5LtzPiCExQFaISbe7GpyzkoRISGX5y9H9OlIWX
CVb9kkFSkfGbgwRtTMTRYXfj6F9S9abzf3ZmDiMjJ69Fsjgl73uspS53nUcvvt5o
bXSoIloqFZjlrKVk2MwLRIBhPqGr6cdzCTgEWU+UKPDp0zW9PM1ZiXsv8NBFkOgk
usVM8BljJRrsyEPVzxq+rb1OuXA2VU8cMqnVfK1pCIEL6N2Yb7pK1fhODYhuLW1x
+lhkpk4pLBeCRkpfsUWRp6fu7hxtY3CVHp8TPmVyXWS5NpAnc9XOVi+ijr07VOD2
yU97BCpTmx6E/txMEXMFM5Phu88SyPKCqDdH8vVu0FT6Q5OdoVXzbH0p3M8YUJO8
YyYt/v6oc9FLUHZdSA32dtpgyfTPxfoLhYVYsj/DrNMmgKv8MaVP6cAIK8d3pY/S
UNkYOMOY1OHPXagqu7iEcsyERY3djs7fhkmDKpfuBS2JPFIJ+4qw1y4MGoJ6xNVV
ih/5HVlqPv+RXH7BPT87az7366mCfuysnXgQiFmtPTyDCvs5zm9iEhqqrmcBaRqd
JNbgeknbML+/faI/+c6VkSGTJIWElAgYiYGW32n3BanLtfK5Fa8ApaGgKXE9SL/Y
ov6EtgvGKgDlDQLCSvnHXUDUM+CT8sAWjB1cKLnC/SiLV6xJx39D9dNJ+sQ4346y
0Z877jS9t6uHUrHs3xaFPIhd7vvhPxYVIrakAp5UyxEnMjUlpxZ/zFwnds6M2Vy2
qO+zakJNzITUQMjCE9pUKG829Ahsqz6n1474PHWcHq+gW+4nFKL6U5Dguymzx56N
evGfxcOuQtHTN0s4U0XbNq33wBS3+u3cKr0qr+HR8hmVPcXGtdcTZH1BIyosForY
TF2ByXTwjKJsHCS8xucIY9Yv0dSxMX064xBXfkNHxx+D82CHzZfIgcUdf56qrNAb
kJsCT4dhlh8XOgabT7znapb+K0ryW6hBBDELhQ/9fzTuEz9U3cNR+2jaCbNxKMHM
e++auNc10PU5SxQVkwoqnub5zT8l8oskMV+ITMoUx5PxWKb9F0ekKDBPaFBGxPrw
jFJ0xk+aPOP4n9hxOIa+s646nAQuKtVxkmY0mU/wNcBeL5Ykg2C4dPSRsD3CMBP5
+EIEATzZryz69vAWnDMnnQD4JLyIYGbspn05YpR6xzgQsC7YMOvSzFg5mM14SPky
S52cj52ivW25isAnuF057TIsSJVcXeja6fsOpHKEvsWNJorlLwyEIZ22lH34dLSc
lY6jLYwO6WyJLKqHm4JE7Ti+ub6OIgZKLzqXLDrnFad+dPmCe28IqEr6iHf0o6N5
se0Jzfr3yrZ9frr2KmEcSH/cUJTXugfJt/Dh7+kgPxEAwhZd3X1dtSxjAVKSGsPl
NDDQ3NFcbVkCTWOQAh7kuDMvNRR87hSveOp/iPU0hIZgjQyVA3aA9ljfJ86KEBnX
XUTH1rYO3dmfhzA0pcKyS5BPjM5G1pi+hnZmPWMWR4FUALUGd6rWkFh1qCJrTFMB
W7n6d+VqTLLmOPuriAFbFZkrjULXgV7txiVpvF6iBETNp3WtxS/w7e8rIo3jJv1g
oWLa/MV2bAtBOnH/JB7B+Udl3ue6QGN+RdMuxh7DfEHmd1+b0zGwbaREhmquspzx
0HkSb0D0u3CRXLE0gqj8ZNq4pUJ7e2p7kZ630O6MIe4HJUbr74QpkHXDsyXglJE1
CHL9IJpIYsYqBcGJ08g2VTiD4xeabgRg2CtQyvJF+jpZT4VmB9lZzSRv5Gsdr53e
2gBfy/y+FYNb+TryOVaXBbVSMSeXOHZZYrVQl5YEV2tJrlA3sCXIiZn5RODf2rgj
muSBkykK6IP8YJ3leoeusjp1NC75nD0RZxkVFMSXbxPqI+pI0tia36y5Qox1N+7P
80LvcUSKZngqH3ewK3mQJarlQCR5JScRnqEJ9X7GNVVmAb4LkjZ7CTIQ8aFML39s
rdL9TTcsLeb8n9LCtkTmgJOpfnKQnN6yDOWNYHrHiZ/qK1rrak67D4DNaQd77VVP
pokyOM3TZZOY4TtAuAtJIO691RjOxLsdVQGPHnDAnGMc89yN32yC4c1E8vkdksJT
oaEOQCneWhNOxeAhzPVJyt6EmKHOvaKqLbhdDTpvvaKnhoYiyeqsjkzPY1SoNeeX
aYtKP9yNMOJt6end3AK/zGRnpxfCu4Ct3EQwOh5CNWt9o+BfAR26z9CIRIkttKBV
1nq2XsrmH5qe9bviuR1XJeHKP28pOiIywclg0ugE6UYZCIpiStKIHLgSEZEsOA/E
1TJCB/iHqqgpVNjJAiFzAGi3n4MG3n4BxVz9CPEzRLzua9r6oTug57aFtOfGd0Ra
Y6Rj4Gs6hTxcbC0jxQkG/h0UsK/tNNvTx8zIRTOl4cRbZmwB8CSpja07jJx0PRwA
vBjWMH9981ekSzoBFHoAiuiK7IKn8kehzMeH42NtLgWWE+YV7yL65CXzr61xExhM
6BdZIfK3xR5csn2Sq4KDDXvvKMxIfRmSn39dJjqF8wnDvTZNneJIyuPRsOBYh66+
969JO5v82muwqGiLi9lvy6AeKLg5o7Q508+vQKH/3kI+4kXM1lvoYqgX/R94rIwx
5GPncVV9vT+e47M2qlm2BKv0WO3XvpTjX+BGf32y1fY7ILa93G8P4FYFx69QCOH0
peGRBfCMmYpRmWvqFxtdBkeu4qsfkcRBPNdYynGUXQpgPgstMPPreZlXVWg6XNw4
DXe+Zm0v3dvRP1n4E9UsRzJZuhLxdo5X9HCwhB8eZhLudIGUdNNfk/MncXLWcuV3
1hXy48K4FxoHxgLr0QfVyTq8JZhYLTeQiX04YEEhgDs0ITSejNFW9yA9kpcYGkz4
9oju4P0WiS4yVpBJDhEHbYeKNedkU+cS32B/c7SiSfQlIkmFEiMKM28U+M5U45Ji
aMqsP/DwXmpE0SeM2oMHPgGselvEV3ytmR9bJrqZsRvXnDgo+eKt47omwwGQSSTw
9TWtZ4nQiYIvtK4CL7sGG0/bjUgtRXUevbAR7hTwfKy+6kQnO/Hhz0McD0hnhOqG
J/ADoUUyX2ljcQNaFBcFocqxtMRLRmsZeAie1QRNfku59DoL5OsTkOfR2HdQEUm/
Z+SumbD0+/m782/HX7yoW+LTm+7JFIQxLvordEuLa1KnLut/hO/RXZwFmQJtmBfF
0AfqPv24GQjk90JcdnmROPK8d51RqUoEHd95+2JQbaWQvW4BYFedZsKFkkd+GH4+
WAFS144SHmeafN6Y+vnL8m7iUGPVOizEP4v8MecKCOZwME+6VxIqm8QSVAK1BmwB
Xz/j+I7zTgyELdpZHWP5h6k0pv7okk6Qvn0xvRCXRvZnUlseRcj9b0WwVt7doEUC
TlRj/V90+oJ2jQqyhOOYJuCpaYqYPBmkYk+atXVMk9J14DEumaRN2nARYV+XofKz
+1DJhUhVfwgFg6AU73Y+WBZQVILHCpVxn0+3IIEijtgDAmeTIILz9lt5+hXqTtJ1
0wTDjjZRb01I0rLbuiVWY/tNH+SlGJyt1vlCkKL1ikiMYCZzwoO5sgUrrcvhO4Db
1+wYXCE7AiDOBjgQkiVL4utpWZFXXw0zqn2MuTWXYkHnXXWx7V5K0RJgPR3VBa1I
rvgTWJjNwC74qlJ9dFIFpQwkQ6OwB+tkeXW3lEG52wXxvlCS8B3qZ8LCwmxU7aW3
Z5/vsnFSksdKtv+yrb6UPCClfHJEcTG1MXgq64lSjZaDApbencYon2/+5jZTZCwA
6poOdoZV0B1iraom++HH9yRjPPUH05zS3h6f3ofbzEWJKSoRsGL4NtOPKzwU1N4G
cVCmbr+WIgbpT1sVkduIa25qctqM1soxUBLGPQJFQxT2GVBQaWWALTvAHWwDOyko
GUU+8eoUqIgkLXK4Mj452CDOwxzM+qwcZA1zVqk9blvkOpSqRnlJIMHh1rfTN5Lm
kGaymJBufcbpjZq8jzOOE9+Ed9NlWVgQ/5uS6L8K6dy2eyo+bbON4RTphlTvi25y
u8snbuhC9nP7K46u8bfCIRSmvvivW3/z19ZYYPXHeY0n5pxgHKNr2nuNxmWVjFlz
W9YZpuTgBHpsV25GplAN87L9fBEPu83lT2zk7hRRxtvlhlnli7LWLx+yw8YlWFdo
vE3kylFB0bq/o/jdIs963UhUzZm+ff78GUNXmGwA562A1M6qobzXhI9nTUdPFF7H
mZY0LWAJLTk1Gbx9SEUnUpR/CgaKufiaZc7RZY8eL40AwKpoEZ/ZdCabreFRjuHj
ZLGok+80JMiirrs/A2JKGMKhKe5u0T/6DLmp7hWXeDx/qlrg3xgEC8HIhd0h7h06
CDNGGtB69rLCskDwWLTadL7jnOPvUhxPdT3N8xGifFBdqzWsQ+hdaIvFXyR3HfnX
x1CnhMWa6Jt30QdGnYMIWkSlUpG2C95/E1hraKpx+DHUbSWXm4I0UU1s5qCo8ysQ
dyoaz1p3eFA0fI3XJC4QpI5Rofbpu3rymH29sUQjJjcTCRx95+GAjOJFg79t28Bo
8cPEy87QqFeHAT/oz/R9fV2zkh5zeooOgE0bRSoASb47+dON2OramG+/qq9CMECx
njD0Ls+BfXhlfTnAFA8qnvn6GHwtAx83AiZ7TzusJQXq/vZqp/fZFNqDH3KWXfbd
u2gZ/RrGZpYOS1+lppyBtpSB3l9ZWTOSsOE0ask5vVXRp3xleuBTDM1Q5UFSWsTB
Q7IPEXJRnWF04mwayHtkTj5Z350c0YpLXlL0rflfORaA3ZDTtWBrgUa64+csTtvi
uFvQqsUsE+SWYstig5RJa+yWnWdIDT2SvYtmw89aqATZxQfsUM9szC6DFwe0ovTP
6tyE68YieaQZTWQjelvMv2WOUxFlXBbowesjg66uKPmd+GykFh3IDeSZH1MwFmad
OC0HFNdb4ew1Cqybvl0apu0HjFe3qa9RXtAfh3gWpjW90zpqCNXL0bWi7ahMhjFB
25d2QDuWyktocAfqtm4rn4EJg9uITc2DWznI2ALZbhBbuAhpKIkwSHYAI9QW+HCU
xlf0dMhHMx/3rFDfjr4jhBVMrKCZEPptiHCErHvehsL0naNI+tPnzRub3ytAk4qf
25j0075DlC7/wdS+bA70owSFoB/rWU5tpqd4gmqSKz4v+NaISf1XbqbQfc7SaY4I
ZdqwG8AMOY3oDe13KcsGPXJxeeyTh5hX5lEraRiKjaxae8KVh9hq4h7nq1PcxCdw
c9aHJIyZrxHrIpEWPlH+CHi4CS1/WohAsItLDFY+lH0N7KViidQZD2Vobt1h2Wg6
2cMGVPX8oruMiiPmDSSAwvQVlItrBatQiWxS4exYBO+dzDM+gHKYKJkbd8YmesKF
e37fJ1xgWGh94ISLhxtAP4+trcnUTr0YO4lLpb+AS/MTYeo2BN+MxNEP3dsjJ2w1
kVslzgyzLMCgPJFWJDNVdZBNcQnYNca/Qfdv+fQkErVKF0KMHgHFcWctgNr8QNFF
xP89YYhUAxfjAiZpQ6nk8TAwc618tCj6kP+Fvfgl/VrzzvhBNcCqdrEG/uz7STjN
cHrUMGXgDtJfVMs5alx6fFXrVWBVfvP4grK2zX6/8UO5bL95s8jsp6QParES+dLP
+i6vS/8oRPru3RCzrYPAufD59OG29voHc3nOXwZgyb/inxP+CMTRWVYqDGIzCzsp
3mjx++JFHgXfRXShXSo2LdxG9mulDR9mjx5HCssNiCWGgNaKcdQDLhKngAvpV0jz
mZn5j/hRYUVWWmXUA0vu8NXxSZKKIsDej0N/chKnWoZCH/xEbhFsfixT9bS3tCdr
B5B2b8EV6nsmXhD2MM0I74VocbbicTg52iHvx8LPIaPFtK9u0Owbqza0DGUeSr0M
AmFmFjZ6gBa3Hb87qqsAG6xrWunk6ZP9Bop7/Y+p6WvzAZpVzHm+aOMw9xAE/XqS
7p2EsY5V+WQLi95oN6dfqbZRFmiK/TXe2z1nPd5NahSdZbBgxvkwsMUL9VhRuz30
eCcyCjrzH1vA217a1BTVBdtzGXntqMdHYDq4g21KkRSGHmpRpaSjitOIo9oNbAs9
YC7Os1FHjzpSJpf7WDSBUF573pSSXAfX0bXGWLquDxO0gbFhpoUK917nAeXic6Mn
dngmSW/BMP3GQ/vf4O3afA8sE5Ql7nYNg6dMBSErJtEGcMNl9ajBYOZ9KsuV1xYj
mLScUORyetJ/uBHh5WVv2DsFr1Bvs0e4cTNZFf6Jb8HTsYZM9Q7rmR2+OCf8xRbS
sG1KLdEOe39Jf2y9HWnJJGvC0b43viB4UdO342aqmWZOOzJsHQ95fJ6si5DCgRW8
WP+Y4EXEi7hm7eUBQcZUr4KStYcR62ikZzOxB9zfE1sMGKSZlewElRJSzOHcWIaB
29sIwI2Gysp8bEUjTwMdFjgOwIxUtgDM59YOr66l7TjVzgbUJbeCZBNnFkkEtHEg
nj0FtdqA/lYd5vNgwWDL4mJ71+17lnsqYgDqRNTd+z8Q4C0v2ldycRF9x8WhyeY1
g2hxLbWgsjKIu7qMbcxebUNlFmvcv4sh1NkNYNOOyKC0/C+Z5xf0EP78ySn1jO/L
EisaElyA36h2b9RVU7BG6s/I7vGE7pVZ8FMcoML+h9rWyhuQUZshWFQtlADv//5d
iHmDy8DmWgIjU9AZdA0C8YHUkWrWN5C3sUurMXzDlAwiL+EcvxqFzFoF7qjSRYO0
WxYqo91i/VQwHw425BZROVwcPWVPqPFDr9FrFiyPnckd3st7IQHO1Dv0S3qhx8LK
Db3atM3MBcqYy9mS159ZmoMfUeXOLOpsybE/egP+GDgvtLmCKIQHeKwRTonNojRd
3l/r70Blc2MjwEdI94vIFrIGjYfsMyfKyPKx4JR7GoqwSq78IjUSYNfpwc2JpT5a
ysxsAimFsE3l+exLfnsat9fsjHH2U5st7v7XcCua8c7QtGLkEUdiuXX1ZN8aEpn4
UHtaVsEt4vms735KN3yBx86Kx1/xpn0U/Ct3a7IaKbqvm2IZGLBMlc2hbBe3V1CD
nMurle8fWtma63QWI0KciK+Evofg9IRE9vhzmyl3OBf2FdtPa5/p9H1A3mZmWEla
reGnlqitZcjZ7+K+5Z0R07NOA99eSwVR6fFhzyyOcGC/gzHacLMLPPxjxTb+Pe/V
CmsyLQmY8oWP1H3YLCgihTAHgotsP5/VyvCpgKE3+toZ8m907E0ZpLcMNPoRfykR
5XcGntDo9fMEnpa47VkUDdfrPfsbHOubN4sDHk/Oz8Seca/u7wAKiMoPLOnymUe4
PqoKlIfoSwJZ1gaXeTh8md2U1g3b3HIaYc0VcMQtxdWAaURqDqJe4M9+/xJ2EpDd
LU7r+UhAEmfYBX+bCpSPrCnYWbUi+J9T0Ohcojt7ej4uWsNc0yLyVnZIfMroBTeO
D5SjTf4Zg0cxXz81CRc9LFZY6kbrvTkv9l4PBLEKN+lanmm5FdGYFj6K8kSXEpgv
2cyLbCfA4/vpjgDBJ/TEXCloTxAgfrel7+n+UEPgAf15xabgJTRSGflo18DnqmaE
CrFE5J96PxefETzHCaYPSlWgfp/cYY9C/Uh8Dw8/ovo15vPIhstfafNnN/ai+pk0
P5rjdLL7rXd1fnSXzQcUofTO1TF8TGEQPApK2z64QKD8hY6/UV/P3ulIR36jSPAr
EZHJVGLIHmO0DWjo9yvtQhF2Il4RmRrMSqXZ8mi19P6p9dBpKIyIG90BfTG966mW
NL7lqHncKurl+bHAC4bNk/wR/OBU+LIg6hCUNukXOuTrUgrlmtcM8Zei9EvC/AoY
nvHrM9DVq7dtR96nNqnbL//DWboCi3HvI+giJkzN4qNUxVheieWJVtAaGoyzo4kS
OYkFufqptdkow7OUD7vPabGqQ6HjhTHw0v1POZhmnmO17vBOG7WvNcxOLSuhAIa5
vC3wJCkvQyV3hmYP00vb3RXxdcyjMxa+ahKzLsflsL3ybKZEDLjanYOYua3vTs8o
t+K8yxNfXnULfkA0OVVOP9Gv2lEW9kOttba1/RV2AN3vj7t5cpqR4QyRp+TCh+5K
A5HcWa4juhrzRj+93oOZKWDoc7EGTPs9YmR/TdjEb5AfmmF7I9PdE4n+RPnfJexp
kGbDoxZmJyRuIdPAndMKtbzrr7C/2FIvsclgA+fGkETF2KJhGbb3LkV9yVzNxf5Q
yYFcGBYztFx6Pmnzb0a0Ewsw1wUUqldSKMVQiMRIXvYrCIA4WmKoE2Ss02YINaH+
xrdyCiHFv75WgWz0x7pjk2waz02+4z9K/bMWSj6keUs2t7eBgiJ49tK1c3Ty4CzN
/rD9j+DcYZhnR6AktricVGMi+sYRTfGEAADb6SAFczgM8GOwYCScbzP1GexDDcn+
TczG2OpV4+xyhklzgOa32TVYx7TWVu/2YUBV6eMlNn2f1718QkYZ72o/DwnlfCH/
doMi/OfUU6O7W3fg43bIyKqkQkiosf5XDj+komNW5g2PDC9qmqAbBJ3DSfUuerri
znHkIScBrb4wE7DBUAA73IRCFq8QO1I0oYcLHmP5WpKAbZz5F3MsA1jmfJurZ+vh
8/eDZV6PLUByfu6ABZGYwCtlh31cceiQtZmCFmB8oxZYANUPVWg5nuIiyicC6cF/
9Ac9/vU9aTsZa0O6m8I51RuZfQKOXTOTvIozQVTXeUtlfGUNhLekb1qXobNQAzvt
Q5UzKghjhsEwL3iaw2O8ZA4DbvS4bSAylzZRQcds4j5QK8EFS3x6J96q+OvxDNwU
jB8QL5bquvXvxN/TT59bB36YrF1pnul1TaQISC6mUr6RznNpWmsc1dOPqBC0+O5s
33K2ynzDMZ5NQFSqtUe2O6wuv1mHz3ofmGATRSxkHfFyC58/OyaVb31w0BeOMrIZ
bSPIOj53YJmEWUVSe7N0uSeWgK/s253GqeQ6OJFNQ33IpxzKChodCnrUVLSLM47k
RdWBrHZC0Njfd64zRK1KA4xlSdJWBcp2kWnmCx2wgUYtsk+O2WZlz7phAP/3rFaZ
+ZkL8vi6+JkoSYjFloUqCscWOsI37rF6I9BrYctrS+hdciwe8jKCoa2vaxTS7KU1
vIPAAG896rZb0OpOa1tixvMfhJ8xZ2PfxHNWJyn6Xr0ktLKxiYEK0c9bJyyzM+H8
Po2Rl2FA1qn96UtPbv6TC9ZwYRm3q101ET8WYqrie6hsSn76uL4L2RUO4ofAs4h0
3eNHcuqh5ig8aeFxwKPDv/0fls/7JLXd2AYyNBcKJR7OnE7QwMhBpxBI88iCZA5V
+1DO3olDLEBGrFBmN7Hln0lLoD6VIe7vJwhf9SAgZIInClc2bYtWRPLArmJ0Thfa
kX2LFrY/kRCZcJy6bxvbYWWwfdGlpLevlfTxX4YwxAqSaM6Jz8/bxrBdkWRtctQy
ZtONK9SKXeJbqe9bNdK0RZoX+c+xTRDuinY1U7NXuc11W+vvwoqZGjbEN1OYoKUb
AECg1B6Yw0jtCW84LrZAVWhbKMvYl1+CGIlYTiQ4Dum3T7R44ln9yXxRnBbv6chO
piObDLZQQvUT+kOVOltFB5CFmU70SOJba/rDbrhv10DdP0Cu+4imwVddifzaZ/R9
Sjn+lktqsBVKC7mqyJr8JTBF32Yf6nD9sPFtqFRHGuwXPnyXldWpveX+4GL9y9UR
mExzLxLpW3aRh5iEElHaKuyllXGzanKqngznOYsIxwQq7V4sX1Cxi3aO1R5jeszS
UWxvbvDXg1JIQNa4S2/oDmMyUfX8mlEiugFRFBw93YdHKheDoRGEV0IUdQvgcP4u
GNR6rla9hzLqqBuz3kTIuDthF6ikvr9Nst6Hm44v8WpYrzljXpPtJaFOxMyIZvQf
FBClNct6vgcb2cN1vQpSjU+50lXgshBWusfeT/mqqEhrBJxW+sDXZfEcCkT8hQrw
ng0VEQA9mUATrJPZsAqn9vNvimKX5YIwPL5FRI1STJqPYqFyh73Sx1K3Oyqt9uVX
1471VhpCXEPICMZL1TatBcCLy6Cz1BwG74FuyqSFPAX2vU4uxFbYwovGk0ZjCEaN
9a2mMJqBOjT5wAEDYMzE+5O7LuL35vvndX8f2QMf8l4N+GqZWWy5pcOHbKsP42lK
j+AFRZRE9i21uhDanOMnPUA4GkJ6mDCG513oJDDhMxgjZkQrCoB9RFHwdq9NB9pa
rbZxW7U1+GjeOQtFNB+SqNLLbGPP26Db5J/7giCcCJLNz5NxBhJFqUQ7Wjd96PUf
TBxzVJRubz3Ra9i+g5bNkuVzgQqRoreD10i0CfQVmMh/lqoYO36PuSIpNBvQzKkM
tnXx3KWqU4nM38aoOP00m0UlNHgEnez29dKArKi53MnQXWAqZTd3q1+/JJyhNwO2
7hjmEx58vmzEuJaQr03FuppfsFptjOvqF4Y2bLOKV6W+ildGuakpBfyqfaYYkk84
3a79YXr69T+ZK/DKN5GjCMjVCoTPhsqP3SNIDrU+i4zPNc38RHE8vQap3PNgJhWE
eaTLqtYbLMfdTrfMAoBGflGsRWtI8Ukoei9DkLNiclKUnzRTeoceIf9yRH7G7w+W
iwTRzHZQiH11B8Idp0CSwgKrDrHwuM4Q/RySe++ETESFh5NGMjy8nptc4iMyDIrP
SCw65SIZFlVWdnMNnIcTVgty2dn2hc3MS3MQGujOwH4GpRWzd/5+pXqpJedNhUM+
speNuYh3EeL5EHFdRiDOp22+eQF3CjeGxRg8pSE9ZuV1jm6QmAtm/3gCBBISmCj0
OWQp06hK0rNfvUBCcib7q2c47Oy9LgRe2/lV8EwnS9yqrojd2VvaUWbY+WbFjoSq
kwa8J4jgyaOyVC8U3PwmMPptECMZ6pSd2MHDleDpeJOnENhOBkGFILbtIjs83siH
H02oC5heQnRaVMHHblHU1n4sW6ObUc5xVTrTZiTWFHE7+gQJeZIFidNNoBPhRnbL
6/yXQtFqy1Af+iEBbxQRD/DH3HxYqkX7Y6N1jXSbeHPFmbVxrso3tLOOlZEtKkPN
O/U4Q9RNYEdgurg85IDOBgdrPq4MqYevnpS5jMnbarTYrcN/XSTIRUNIRUmfJWNu
8+nC8eKthG1oITEPacQFKC8nspqG+D/BSpBKX5GPepbObitfxwr5x5WbwOLa7/EQ
Nma8NhFHRCrhRkOB2GgM4pFPmGhxVwJsGwkJzitd80NOHRLEHjrjZVONhESvmkRb
8fiT7vJXceilB08qIltqDayxsGKRkE7AQiU/kOL/Hf6+RnlQmw/8bDM5q2uvXK4i
XC/NT2nwU5L+V9tWaGj6k4vKFg55gKPSBFdkTjjBlytsFbGc4wOakBTV5r/2aUOl
Yg5Qd/W0ERc/N8hUt/rpzu9Dj5X1zQkGNxzxQKQ8uIWqSEkux8sKRcwBdHVaqHzH
JrkOGcME5C+MRxIE2pX/ONUgdVbf62NAFzMb7iZSqaCzoMzZeAqGD8RYbX9qyUeE
NNh84rNK0qrAgPNVSpM4rb1oR63DxTrqjO5oVrHEasifLA3YHik021Q1JIPrf8ec
63/TnM2UCtRTbZj/PfFV3EZPfGMkDhHUm76/YjL/sarUcdD69d6OMfhcWpqIwhZK
+8GTYVbgBA2f/ceQgKOE3nkT9kgAmISy8cLP4hXHBBz/PmLXYqEF3iaGFMjl9zln
dOCzQ8LNpA3aF9aLpZoeWcgC5w6gWgQHNitbrqM5qww3QpmepK4hwLcHJI7PwNUo
TU0iRNmPKGsrR4+Iy/0c0GcQyPV18iG4ko8Oiks0dzmz8uGXcOMB1/cUZI8nFpH5
MwwgjC3JRimJsVMceFr6rruPO3aUAUyBNO7OtyKz6anu3nrE0DMnByu9gYExmJ+e
aP+yxUYEa4lUHl+dpGVz5Fwz33VFCdmKONDjPSX5WB0bBwhQYpN1WVG16XriX9hJ
zbXUGkGoakq+W6TF8fxecbqc3W0y6haXkaQWNjdyDjAfCx3EyKVDK6IVP4n9XBp2
t3BUKNMWMmHgxY1oEPrRIi7BUIndIULgrmg2cAmtY02J8scV91pI9BeCWUhfCb/I
t/ykH2fd95UWEHd1TVU1u6GvCQR45SJhfGaKd3vc1FjFgGhNg3a/3I5EnLpl0+1B
HvUHUolCUA5Vao+pzbIsS8Y/UWG36SYbHzAyNiFQNC8lsXFdDnmwq6X4Lt9g5o5Q
SbGuvB5eG17ySR5/0Lz6rQWsv99tPHTYNUQJmLYiKnOS9us76646D47+qWaqkVVe
EHuPKoQidxMQZnwaPOQl9TRCAErqm6E0TZ2mkuKTHptjXzX64IrtW26cLeVvYGEd
OoZ+oyh4Yl29/iAd6IMnGvZE6NvII4hmM41mUFGMsI6KcV7HCMuXrRaVJ6sSOymE
208K7RemXlUZNXSTILYKt0VCwj9HcjGY0MG0DrREERYmwOMtId5pRQdlTMEz9Mk4
/CjJvefskKph/tuY/OjQTVl8s3qFqektTGo/1JDtLVr51YUe7R8/9HSNo37G/IeR
Eg8igYbB6gPLqxYeTYqStTd8krOjECKtJWQBmT7a6b7QowoSfiujMAEosVXWtsPn
ZDbJvZaadH2m4WxhLIXSLlSpPsSnqPRktnEhW30CxewU+xch58fcBXt4TqepbyOc
q+H5HSOExmTDiiVIrojpHzbh2wlyrWTYMu5c0Xjs7/ggk7MzNAAvncZ4qDhhUlv6
gfKrtYHApZ7IRhHs4rvaGhS3jvPEwDM8Ad6kE9JDh9ka/DJHniptDSCKlZM5C46H
qm4yH+VJc3E1ulfCuNqTSrVCG5u047eLIRjml6+IxNBlB+b07OIa0oiOWOeaeBqh
/sgd8mCrz8BEGWyQGwj7nG0JcNtTDiyR048wzVAx/FWdrX95VizT4SVRhANQzk2U
JFjjKygr6m3+ITpNzGgKaCDEoYhkt224hfBR/Fk72D0aLdibSLsobU/8/qZ7bXEi
3q3cJZWOvBb0qwfais9qF/2uprot+yDpb9R7brGRz2C156lTczGbLF73MaDaBJgT
MPq2M0/LkekYZ0T7tdye+ma7YpGrpMMm90avjq0SPM4Ktnov4J6D/rVFy4TuV3aI
nHlaVI1vIK05fKL9kD7JQNRSuVTmBV6wcltpWUssxSw6PNMWZrgywnV/GaSnHJPP
gu/QCdKKy34TEk+susFeOq99Pdv4WLUmpNegH3kfWIRJQxuTleOx9YLSZ2v5MD+R
HkfWIEFxY5wvck/zN6aG80/G00b8PgEueFjPquaSokMZ3wgRT4An/H650kjPQjzC
mRZoskhOArBUXtbXiQDLF7ZQP0RuTmzoLDFgQwB8slDM32esVEgQ1OBuJeNJvYzo
Z9RoTIzC+7UEF/zjkHQhP7tENHWaGLXoMcwLJ/Pwox/OVp53UjR61iIgKkO4tZfC
8hfiCLOuqEtsmE/axFDWOwLaIdvcgyT2astbjeBko85GBMGmFg5I/QOQeUJ0OmVB
rOnmy5LiCGSO3uyjxXTAhS8oCdLGodoL+R7VEY0ahykmk7vSiRj7mmS636vpsYxX
fzLq3M0IcWgyLmzpZ/TpxQ0tTqIZ3rf/8Id+WqVCUJu1Wr+QYr5stLWhGTJvsTBe
79qBJebo1Yx33QChfrRpEoenNjK7kYL2hm2uCIbbI8zorBbhT80k4lVLp8Id8FnH
R7omgBnUqOdGyzkzE0a26+qxdIYcTP7faYS8C5OHKvN7USB8/MCtOl79VCiGJkUB
YreEeJFGdH87AblqjP8J0/Ej1EyI5NMj6ZclqTPlCe207tMB44sqlRXkXiR8oWQi
xTK909RIS+GrELpg1X6qWZ1euXgqRYOdOd302+bbuLsK04Ewk0AoqxsAE1g9b9CB
Hf1nQYDG/qFu4QUClZ4gvl5hcwdBm3IqbTk1mc7v8xfN/F3U+0x2wR3ew13mJrTg
rryUaPMC4PoxfHtdAxdM9Bon69pJpNYmbfviFn2tvQ56VdXPRPWUpedBnmEdVnxV
iS8CEKx96jCTZkrTDz/ZJp+D5G5JPAuRChSB4xia5kgEX2P++LVmkImMwwT1Kfct
HEuI1MxraUATNppXsnNsq2+pPFpAFZTiexGwx61OHjOTEklXwYQdPAVo+9C7prsG
hrtDITf2UiAU8QcoXCa4Z7PB2hoj3SBZpVsnIHaeEdLwq3axP0Fxbp1n2BwczD18
UcgzZ97sQpfNn+f7aC4MGQrO1PG6he0Vdmv0j7T7WQe6gzMe2nZJt18Y8VH0t4td
oqt0rhjr6KFlRnXX8Rn6YOVwiLCVX6gj0oUcAlDMw2g/NwJinUwQarAKqZ7YbgS7
gUejsln4y+E9i7LMFJ95z3HWMRaK84MgCK1iIR5rirdEqBNVvOLhtsp1XvbnD/Mq
FxRjS+E2C271c+azc6Gsn99RHFJn2fGmSpY6AkZ0RtONKMH4GrmcgThNxev5frEW
2W0awhMxe+JuBNXdocCClQkZ9/iQq6Byt31ZKlWaTgNE2yTqSU9ATDj1i7ncDFS+
sW2NHPconz806/a5OwyP7450V0I2azTCm1TX/oOaVlZxsK0/moMMt37Z6RN05uWD
B1UK2Ic1wjMyaHCB3HCA6u25djXyocs/cDM0UvxRFwRMWw8AcL9qqhonjRqwADv9
y+GH/eDFR+06OPy0TZMQ1an4ZLHZ4Ntp6yUgdy5P+bQhufdEFsXa4v1IfnTdhgUx
1fgnIXrfozaBkBkJxAxgdpEmKqxQyuiw7aruPTRVXOlLfRM5x5sbNLSm76MjmyrO
+M1+90WiAcwzvmQJI1GVlgpXGdfQxL86c1pElW9wpJKu12MzDV7gj9dLJc4DP4FV
tc6Jin+5imhhzKbIxlcO2hgGGqjo9N5QtOQZJXXsUyRa/xCbdyqnkeNNLLbw0uyj
DVb+32CXLdObCVe7cjGUw+pUbzUQUckkKiqDULTFzeYFIBMBuFvSAflXnD7Mv+F9
pMXNCu5CVeSBF5xCXX/YlSxek6GWXPO9LyqBwNc/GHubW2N4ote5PGp7ZaV1yfas
5qbj3tUHQ2sY28WlgCgeBNl0iknpzAw0mKzhoIQ2PslQfVvCzIiNMlEzDHDwZBSW
HGfu0a1cb5jwJCUJo5ntJKoOwjOyZWfgEn8EjnheL2V2xBL7Gl3N7t/ayLaEF1YQ
mcTR28gtLMWty0gW5AAz6txnEFop/TpGwjxqStXVC91W6VevUm+b5GjYa58kRm9s
mW26zHPu97/0ojYTgqPzL8lifyr5ygw7EfopT1zUham6y3VVqxGqhmuGjrGngY7L
BDIctw2TU3p0Hhh04tPsHhIo9ZIk8bPg8d2Lkhj2mj+sCL3CeGZ2WoCpMdnnJvPc
CPpDAPTid74x/EXC1NUNFCt83D92BOpbF6Hck3mozMHlVkXE5MWeOV9n3bYcdktx
NMy1DJu+ngc7CEddJFIDxuPJVq3VuEy+C9fvYSh79anOll+T1GqAdlk1SPczWMUz
ZilDyYK6oSdy5+68RZue5rE633UZPcjGjKVLJAwHI19x4pGqKHSGzcXZS2gD6qup
dZzRzvTz5Rr2Q9YTG131lhIAVVVKSxYCMp+c6bld27rFKMYdbeK+IGkkVXdthCGW
34rbk3Xb0PvxbBkzcpuHn0bTJ83fcBeyuCpZopPwUHyQ3sBXcbtMXQ1hyPGWTVXc
18VSqUsRy59K6PVNp0az6EHoFJrixPYH5b4VTdHaAjSlZ2noQkL36AH01nIJ/3yt
OUi4rcw5R/7BCxb5VdaLNFss+tDD4JA4hb19WIw96PHAfocJVd5t0/OMY3tXz8v1
hCSx3NM4vheurUkd1NF/MoDmzC1i0v9P+rB+V9Ueo4XiJq1X3oY6FhHPLPWtTDJC
JPHPOYi5OxtHrdZFB1OuFyOyri3Rmv/gyCHGPaC/hP2PJ7tB9S+sXLYu7q+kWcTw
jbyeuC2lf6eP/S0JlgMI9sMuhALQQlnI1CNC80f7yv8NBAvybWtrc4cPFGpLIAEM
6SCpMCdd8ePsb79ZTz5Km5KUDj/NbCoKWfrCEwKn1Ixr44BU+q5i7P4faUSFDA53
zuoJXJ2JcHAzQMqsoY65Rx9pi4uHtUmAQDIiwvg3KbDUD+r6/k1SW7bar/aMzbHm
1Dtto4aqJJLIU7b+NzSmCmHRaROpOCaw+3x2yt3x+ETvjd+ErBSulspLasmA5w2/
F60bmFzlQosXMBvUVMvH9i/oxX8/ALLAUXmk3MLNiwbwB3UVGY1ZoUaVjuObZgUL
q65XFiChafNT8HuQC0q8FM4HEnS1GWBfzHF6DtMSorpl2dNvhc4/6bX3c7RN9pSS
Z/wTt9yS2jXQEDZmkrn9771YKppWkUYedkKLEnwJ30uz4fH58KQL0e9fZ7l9RifK
N/6plE+wduSZ/QfH7S1nIAH5RFg2GFV1tKQUteHHQmdS7znRWMMoO+BU6t7BSnGR
2tNIu6QGYSgFxjwMwwi2dYZ3xA8hEIfSwWxajsD0XNQmAJSL9/ZEYmQW8U+oWYTI
aVXAd4A/c3kOY3KCBipDbyHt5NOGkNCSxwMOFSv1JZYqjJ8wwNfpYszForTuCnmI
iBmhH+U8qKpNewt2JmiCvuCbtJsoQexxoU4SmNb2zMx2qRszNyDh9yG6EjvRmhG2
3lNpvDz0OMOZcXVisnf3/cGu2r7VL+L9wyv01ltbwkl7xv+9ptJmao6M4j3jUqV9
PXRqDJ8MbcxanQUj+nFpL90bu5JaYLvs8VkecjAvZv4rcwamgT424JqV2N8VfagN
+hbfbCjmGRtG68u0J/gAa5eTXt0H7B/hgOBbzm9l2YgSFC9l9XCUs091wPrJyIAd
Jkm91yd0YnbyXEq4XrZLdQd43HkiE3ogDUZRDO0EzM8Gzgepf51mfNuOVMRzDafe
kqTYk9ox8ke0CFEzuVG8A/51JupmVd1gyuzyZi3kV0rjicwVZtP46HC3kxTP0EZj
wt9Hs/ijp1Cx4pbCpayX0YnvoQopJuxLF0p9bYFUfTvjKmEH4YGi146/SUbb2rSW
Cdj+kSJgyVMxEC1l9uGg9QR0e7upH0K7kUFx9WBFg9QbdhhXKkw2XbYcar28LJm3
1vZHA8Njh9TjZH8f1J7UvkAmCDTXjDyX+PZ9bm6lBFCgCjfjGW6GwsyDqPt//ZrI
IXP9hThT3Hpr+uyzck6I7v3GZYDgV0jYrMLcgW72ZXfHrAS39QMDUW43R/AeqZ2q
6gMO+RF1/CgT4xVNJisYFBsDREKDiuonFCSOz4ItGMh8GCXc4bB1/AnmFneahuo1
3FoRDbwsthRm+Mw5QMsP2Y6SpGiq22h+o5/YLAVoO+zMrrgz4rv/eeOpf0OmgfIY
+1MVNO4iLw0IjfA3dPTi1U1Bl+ck7RPfFpp9qxnulEX0zObNH63+S9hYCZqKQyj9
rssQYLkRwMDQzoLJZoDFF+TW2c3/ndC1SDzyXr+5kPtUE8JNViBIVW6utADiRPD7
hMT6XgL1HF1/EJJ+4UHUcrpNjU4affLQHGD63J6coPKMzV81mW7BwrhUN1mnD3Hw
I6Os2abM9XtrF3MJYp5cu1i+DLQrm79zYQl3KHV7IUQ5kK+9hTBcyhxpywnWyTCv
6Pc8MnYU4rEWRX0mX8/q4Kowwan6aGHYsIz5c3g4QG9NJbcR8vbYbfi4MSDUPqay
uvmE7G4ZySGAoXN3XccdolfUooIcZ4oNL/SURiGa9d3DQvQF7egYV/2fro25/PPh
DwCDmdpPy1uJF3WPHHoD/C3JnTY30xW+LUcIZZQ2NQE9+LbbtdXT0F1xwB+FJbQ0
p9f7W7rwuRoD2r4OSX1EC4GDJ7O3rMDod9LnpH3ik7P2KtQbMof15H+NmAk1EhxH
0C7EULshjNGf6budNk/gbs/3c9Ul6x1U+y9kJ1/+oR/XdYiiuwBDYBRdlrTqZByJ
DnRdW93RLMnCCtJP4KuCtcysuY9tG8+SB0NGYOBqk/ehnZIxWG2vD10ShO47o1OG
6Vv/agP8BrToj4fNXNTySrHNgkI9FaFJ9wcqqWB7/2fXdSknSp60E3x2stSzvSEb
euQU9CLEMGie7sKMyIu5mWoVAnXi4vQ1mWLBXkyiVRcRMRa6e5Ss3uDqbFh2pOKh
ykSuu4ryAKf/NvTlZwZ4zH2O/8wEMHbE6hK8ri/31D54gqTi5ZBscHwak5aQ5ZRA
Pee2/02K1mwqX90FS9ZEv+qraecETfJPXXi8YzD3wJYM5nzMyjXNsFlug3q81+/0
61m6bu5sD1mTv13WddAfmdod7C53hfqydm5pKiH/tXW2puv5ZNZz6z2p+apzwaEH
Od41lYBEK2FzkC8Qi1hLfUNZSyl0eyvKRaMtCesz2E7GTQf4LJE6Ezmul8c0xDLt
06woz+Cu9pKQJE8k3Mds+cWnOV5MbDcXHeVe3vGpepnoMye8r3m5TsoByTf5E9nG
ic3BBia68M6JSOE2xz46o55RMHw4/g32jhM2LVMYX4Rv45zQ393kamFPrgKkAhUo
RimALVGmqjlAJb5dRsYwQnINAgDZtyME3vzb3su9lhjXsIjdAD/7elRL2KA/t1Bz
38cx5h6x2cFuH1QfRh7FaWD5PQAPBWiZ7dy728pjc1rzUGQGL7RJVx8EaA7+6zfq
HzgWazMHxyTGGQjAk+LxBGChWLOnzcKtiSrMHbZJACldYzF30CPoZZveK8H7u2fi
K5B+G65u5BNkze8VNlBQoVJJaKxpK01ewz8fHExP+ynJX+SpsGQxHgWD3iRv+85Q
XmiBlVzkEEj7D+7OGdLQ4VV5AkKLGDaFz9JWqpNKhU8UjsvGxe8rsX7503dMnJ/Y
h8zoEUrzV1XmhT+Mz+mV2n7rjZYBj23AoL2dblINk8Oig0JApkpoLgCL7qYbj6pR
GqwaFfVnNQnNd1qxJR/tY/YZYz67TL49vJgaMegVGHhZxgeqVuIVEW7zadoo1bC/
JDzcxE3abgcnf7Oju2L5LbrmHjnlrXf3piAdfa4hDBgjoC7zaWkTVA6vaZe50aII
HqlaUL8v6YXUt2SHRCq2tny/6xI+T9+er094uMaurhLnaenwErQh8brFhbkYFfHJ
SDHLZsKltVoymYaSZk8o9wbOscm0yHpaI/I3maneFRGrIvOCs5TOVhxVW8FxPnni
dSRDspcx/EXv+0K2Ql56spOaHrpUDKwUuvDK5GKwLIHKFP0TirVz2Hyd1CxLMp6X
yL9V0No1/5L8tK6IN2ERK56xUPOXhehVjuziCc/kKAgEtTD38cgbgCosyBxkmOLm
3qzReuHrE8rmyycSki7WaO6Mq13cskd5YiQI3XP4i78j8kys+Zhcd+Qru+t/KBIt
mhJZVXo7vSvpXs7TvtqL7Gj9tUnRf6URMLAklQZ+u8QP8eoMp6Ql1oC8MoyizZKZ
MXbIb719omZ5DPlehoefiJ3JX+nkm8k5NlU+rSB+krbkIZR69vN0z/kIiZEImwQR
ibInQfpiGxEdc1LbIc63p5+BqcbK+dJ8B79U5HwgIQOliwAJBEUi94Gzp+qY+Ee8
ASLOvQZpeceqR+pwf6kGlDNRIGWTSDfykJkZFWUcCQnmBdrdhCztLIYSzCCIeYhg
C9mYH9khjqRm0FdquRjDpJRm63clpE793VlusLOyaH1gnE0j4BEm4hzX1L4Vfghh
28oAOgv0o+6h3L20W5NltF3nmjwkfJ6uBze1IItt3OTzyM4LioYK9XZjTIR5OVV1
YYkRWrex5h8knDWejCakX+IzpcqDLIHTsoMYplyF2RcR8Rm2Z5WaALeIVifyvcnl
mADEWwbL31Upp8rVC+chZqwOqeKfo62ddZ/CIHTPuHdM8ougr16jFUCTxSkAr17R
DcEmzcAGZ/acg561jRGOBuw2FW600YX9Ar3bhx1spf0p5zbOWL3fxiJbyimvj3V7
GScR0L3L7hzmPdUKYzLA3a3lkdT3rSbuFkLZungCLjCdR2zXZkq7jEBJsGcOnvU0
zQiZ/nsAm9/yfWAwMaU7OXQFJKZbwApW5DD9jyDmf6KJvk1HCdqkxn2FpomOmZrU
E4LjoSXHskN778mreW5aprV4Tg1zzZAJE4CkLl+2Judx1r4a6YD+vIxZX9ayn8B9
cGKP7ygNgRga4vfW/RCwa0pd5UMTuPSIoOjZJq2ivUvmobym5M4akQXiV++OZZyA
20WwT3GIsJrOGMZIThIlOY/KFQrSVV/2wsuELsK7lvmLe6EW+VkjB32TXilgC0sS
bWaOddBozZ4B9rgYmsHRjAIckkiUY23EY6+q7FtCflOSKVn91DjULbhsEAWwZkH0
h+6YXp/5556nTMhwowt4PqzP93nKSwxzlbe4PEZ0vFhdz7XbzQUGMBSKdEuA14Dk
vbGqplSI7jBjpeoKq2UczksygBXTMUAfWjiKLv7PqLQHlYvbxPArRIoWjJ16YCFc
eN6ekfm7B7V9At9cBmVBbgYkghzG4aWX0YxgxK9gdQT/ozn7MAJrEmCwd2nImum8
lSMuGKZMo79k2svNjAto1MP4Dq36mH4oVOwpkAmS2n+mJlGvWxdGVp7t4VURqOUu
f6j5vf/sY6y6HxI8CRTe2fqwN0ynoxtRPDdTsVEyNwv9WavuvHS+YhIoJFz6u7Z/
WEpwQXhrAAAsB4uRRCvk85q9w2idKxXGXOOpVqFoBymoFUPLt7feJ3zzk9td51Ei
ZDEPm1ozkDUOTznTyy5PMTB4ngTHgYzCm5SDPwIu3o8FVtPme9Zb6PAZ7OIYJnHd
X9dLQ02m/Q+I/OAR28jcP6oIXqG5O8kD9w+H6WRgUWPd/fSw3hYiundejAn0UFpn
yYMbUfhGJPUAHv+A7k6vcfa1+T60TKKLH8uQmGGUOPQZChOKdAZ2RMCu0bXKd0B/
96Zeq01TLlQu2JyrbOmK0FdPnjo4fUsf8k0G/1h3Mvu8gr8M8QAQlYTnRY93yNIB
MI71iLcrD6/W9PnlZPUmbxayKwiD69eG+8pUCfwJr1SXEsaCZQ1yLnVRbTa0wOaJ
wv7v0WVoP/Nzna6VeBpC8JWrH8SzGQDUB9O5TAgsadwtEW4nkC6/rRyCtlV6EjBb
h204x4g2TbTZtMO3PjRLi0rvQCn+4uqurbR3TGHLA69zyZbRDn/ijXf2ckrctGwI
s8nmz8k8qnb129mBJjKZmOj1fnfIt/ZJeAOqN1+aywF3ucxrtc68wrADkFd5u4cc
uRfgs5HxDao3HidXA7jHUj25PwE2XSihThjRzAm8ZT/yHLx2RMsuh2Nl619CGSJ/
TGnUz84WBkB8Mw5nnRa0U7mCq+O/ZvE5vGFYjWnpF1uFTpz6BvoZOModldGWb5/1
gnIjtTJBBXWCw8oXM/X7cV7tXuI0xqXT/cUdwR2kId4Z519SekYOxywSd8gL441y
sLBb5nJbwvS5mOF52dTN1IRIivPfJi0qchM8+dJ41+edT5Ne/pdEQPcchOEWel2o
tdZc1Zm/PwnBmpRiZSlxAE4RcOJKkjt3tzZbYzb0EJF6mJcMaiw3wW3nz9GfeMs7
BeMlL2APwHWtyxG8azXisaxWVo9QsWdLLSV4sMpRXzD5mnWCT4seeyje/QI0G41n
mO2lju+nibvLs1oZbRedX4r8f9tSYvEVq2orXQJm6hI1ynKKt8ASiAukxYLt4XzO
Al5X8btzZDhmfMWsQM7UxFMyD93RyAf/pQOz5RhsoXRKH4PPwAtvBc0nNcqtmMIF
3xuLfFQiTJK0kEdhDVKjIX76E6RKBiVPAqCg1ju4TgnqPKHfOFSDzKjz/Ulactjz
GK2i7k8Ei3XR/wfq/QUVx/ej4qKLDVN3pBAPKwuGphhkzJUHfpieSAgrJzBCc83x
hCvJLSLu4/WKWIjFDj3BSlow0PR4Upu1CFtiYOv3uaZijZokBpNPLYNLDK/77JTe
74E3UXjN+2B1sNNAuvK2tJMaCyTxLie0eEeZ12aI9pgnoZhwSSYmRHzaNgsXnnxi
IK0z8yWlzFesDdeHXdMS9KYGvMrV2dzc+PYgHLSK35E+tEswnLDLI2ue5SlBeLAQ
bNBSVNZEwi80KM6h15eCuINKCcDVvKU8LE3/4EOdKMT0MIxfJrmhhmprO+sqI7g1
kuzQ85kFK8M8h6ApmkKWvVHnHc1uIGxj2B+zPzWe5SZh+synDqm/Aakrc7f3AquX
jMpZ54rHZPngSAop9Twxb+K22hLZXLHxLLIy8o6bPBiaRohrcFvX/iEQtb+Fu/MN
vxC3bJH/45Uw1kuW7+lJbIYKPl670KJgqHlbrZNN3rM56HYgXFappjrHpjheKBJQ
dJhBznx1MsLM4FSOPwqHBIDFauPlH28/x9P5kCizWjKVQkKIQNd9e2RRnPz++5BB
o40ZXIzy18ZeuI2t+ull06zEc/u/LC/7sVZgZpMJ1Ft0EkfRhug3HVj3ki7BX94k
0QXpiJ6rgeAsOv51Qdcf8T//CMt5UrzNVmNBHhVWYTUT4zVNDSrNWw5wrNmK1NCI
GzeNPBPypFPha9a225sabElgH5zKr/hBjExAB2XH+AJkF72k5H1ZH7/GgEWa+oHi
+TKZvsFbAy11FzFk8GuDbTkhB0fcm+D4DE2BDMBbeRwY5J2IIU0neDAQBDOnmJ4q
trHSjB0mBzpYtTJUVhNF2iFQPJZJXSkBHP6KHOaXw/W8PKlRMjCl9VPKBPuoFcFr
51U+6qtcUlEGPaFdbm70bes5b6Wg2pxDBBT85hdTGPDmYGFoGPhcwougqul31EU3
+N7vWdD4/3FYLtrdozUlZQwUzVUqWlVDsViUrxlA/s+qqei9iJqlTOZPFkA/TQ7t
KvwSsGIfkAKyBzog2juSDR1S1JRARxuuagjn881c90X0GhxHNJWZphUCXZ3vFIRn
diTVe3PkzIPplBQcplkJLAF/GPOtbM3ko7WnBIw3nzDOZCpgNFB+8jWoJAUmra1c
NsGBIQ0N4WLfMHo2mqWb8MIJCZinoJ/izP5iOCp9LH1JaLaG8bKF3EaifQDpaZNQ
Cu5obZajFDXQ+MnxeLKuj657Hn3vfWMilkcCYz1wdZhVxICrymDd8nHuFqkJdoKx
e30DsDAZQzxHrr8RymWz9qaYMy8EWCDVxpHjKQnSgRvI6v2KzRJNlxOpS2YIocjl
8PP2xjeotLtzHMOQSgOOmS0qmGMuzzotsE4AuG7ViW82UxncE3HLdHFaOx/mLZ4f
ERKmThimYxyIMRP4cbqEhLF0QhWSX0Ib/xxfEuXgPeEawwaVY1SXSGN6Kl9yNo4D
BnEILvnUMn8I1ZEwvmAbwyxBizDzzewr1sp7u1yUtBx0Q1DTcOBuMaqygYueCYLn
QKzTWrahFg7MUhN7lgr4lV4zKWFuGVuL5bjShzpU1fL0dnAVhb9vgxRYS02NmYVx
6+Yjro7B+cWK5pf3khyROQiXaw0zWY/iwIn9z5JSqo4lYmWJKZFiMhBlUfHUpdM7
6dejX+IklGE41T9MoDhpktbGREtolMURBdgMiA+l15pxgidyAxgKwAXPzcU9TLkG
urhHPB36DH+5Be/Qrh03s9BbnlOUXx9dXmD9PGg9QMQdPiUk+A+Mh4X/A9ZMQgIs
shXSgdWEvC8XGeCRsBch9mRQoxs1Ph4KZahu94HG6Qm8h9ahKzgbUCKhHMYXQVwY
838T1tNANa+UCjxPyvgVPmTplUfqVToh3AqRwgHIYt4GaClWGAL/nDqDC7bZJdWy
9umB4n/L/QeEWDHK7fOMIjVKTtCHbXV03mNOmAuGVPQLP/UAx56erkf24qEPLqDR
z82TXDufjsj5X1lATUVVs8tk5uIGKiiPdK6vgujcG4rTnHn1+iEQGTjzXM50JJQx
mOMO9z1fLggv+iS4iCgKbSDLcujcM+zZhPS2isIESNps4fE0qVoRddD/urWxp33k
Df7YpG+kWJs2vSZ0pmHvrfx4lqSRPIPuybq8Xdv0a76qzBQc18QJ62mscGVl3rla
SvBjcAGNdfR+0Ux6hE7gS8eHd16icZwNvdJhCcZqqq0F7CrOf2kGT2qh+IOFNZg7
BQcvu8WY/GQSeBXNqC9XLg7CoeAWf1dXrsDeEk8w7gOfSK8oiUkz1/pSo6G3DM28
J83fXOyh6rWAPVguIH7ynJftZ/bne9uvy9EOVMHWCfBQzlXDRBHCIuLWyMqjv/uW
ki1TaREdfMbbbwFyitPLaU7M+qNE7/GiUgFAtUobJfvP1lgcmu77mGdaM21R0zoD
mVYS+3HQfNolmtBN81OaKFlmyZ4n9uwXvk4a/mh0wuMwd1f/jWQxloQX0ht68cAl
QvnZUmwnlTgA24tMk7LxfygOftoncokPGuqMNdCZhw2qjV2r5cHwc8FJX6AFmNbg
OiFYlzr4lPJtudbSn0NwfsHmWSwOSoWkAviwjMDwRrPCUppT/01f/32haK+JZhth
Endq0Ps5xPX3gnfq1NkkwxSfD7yIk5ZUnT0jQ15bF1n6fih3/0fVtS9FxZkNEm6x
9Y9tFXHwy8grxfQzD7x9BzpS16vmIF0z7IWBMC1mriEO6YB6ZgHeu+N+6xPd7Kuw
7IMQ6ztE3OcDhzlDZnchFOLTJFKKtp1+3N5GKPBqi+/B9/WmgLW9O498EwiYl55g
FC4dlDmazbfIsvBgCsPftZapybuVQ5IGYuIRGKfcC29/jjJbrafarCAJkPnoEz4d
Yd36PgHIqCU82i4DEpaZ9ZjFZdB8hjYR9cllefa0Y7UT27HOOEVsbtTwm8w+pEIi
OZzzGtDr1RDep2T4iRlTaGLrWzP9O0z2hE41izdLyzDoIh83GBQpia92R0El5XJf
JdNw71jj/xD4AeUAHOF+51gZ7t9IKFYmcESDdEPfs4e7fjvXasPsEza9KVj3NX1e
Vw7039iCPaAnFXsFjuCLqZj7SZ+ViE2ZWzGsphFaYjSaKX9Y2pvHb54gvd5gShuu
UhizUBuClDQXO74qC3iolf6IswzHSACRIBEgm1AUzGzZY+OLfkBmJw8v6tFMFsuf
nzz3gAispXYsDPqweAM2HoCVB0IgWyvUNfaIKtzR9W9DIG1NVmuZvW2fOMhNLtuR
akOpXCovAEj+3iZAlS0ROtmUrBpO+cmt3J5zEYy2UWqeiH+a1VMeG+OWZ+9gM7+G
51Y9Of6BnK7Ipxgt/5T4uC8xQd1IU3NWhDcy6JBp0VayorSGMuOy/zukIpg2AqGn
sjjNR4qkfkYcI/qqso+oGH82j+u786Uf1lKzN6GrctWh2mDpg3nzPdQ0YGS5n1EF
8aZTQm9TFXqvzuwldX/vad08SzbHL2uekMqYGHdssZhwO0qa1/G91segAxi07g2Y
BgLlF70TEbYI98jOliszci350A7arcPoVs6bx8otzlthgdnfbkyPwibUZLEekaPn
DVS5HF1pxFXQRrSkI2hoxUB6su72/spJZ8a3BVq/TB1SSR/VSfNAQy//f1cMv2kH
2uVnc5fvIbXRwfW++pbJb9WrZ4XOStx5JzyHtnWaeEDADx/vFZPMqfhIevhCCFy6
x7BW02z2tkerf31z5QA12QtfP1c5YKvkXQENV11gPU554ZyvaZ7Kthp9PQG07z0e
aQ/Vmb7Yrge9j7ajPBXYMAGdmFmpE0kBd/AeJqOtGUaabwWC2cCnQS25KNRFKE1Y
D7tcVFF9FDspH0oKRsSbFeOEbWC2S/olbfi1+alUT76zfU7+sHi4dC5VD/Dqp59y
3yrsLKRrnv4EUHeHDe1j2nH1pSpSK04rr9JdWkJjQNMhaqELTZ1yAK3tDHBWdWDO
6YslT+KBPLMGxVP68J8G5tjOzO7dLwnEjjaTMqMOK0mx30tJO/buWfUMzY7evzHN
erYZGLitjlKd2qCHywIV16L6ZtStdFPlcf6lRfwl/1IKdyj4ZnnW7jU4WQ1vTnU5
KHyEqYOCpkaSTuXyp6N0tYhmKoOnBbGcs02niH2+MpYu8V4Qakc2wKr4sGlSMnSe
vHZxxisNEocDZixVodOpNKOrJf1DtodVgikR1cPvVwOLbytjN9I/U3WnRX4KQJKD
9nXpbQJPVupRLP8pGxl/sKXKfcBsIMVSjWYnGRf8XYih/GewlUiIeNRuQD9NHjIZ
7pzsX3sJk1VjMh7/LkPoB+wWPEppTHrEoDT6mnKB0rajgq7hFUL44XnaS7/K2XCY
15n/2jqvO+rJbhUMS9UgLNqy4GKCUGYyFz/kMWwqNseWR1MC1v/c9z/BnNIZ6SjL
w28SYQfXvYioXCxJBAdaEhx8IgaGbPBxsJ7pA0KIhaQz153/k/Et1Xj9owY8m2uh
neRlNCTlbqngeOUgNz5XP+2XGRl9/58qdQ+6T7e5RSkFaXMDeE2T9kWATvu8jZGV
6d1Wbh6TcURIRqy+5o/0or0z59IGvSidKA6Mlo77+kfz/aSR4lWyH7k/1/pMmWGT
kysUwUPL/JuyV27iRIzCgc7V2K4hcv87jBEHBTHuTU9/7tSnPCGNELy3an+rhlsz
1rDknvJfBtiYNKnrEin1XHU+A265R1rg6qr9cgmqlBpZ6NqdyPO2gQTRDRX7yRXm
q8fDaPSEZawLhao99vAUWRTeWndaxdBL4Wg3YBASaI5gRwmoFB/WsPtxk4IW+8Vp
pPCww2DIoRcegqp2h1AOHhqbOi1Zm9D7Z4v+aNje4qXpLfPhN6BWTnFNtb6zEq89
dajVMGHKkGMHz+R14nw/Jm+kHMEiPxzWMDFf8/CVPoC9INgBIWzMzDRo8fGTCNhk
txqKva1Y7A6HrGm5Zg8wdgUfvg7onog+e95un9vcnyUJ7N3I9yrHsr9hl+vik0B4
pz3tM4N3qER7Rgq8V1ZytESnUjLF9sNAYq4w4D9OYHQzfzTu67oRjbqijLyXAYCS
0AFruVRzBFEmdcCmlWExwFXtCidEUE4FBIyyCh0eVkSJ+2ouSOjeAaJ+o/iWj+sj
eo4V6OtWS+Qp/3EgDimN7dTxlYtmT1NgoKop78ElT54ifxW/3+z3pUnRN1W8C67B
P2B4+QbPsLB0aCWMQs2+HLEqYB7/yMwW43OIZtOxtY883twtJXyu682d3JnpxoXJ
6kLN2wK9X6F5B1g69JQSjRWpCpR0/KvSTA+zYbQHPhPJtK4IAxVw7O3mPUY2vAqj
qNkEkpVKy+qCICoZzxC6XWHyAXVDpDgELdbU8axIMGg9A2XhLcljaSHkmYlXYd80
JxODDo9GNE8gAv3aXfVJZGQf+iufbkSihGDUT3f5wqU0o2TAen+eXONafuBMuDP2
9AuBB4r28lF73PKgvImlD62DZcyvWe4c3xTyyUWKFd2IwI3trw9cDCzbuRxGgsaZ
GigJcR5be3hGXJoBvs9yJrbZxztkmzFvsYS7Qanp8fxPYkXYoJnLVW/R1kjSUqas
ur1oxSunG8USZdKcAezE8WGhrzQwGIBL9OsHV7V62v/k+Qwf9VJicCMigIqZ3ZQJ
JWsDEcj3TfV5fLUK0E/rubztBATE8DmSXeDgFJMu7E15ovog2pSlebQecNPctkHN
z3h3pRzbkZ1KTdj87WCzJCfaE5ttfJCSwsiQdRPtnAMccSGW6/h4u0cQAVjkSrhE
OxIwvAAdkCTtpDsIAk6fmT8BRmuHUL1fuxtNeB+dD2bdyJ1IoU1bMI2X0V1U2nKz
2He+qHZgKXOjRFmWEZWKIpK73KJDqMTu/XsPsLnGkpJ48EzQFkiPi8LYbvwEWj1G
Ps3ZR6+ZEXfQ1zdtjBAdFZDSy1qF5oWUJdMoFmKsimRXKkTLpVrpRCedECbTQfCi
Cei5whO590JyjXVHrzZjhynEPiqx/o7/7lvU7HoUH1bSBrB2Xci3U1/EzFx48y6W
T+o+Wxi17WNF6Ri+49csRBz0OStmxTc29l/XsgY2kGK2NBArlWJrhDdGMq6dOusD
vSbj2wR96QFKMlGgX2g7gKAO7uLdpe9Lj3dFPPDr0ufzsoQfCBUEdM5B9Oa8Q6BV
wya93oN9jIuMfAyLM1kGTZpuz9Eptz7sPJwFKGvDDBr3SF7sRWi7O8ex25dQ7hpK
x5IRgeZoMBXRO0ODGBcyXcVuZPIF4DZTxWtw2sMCRp+qM5vn1qIStvZZ7IwAZTuQ
Rhdkavfq8VTdzD5LkL7DkNcoLD34yq9N0ghblg8zE8kKQPfR4SB4MxKQw3FNxGoz
Y6dJUlnn2mELE2q2F7QtDQjl1VFTJBgP5YOx/6p/uC4U2FWzt3SjG2Xu6E+zo8lC
xyfjd4iYV7GIPbFd1AOmD6hy7LiqEn4HuCVVKnZDiTL/yF4K1aIp3PK3FWMX4Qtz
a/bBJK3vrRRTuiiAH8KRVPTMAaNRNwTuKlWqzkMgxUCZgXeGuSLGDW+iLO9W13YC
SHM8zfbPstPcweDZb2gZH77lyTHvbJn466ANbKN6cKB5GzUQpeuLIZCpDp8OMZ1R
MbqL/o0evvPskkw4bZHffNgyX5foAJNsChXPRVPRNcMPHJo2bvbnm0GICvFYcdJz
zjesxDEgk59wrzDDrFeXnhL8fh9PKM0iE8Q6cAsMnrf90T3r8nQGqRjut7iPNT0T
yxGKOis+/mzEjE/O0Ms/TCGXz1euHhGBuoxxme6FoDhCcWuZIs9XXXJnA2RL54CQ
Ktm0jjKKY9Qv26OuJjxjc6ZTvax/uohXbH5Mpf5sG2BTjxP37J0DzGH37ODtzVoC
FgNxKxk9Nnd9Q6FyxYeybTrz4tABb1O86wAtqwe2Su82kHfymeeXYJgngdGDq0UV
6+QT9htQ6+CSE4OGCzwaOvSk72CtFDt3qI2bA5h/2CHLkYhMrSv0HoXOTG+9/4Vz
NLE09dbZfXxfx2ZpxhB0EqImSuGMH+0cWB9FHrNjyCsp1lndWFayoEuqo0Rg7HLh
4gBZakoHQBZYMYpw1IA6BJqT9dOQTwQS3iaT24HbgmGuYggBREFu5ROwkM8cOftC
IOSjQ4/HorF9OURQPeOKhor78lakA9vrwNIVyTKTpquKEelwONWFSn4lV/BI3s++
3QgfVffV6628z3LAsFzQMCkivL1EIDKOFCL0hOzCxhV7Y8vy82Kteoi/4udzitSd
eafxlYUaBihvXzmsJXMGpzXHNs6t+qd+NN+M5abTmpoEj98RQF3T/2sL+g4+fMp4
mnE/mVP+ddQYHQ+jtfI3iQqWJjBkqHOroh1DRcbEKO5zuu5z8Y4w2RexW6jGqRt5
L3Xs2yDS/tnfWOtVPTYmuf6zpBbp6wIhepikbYnewWkC+4On+66j3FdLJaTvcJFE
lRAIOJWiJ5Has/KiHaUW+jU0vJVcCiWWLAfuBGVUQJZJsgOuZAeccyrbxF+5YpBl
uxL1TDX+3/ZVcFAaoQBlPv5jecFQHHjVEIoDZ49+vQIyESwdiPFMe2WdWsQXZX49
7DXTnLEW1SV3MauU+17srOtv3wP52H5hlSLq3BmttCRteGIfjG9rXyg5Ic+7NZi9
F7iyIUN/plPtLA8L6fK4aNb07YkXNzCrWNDKXEV4vBQilIQv4RVSEjnyelCiRAuP
flus9c44OgdU58Vchtdgzyj+rbgtPEcspGKDGvfl9qasGy2M4QVYuFBVtDNfbQx1
vBVZmZuGwuh/KxaRPDEKK3U9xpTVn/+9DY/1cl612ew0e6HGpTS0WsJgDVfip9M3
S1r0b4/68Z7UXphOEl3yVEI6uLrrcV/r/hn4/+igHbz2cskGAgQ5fwVDEA1IRJhU
2zCmyPbBlwDfrOsGVMFpkfNmGFpqbLwgXLXczknZ0PpPn0XMvhEq3nFcSqvCHbwJ
vDEaqzcVXUBf1a3PTX0TCOSv/Z8aVS+IlZ2V2Jn/PhuDKV/2GAYqNVFPAS4gKA3g
NAp6TEKdIAvRlWJ5tBz1zIdJqDiPZNtnvc27F4e85IqRgwye2FdyjQMgrq/ztDLM
UjhgtpamHxpP2oRgB8lLqfbodir0MMfq3LXmgp4prLKqKuG0iElfU2dq0ebRoqYl
qDHutt7svoVVpbiAW8DQdQJjOjxCP63iW/CKZ8c7+RlnvvioTiduj0aez931UVqZ
bIYaFP0H07pBUiEgs77xA3B7VhMquWFDacOXeOeqwugg/+i4Mtw4n1FxIMSY8RV6
z7et1IzGEUyvXR8TfYlIkc4huv3DGHa4wj4RaR8bA6/zJG+tDzPbRmrYS5w8FJUI
UW/CejVAL8JhqkAV0cHNvjan006g/gA3sKYGGgPB5QvkWrhNeLEjdYtpP7ilpB5N
Ok1FFXvJOPPRfkaaz56jUsLTeuzIk3rkpoHQtbM6yqM7W+uLGLoP6+H/1rfUSBot
USZIHLIfevVmWWqzbtCZiP/goqxPfCPUQsft9pDGLa6fPh7w9RBYjwbVhOKN7xqD
Al1KH3H9YeAaW9gpUkb15b+mZTajP7eGlK9pOjkxxzr1/ejW62uxqXRdL6oNJbfL
dfjR3ICHavYc+35iTHnmmamB6iTEPaxjkx3CUo01y0MJQh61o6Nf2DPrOuNJ7XIA
U0XAWJduWvZ6AmMWtIl9oC5fQipeQAUQFTd9V8X789gzXcgWofZ1Mpb6QQhxbpcu
0Npj6wrx7qXI/A80bfiereWYOg3EXDiOjvsoxq+jYy1R4J2Z56cGlMgndaeNeG+/
NPMX6jT0b3uyrTgooq9IqZlz+BSv+3wb6jc827Gfuoas1Uv/CJiuIFHFq72sqCrI
QCOe03DPHhVfwdc0odVDaHLWmFWCJVveeUss1wzxeVn8R+anux/Gq2AXivU1GRBf
BmWd+Po7oF2ACq4RNrI4Iy4PAMLg92p/ebBIrIdovFQIyfMsWtMe+S6wwKjTyCCK
xt0DTejO4gdHgweSePOAo/h2vl+bOj399wy2Zb6obEcL65U2xT4mjj3/q7DKI1On
msqSMM4LPwcx1p2nlAgYTcjFkMxZ2McD4zfvP99zySl/ZWKrUH8NweR7DHyy04nA
6gjr1MLlzS61z/A9+DM6aPcQL1Eg3eO2Ez4VBdgLWCIJakxG11sGDsdcpa92OZm1
D2UPmLSvBHI4r+X0xKzNPK4vHUQGZb0fsiLJ0J9y2Pk2YM977lPuWT0xutvSlGS9
nCn0E3WWTJYmKk5aSGn5Wg5DHKrkn9ItPIjMxpCmlUhdWyiG7Zax9lI49KLlzI3d
5GqEeStHpYL7LbtvsrVRuU02StRFdD0kdRjj4VrgLgTTp/zSJqqdSYJUY7drWQnd
AOY2t+LrL5wKzv5DjhvqzxMwbramUR6/79TN7YsFt5bXzzBZJvk+GwhdN44Bi39h
cWrkSsev3VNOut+p8xxD36BK6gb+gQUM8qSvOT+CNxp+/6e57unBnJx1hD4T5djQ
5SoUT5jyuWHkTDtnLq5grO+yPEQ8UcMrgO5neAzYosZ7iKxy9Fitz+5KHZxchq5a
1A3YT2OgwDrwAtvsxg1Z77xkDKfYQT8QSFIXjadejbQgCfTv3pmDoGReC7h1As15
id+BrIIgNj08XtV3+eUESRjqvqdf9kwFiMuvIywenHzwwTCiGFJzZz2tnZztMd+p
sSp/BdzZHd3HMCFET03k9GyrIlQn/dxGP7kxGEqZ88YfmFcog3OCUL7rF5ymLzGO
53ydtodC/Cl2ICohyH4hn5z4OsV/FB3+UpvU0G/3WqmHDTQ7MzsOG/7oEYoLuFoY
ZLUcSRIVXQf0vW4Ye7vCpxKlg7XSWUUo87/UNfZcKIBOarZQ7p7/jmF0oCe5ppvu
9wXrPFKeptruamEhWn+Li9XbiOWSQDynt+d2HucaNAPUw8EerW2Y9DTNqzgEHIZq
0A1XmwUfeTKn+AdjDUeNKKe6+C4wtB3QGof4MfLvoJPuwSeMVsHebf3tgIm6ahM4
PWCp8ia7C17tEyNEAcuJ4zKNIYAv3C8iR1ClQyywaybm6GAjbfnX0QroiEQbCSUh
ZDEOV640t0xn5PI0ppWtcOqbRbtPMThT0qhWiuPY05Odh33JH4rQF+fgpFZTSts+
/pQG58he+rwk6eUXswWNqNqRa1UvEhR4WXXn6u2FdJHzMXfSE5fQ3wawCIYbuqid
rhtWFRiGT+urxuDOnSy/4oJNXhwKeqq2L3UPWmpX130OUQiYMKp18zdpuI4cEsgq
LFCPhmKSMB5bPfndPNt+gl7cJ6KTaPqYOvOfidSjDNNNjhGMKlUhftJ00zRaOAbb
GVH8HPpqV/rAOdJ/lAmDAgVxs5kZzAOUHzRDcd8ZKX3bJGWvtHNZAC2tuLnptSXs
ABb/cTvskEdFvaAPKNeigC1heO1fE35Y+17JDRPhZP6K1yrg00rx8+WUAnQrgTgE
2UnKg+ibSbWoGSCqwTFon9g5XMRY+EZ7Z9ke+fC/cwoQdIyfSykSIfNyhZMhZFWQ
r4EemBqVPyPxMxXUjdKJAaTs9gcG8jrm0J7GJY/VtspHpPugBdSmzx90VAmEf3y7
N8GcH2juEpmk4DODA8YFlLx8esAJu1Ztd5v+061y0fYk/F7CDUAM6vUvbQour3jW
Z1HLGDYzJGq0e4H5kTVL5EH82IflbA5BDgx/dgOLoMnRt0Vf2lDWXeeW3G8eSHZB
bmOmN3aROz9vXg7N2lLyYVhvbu5t0+cl4FEfI0ZM68jLWQ+ewykklWZnhaHCNwBj
nWvSBI4DRLMyXfdScmZtMRz5EMM0vIog7MXlMn3/S28MsdUqL9s5srVcQJCZJ9mg
9sRxzqevq1A66FRh7FE8777RW3DOaJCI7Eqel5DYpQcJUHPhSbOumXDT4+sFrj/c
hiJ76yM7GT7b942QeqjXPgjd7Nf7SUV2mT8/w8wA7vwgEoyuImCjtz9yQKNF6G3i
QK+C7pgoubDX21Q2ekjtmO7p11t6yEdHVFAZlP0r5tVa1HZrLbuLy6W0cB0Ax/+I
RgMDfO0e79lFka0GeXYPaju/++PRYYiBMn1woqEnWC1+pSCKwkoDkfd60Mc8EZmh
ZTnLvezWyKKU3ma+PgdUaSib5m13AvKm9s6Ewf9RW5HBfaXIhT1fJAKU3tk6Z0qr
7ZUWVd5SM0XpoQG1BH4KnKqmFbsdqxb8pe8VZZhlmuCnIJkdRP+eZgEZ4gyTtI+d
gmiDhqwS8LeliHZynxLwQCc/Yk80Fuh3KdfVTysJ9V7x8oYF1u1CeU3xlV2qdGgS
RhsLPafxv8Y3NpOg19nLFf7oVKT+o/xVfrn2xGhWeXt+YwlZLRXFoTGlp31s91U5
3MIzF0ENxXFp+tz37ySltfZMd5Iq3Zz+AYFgVvZh76PqvzkCsOTmuqHLh5Ch1qx2
6YOY1B92Pv+L/RWBJNxIgcICNEaeAcmeY5cl857ol/szsLUSOIBXkrNBqGDYzFkE
PX87VP8Zow8SAP6gh8ttcy5STwo5A+ebkY1AqRX3CpxBoF7okalFrz3jtTfqcJQ8
Y5docpNn5eLoM0DA2I4QL63e76zclQqNEGeRKOPQ3SkfTKsIhc1XAhcQ9SfHhFxa
LkD7AHgrUK+feFTXqkxcvnUwnS5ggT9qDfeOob2wKfFiDwnfpw+37/TlY8yH4Rl0
oGFg4Sjq+FVAsJg7XKwFBH2EwmXLGY05SED6V/EAK++HgbhMCk8YhEIArY07vAng
F1PPtwS7cCMr/QP1WEG4BjDM1ebmSMamHc0BONELJ9qT0KSiFmgoMFZRBlS65Uex
6HzVgJRuvFvrc10uzqdW4zGHU/MJ2TKGx8cLQQ/RI+ToEkJpzvlX2CeFp/1XQ3/w
/0Li7CieJfaAHzU3jhix3FyzZ/bpLjepB4KFDk1nGjFEn7sCviunvp2iALSgLpFd
W0Cw88IB3xWp61gvlxxqxaWqyXROC+qpx86FZJOVzZ9aynU4a0TWVW8eiksPKUiF
1Y3di14gJpCQdOtONxEuYa31VardPzf94C1SoIlYcmPFPjWTqvJ9H7SXeatVaJp/
idcq/AUJuGTp1YALMuUItn3zfwp6nRUR0T8xJnaOCkvRYJ0pwgWaOH+WZfEniCJU
qPHMnkti9CBgzMZRqBeyHgKSMO//p3ZrIkQHm5SoB9HlUCuC3F0ECTstuGUwdcCD
W/7v3sTJbZCpLKoLuJk9DSCaQwbSK6iq1b19PZKtsMQt5FGV9z8tdZQK1zm6ySnF
OPcMUVHQzQMyGfDqorbdvR7P9tSNaDKszEH67DsTlRcjBShbPUaFhJLPTtYND/6i
3YqgK+cgQeYZyuH07YtB8J9QgdFfN97VY12mM67aqd7agENMmxXBpCGCIqDE0XUJ
6Uhbjhd6LZTCK5xBpTAHsYs7YoPMS4XltGT1GEWiDsYu5ES2zz9YLl1sh5TBkA0m
rhymrVOfdeYBPff5cogVQ91Klb5QMeVc6zm1TT3NxJJ9YjmGhsrCU2dGiUg+ENEe
xw0dTCWCIUMVMp4nCbh536s7941SGLLAPJOwFw3l1vNY47WsYZ4d2Nx6+XBRgv+N
BkSdlBJke42v9xUEbhpCetV1HSjFVUkjX5HEM1rOahTVyoAUMK7tqdUKte5OiN1M
LGobYpBf5nRYJUbh+AVNv9uu+cnZhJ1Pg93zlM4n3cOGcBsJvZHcuIziP0oDKguX
2cUzdD+IT7M/K0Pesxc9RRckXuH9RSPYyzWAeAhldgvs6IY68gYTZTShBHLb5AQq
su+ZbVX0ZAZsAsrsfVxAjHuAzpdh+JMQIudaqzTl55Hl4kK+EC/qEF3vzaHAdApU
s5CGiatJDf+6YMKw+0k0gp3/i56N+GZrMLRzUyoSCYEHH71PAyFblbVW/As9PQ7h
aynHcxmklZB+Cf/7eZUSy/VLDIijwHp0935Xuci2KAcUlZeMCdSmDSxgCxxWBc7i
kWP38zPq+Ypbu4W7l/dml3XYZQRRKFwgboA0AR8FT4VJ1ntCWKgMBzlkjw33/mC1
4mBnl1KVu6/ktYRrDdnsGojFQBAK94fDAVQ/dosCbizKafL0s60+GrvBa4jJfdBJ
RMGst+YBNhXrIRare0rUHlWgFeFOFNF0jPONc9debpSHhqOA/DVaZ21tFLM23G+s
yS+VI1qYrT48OdFjbW/8S0gZIVT/sDOREjPj2f2UncjHXopQAgW2V98d+HiLSYYu
wK972cFWweym345C1HCnGrN1irmDwYitHyUPaJG9SCC+/aucYuui8pFXzZXlESGK
lkA1iRLIUOdM5tv8We1DA9XkX+6OrxF7OV7XXlbyHuubfyAfSM11Y/rdfcus6HZV
HWY21hY82pzQqmFviMGMTriAbjTQ58lWbca2CzyNkm3P7Y7iHgiiiDpOFb99y4eD
cafN7dwyn1bGxi+GPaMHFMzlWV9QAQqN11epMyvs+MJvjI8j9NNpCq9lWozX1mtP
70WwLpvhjjFO0aDQ8QYJXzw5HxBWxLJ5VhcXhHC00bXLrgQDvOt2B1ZGg2of/+Lg
nfOWwBYgjboe/bGOBmOF+aVw2regUJ342RslyUmp4vWv54yHWiyPc9JZzczle75M
JoBGlYy46s08A3Ii3ExhBHS9uERKFcd5dhIKwjBSpAbpRszz41rS54/DcoPWMlAw
6Mo0VlTn2CdkRthE6Eh4d8++KGAOgE1wL/K/So17+dv5D/zk/G/4ZVp1Z3++Ylpm
Q+VWHUJmqX+jOrPbeQZvaf3hTRSPLEhCyKDAiLAA0ofM+ujgMyDZoIQtfpQdO3dZ
u84UlpH76NvsxYnqqeM2ANDok13mfyLhevQzANKqm47I8N9urntPv5rELLdvwimx
QJGS0C1AUKJRy/i2qjRU6kOc7XlY2NyysyEPJZdM3/XQMrAKg/wv54R8m3jJezLc
u14N1Ha8fhzYZ5kvsKhbS7lCUKJPAUZhgIg4kAx7cU0R+7/8Wqb2CJl+iBAFgLxD
U+C+IqnUD0R6FJLH1FJPObxi0SFBEqG4VtsOE7NPpvsDIBvi8lRHCvUl4mPPD8K0
PWLIYR7tysPUw5diLW9CONG8jlW5AYqErlZ6ahUeyGsM2TkOgiVl54dA+0fbWyBG
ez+FS8gT9uFLxF9oyEHRI9VVPlgF+Yr/LZb3gHMXEsULE5UTyixULb10XptBYVRB
6x7bTNg7vs5IMYzPEWfEQNAdPulBDX8yQXJJD/JXh31nPPnWh5FTSpG5/zOPQwJe
U9VsujnH5mIX95brt6Q0vV+QKbGy8g+8abmZ45bB8pCRW3DOdCTn/WWOJZeK3X+O
4mz5Re6PZ3SnI3qIFR6mF/IyLH37uYK27F88FaJTpoZFeQBDCp4j2A8zX94NLgYc
b+Gno4IfpNjoglfp/YUNHw7pvIpf2VpETcLHzrnE9efHYDapropJLnci4Fte1x6B
kown3za33gOKKzIeRgcQaGpFUvIef/qP1NaAdETAHioz4LY92r6X7IJ9oewM0yTm
jgqEi0TWc0Mp0RoXwZpFr8halaRfPevarR3d0zgx1z8eYWXuvaTcxZj+u/EG3gHE
DNi4hkjhst2nP2M5OfvgHOzWuZZFHkxqdW7pf6dUxOBfBuqy586LUHJzbKkymHwM
zQJXj6qqw0sKL3Dxb0r8/gEOOdIzLFqSwJ7lP0qgXICn2/HCuwB/vVy6bbBWIHfU
+Cfl2l0jyvrKOVFn77Oc3TYvGhTlH1snZoeysc3Ep3xbK2d29Fa2uzGI8+SfMbYV
JPOdw+unrtSXYg9+WNVmxMAj9l7MEUCUELblIUgeTKSsd/CJqb7aIudsJIq4vVPm
CTAT+qb4Gi2kZcKv0LSbhDUKiyVBncg8JM/lxMyw9L2sj4QfDf807Rjqa7fDi73Z
CyORQDHd5vXfsnkvOPujvulE32GaYHyKsYLoeR6qvJbBP44dfOStK51IMjXYZjS8
C4knBuu/Dp14PLhBV7lHvS6hySErdSS7iSUg0ZGLqrtA6TSU69NYQ8G2nf5VMjQc
fT/oT3AXnEgX5HXtZIK9jjn7Op77nVo50hphGxGCT0CcLHjH+pcYCYqbVMFthwpG
sxQQq0bk78zGWTIEzqWsbrZFhA6rxV3lRwg6fsQmU6VU/iWrWNHQrw99iI6b6vRx
Q1LL10rWCAKxexUy8SIxW9byToRj2/CYxjitL05dfQTvpaUqdtOnAiRHwHGIl5Er
X6/PWPua6n5Zk9tsukpf7wNhgymyEZEOteRUo+TKMgaHg95XOdOyihHDucj0MYQk
EObhXwgbHJSO2QG1p8xSJXXjs03Q+j7CRakhoDSQuACK6IZmD+JKsrk01FIA8jBX
CCauk+6LODHfUFJK/Xq8h0/IpdSObocAerqmy4Gs20ETFRPHaGQs1TiKDGA6Zbdl
lzbY5bg+FX4WOPqAm+mR57jQO8timh2YpXXouOxkNcwgMMT6KObd/qQbZoEHai1S
Oh7vrezaOv09Jxxwa7Q7RGOxt2diwSX9/eShDXjBpKRXguqXc6iuG/cBUYTM1nmh
KvGK9366S99kMI1+IRE7tpACyUISUZdMESZYQ4YdymZNixvp1yFRzRRW3QWTivJ6
QB0cXb0XHmTALZWuHZ7+NxZitmit/H6aZ0ZLGAZY77kPYxW9eC+2uk+QPHcyh5dv
uclb7RECHAQqY3iye8QZruKmhm8wGDQx6eZVPlkin84Igg6ap29MN/x58jZXJxCI
L+1Uhcg15MTmKFROV9bvjo5C+qmUobTLUEHnZ+fqAzQ7hsMUOuhxsE5MtV0OgRzF
fPlUvcUdfUQagV/UKk75TWi0UpmN4kTyvTDj26+JV8Mf0zAxxYqZHeicWQ9GlgM5
j6ai5HDqWlJNNqxDGL/usTjZIsMcaJ/XAN69Sk+nSQC+ZJtJQ1/CHmYWL3vatPpb
Nd/T0BvmEOfvdL1gVbJ/QJtCAHOEXk0okLBorYBGubE1ntiex1n0izd5KrwOTHYw
j8WcAWU9M9+7Vw3iKW7rCXy0GXhLVgthZtFiQOJAXTk0UT7nLgkta53lY+kbubmh
ixmJFhF831LHVdoy00UhGg9QI9teHx/jvOw6zzg8NC4UWBIVCuqqARcOrxTyCLot
/6/aV3JrjPg+U8nhpqAxP4YmbLNrA9kUdCxRBQm+DeD1yOyz69Hsk4MjpVrnH57X
qWg078KIE3j1b4wZdJJjLApOfigimzqzmV5gLjiwEPVUvP39VWmJlAH0OcJL4dbL
zQ3nTOkHt3biIhl1N4Su3kxpBADG55YoDb5J6wRkY6tOnYqn2MsPZIszBrSridn9
rnotFP2gp9T3Ec/ED2DAz7znNk3jpE0ERGnH3rZLKxN805pHGqNjAx6iCrQTbEZ0
ablL0P+g72QDNS5UXfUhKJA61vS7IwE4ViOawW53oUYiVxRWxLob5h6a4gU5MecB
rud0nGCsvwWQ9FGjvySPMEgD9GY8tew0tTpMfZ+ipxdbzdvCFuMIbao6rr7AxEdn
448qGdsgWxDtSq0h0fnme1MafQAA4njCwChUwqXhaGfwg+irKuQ9sPf2I64pIxoI
Dg3PZkVMFFA+gfF6w0shn9wo/wsfG+b+xjGalYTcv5vSNoF05SlABXIvEANDFB6n
umE6nNhECbLMk41ZxKl/7TntPfWudjKHtkyE9VtWYFvtKlUTBZFs+FJyY4OYyr9p
gOKept82ZtEP3K40VKVXRM5hUBH43A3sMT68Ifkv7l1/1qCWTHBpwEZ2puDg0f+d
LGDOPO3Y0B/xI/JocboVABXbteJJ9nqX4pagvcql1RdkY54vfc7LxzWmkPeBj/ON
SMC1xAP2C+LDQeFHdfxrwoqiFYAwmxfBg2PXC+OX3TrbFHpzN123XBcrQhcti4p4
G+KHfT03JAi69iCMz897mTQdMKIJUXJG3cikwPC+4SqQ1RMcWVmYhASCjZnYsUsr
UJGhKDQpgT0hfGq45zn50rIOecmpAEuvb7jId+1kxT9Jl1iOg3P+VMdkR6iMOzLe
loI2Nw6AW6/luNXDhqNQf9wLpQc9csyIqDyGomJZiATU9RSUJTEfQJzFCPCQKlZ9
K+YSbq6Jnag58Hc/n1xmB154CAcNcbJ/Egq1Pmmvyptlf9as1pcQANjloZs4fUzq
9PXIBLmdHxIPM8sBpG40jcXLUVtAkdvsAZ6fD/mHga3REgmETvHA3gfFpe6AIVDQ
9Z6/RPVJXpUBTppyEc1gwe9mKtgYCmc9OeX2pqhm60s0sXnptZF8lXsG4TDjRK3i
yGKgPbnRPMifyCBaKeqlkAilOWTAa1obfiiihJnXYc9oS8eADqutHnTpGZRDgvCW
RU/JqEIvQ3vPOQ62r6OPXQJaTMMqmhs+bN77qM/vOBIa3MetNUAkWM3bsPnjXFep
0y4ti2tZt3XObg86gPAWm44SpOAJMdQgnija8Shs3ucxzjJcjsHw2Oc3rnKdyAtz
Bwusbh4RMGSU1bVUlqhIExfQDxAwgvyXR6iiw3C43Lqw8B+zmMe8UivgU7H+1HW1
urqvHSWrzPwMV5DpyfNIx3xngKlJ4a4zZHGuBTG+l8/tTepm9aK9h4oPSluIbjgy
mqv2xxVm+7rVuqnC7h9s7dO9tUMMLJhCbEno5rv/HXZoLtf4CQzDrj3O0GQUg/Sm
Ss+C4n9y+JkWSFjvrWcG2TFnrsxZEoQQITmNdVHKdLZJvP6e4CqNlHUX0NEH4WIH
VScGtn5BMu4kL0DV7p21qCxbdplMxQ/sQ7qq78u9B/0gJU7Ol/iaK5A5BkFAhxre
cd72kz5LTiRlVQzs74uLEka92+M3OrEMUeForcFVr+68oXwMaw4akrPqAvfHr9XO
64PG9NtdlG/IG0N69Wgtn5Wd1eG14Yvy5TEfQ0UzbuD6bR2Ep9JfC96Z3j/mfMFL
BqhTzhz3oyfPxBKDqYVvR30sjNBBUn7UucOUqtFffbn47cU905J0PlqfWjsIhHLm
frc1cinMqGoT2C1sXhf1PV6oVKU4vyD5Xvy5Aup+TIPRTdvZmDshTMBvlEeP+gTm
YPqaOza9q7+AFGE2rANDTFPruR60b89W9rcZe/VpEUzzSIK5AfxwrnY/Az0cC30o
PSy6oHqKoQPVV0WBnnuVVh6idmZ4AGLKshFmorkjLfbzP4w7knKzzsEdn6z1xnk1
MQef/B8szhRo1YYlIC6HXDpIe6bCCCyG9Yn8CsAYxeAfbX/4wv8eAXfmroa3V2MO
hpzLX+6e2d1cl+CX3ReeanMzrD9roUoPvd86bRPX/oqLvrb+gcBYCYMx8iqT/qjb
k1MZJPTLoEDnhaBuiHAfGl88HPxgbEMlu1ITbv1WinAunT5eWByQ6xClEPXjkx0T
zXbICmnxvNPLJnqSXeXHu9txbkQlzB2AqhaUos6vT6BqFxrushmceU5yCGLai16Y
Cx1A6Kym0LJm57BpeSnwdMeGlL6NOXVKMgGl2z3+dLOyggRlN/fJesDskm7oo3vE
0+GqFtKmgyepUqZ/Ib/AfhJbCxjFpbMkadYxN1NT1gcZjLkBpa1mHsbLcrRfD+yb
dy/TNR+T/PTyXRzz40oF9wSPdWvhMNvhBvurqmTEY4cOKWFEOuk05pNdcJSlfE8t
SFrKMK4MVifoB744KlAeYAYjm7HHDJAi2mPESoc+kFNC1YcVf4noG4eyTjHRlmQ+
ZBLuo3PVX1dXKY+R4UIDfyhTEXKUBLhGxHhjluje1UxITOytuSMrNZvgOvK2MyIG
mUyj9vnHmkqU/4XuxkWjclGsGWqQ7F+fOTItwNssEpjmeu2M4SQcfykVmmwNnXkU
abdV3qvaQ1f85hBMve84MypABB35gKWljH9tdftRlvu3v0him7H6nKdNcdJMd0rR
pFQLIbnb5k3jNKWAy8L7MAJJylCWDqiNUS13tPHgOo3+rlGhPEa6FiiVvWehgMmk
/TMd3wnROgY6kBLLm2JGrzBS+quXIL3E993m4mh0zEhHG1OXT4j2za/h30g5Hit6
X4zMMx1Ycx1RzREv8EiCjn8VSARpHfvbtt8CRe5uxUY3mPswHUS+uvUj0ebm5Tq1
wIrKVlny5oebNPw5vqel59KEpGH4/pFgNhp0NiifOiyOvV10JsUVtTepOeuKsPAT
RwO057le47vnulYp9uTaHz9nDA+J8ZteKp0vInk7mFX9pAPTbNnGkwU5IcHQx8dS
Y6rK9Z148+e0+8LmzJ/0K0CMZ2C6ZfX23O/qK0s+OgV5s1ZdAJ7MjdI3PCdM2HOh
3fpoLIHm6BpZ0ZiA+VkeVBSOxdTQEkCkPVkbpakMM2rXVBX7UFXk8fpygRiHNkZn
vPtnVSHC8MTyw9qXkm7wt4KgK3L0DS2ax6iLorJFIBSYza2aXfxOecn1cblRpA9Y
YENuylg2oc6uy6VNxbEJra38/Ir3AwIEvoSwJD0lgJcjq+QFY5JG+dqUVDxTRLBI
artZ1WXZ+ZnIGL/MX8DHpgKh6w/U6ayPfoeo0//lRk/G2XMpoU5RslrC8rxEn3F/
lQoSJjt6L5+WwMbFFQShCFChpyWOPQq+TcDlTrRT/f5dpoXEkmh++Cr03GS05kWy
3jyFn55le6eKU+SfY23SmXbA1kjVqOybuwYgaMCBaWxgwJjsiisLqU4g+1rkH1Ox
/Cq8NS6BOjewFTAi1zVhGjaa0NRRmQSwKOb6neeBpmLX8KTkF+gY28uLq9yCuciu
nriyXUfF6eNTHzr7VaGn9iM4hCjma2qw0DtdI4L2LiQpJopFvTAQ4G+EvxtzxG0C
hYwtWOanZgyW5ngHh6Zj/Nx81giPVS2n1NWHrlQEiuvWKgXY9nO8AgJWUtHaWLqD
jrqI8JzHuvGq+EZV/Pta7hl7BuOQkfpEUv5WS1sz47/hvjuFHh/XHdocpeWSlh7a
IXaJJ9ZSU17CvXRr+/0Q+WOSinaSKDijWSsrx2c5m5ykjQOPxJ97uBTqHQh4vC8t
PdfznQyJv/TovY7N83JQlXVm49SEM4cynHJV4t/w+jLAtaU+DMGzjxn+XY+L++3n
C70QRyQt82sIHL9nJxV0MbXlH0A5nvbBYbbkYBLqLZnVF7bslqO19c63Dea/vOeg
opY/RHDqV31nhuwh9TFn1OEgmGFOaKQZnDTwbZaO1fe5xEBXIADfcyRpFVuPdPny
JE0zIQ/qVDtPSweI9NT9SrXJduqtQcLH6eQ2SsBvxvwWq+xUh0QD0uvE0tzXZ0wS
0VKr5KiBGjoqtgttGPmDj4V6BVc+Lzz4Nu2nJzOVK6BjgZIzY/iUi+8poYNmZVwg
nq4beWm8Gi+iK2jFWJ9XJ5WpiSNqsJ98o3ZGgUPrB4CCGmLkwsl+dHt8xXeft3tY
d6SrkKkBWOWB01V8joulvdVFy/lG/NArGC62tz1hBztjFTwTVGypg6OXfwHCohdn
Bq9Md1gPsL+mtG0Q1CeZI9nIJoQp/KSgKqBPdwE14wpdFuJ12TSqoRFlFmKamWpo
R72RKD/Y4UaP/3h3n+EGbs7JycYNMm1KKLZ69p0/6/RDpD8OidX3Oo2g0SUzKFxA
Hqmzb/oFrkenmpuBhwWELG6R/Qowtgz2knNW1i6pwRTiA4YN297p+0JtwO2DPVXX
VT2e6pb7qBFORbUuVe7cAkz+CI4U8NiglTTCIC08xScjM9fE48DUzMLSRfv38vtu
kMmoxrlU2AeVMDqScSUDB4OJGudW3u5NQajXtgMHd4Mprmj30Rz346PYZoFM7ktv
SvXZD5PyGh7lRbthJaYe4fStTOY3IRhFNyUg3ytHBX6OlehRKH97ahtR0/qdAyLp
f9khWxPCB1NcTG4qmNYDHvimJ6eJVA4n0sK5b4Jjseryj7fGwZbvfteN8h9SC8Az
nQoLis+3Cm+cpkTOH96WAV74ulcdxpUaxERAlx/AtAn5bbi0PP8ei+V3u97smFtJ
XbX8sq3ZOMYHoUMFYWNDv3qeQvNN96o2aP1msXxcHpRPSGHD/aI11KbZZdwo/ZAW
q/7lUMXHWYXFNdyN1R50Ge/er4kANfF63SRSsnw07c8xjjXB6xseBVIHeMjSqhdZ
aIapHljsa5DBmikYh/A8W2veW2XmrliBO8xSZy0RqbBPbL4lXeKPWb8+x6ZmLXsr
balPmsxlncf44ZXrCe+PWO5LX134WLZ1/60Ix0eSCwkYFZNghZkDqwE/v0SsnFUm
NyKPI3jJeFzWyLwtKx80B/tpDvshAtqVzDtf40pThoipahdT36Ctz9laAY9OVYK3
zP3BtkEdhxl/J/tUU4XQyznS39oDyj0eouF1mZ7gA8t5/M//Q7S2RfzHByIdgGyG
7mc7ODUFAayUgIz8wKdSQiMYUhcrIglqsAqOuJ9mefmU5AbO9Cq2Gx+GA0Q0F2l/
WeLpZuqVv1SwicqLHxnkKycZxN3la36XG114WRng5/DndSFpCQgpc1UynrC+H1T4
pGd/32WxPpWXA8UYt2NQyuBfW9TffjTRyag4nHr3jX6h9FvBJzAe3D8V8GrnBu6D
pP40XTvyW8on7fiiHQsCZUOC5qHF2R6M8mBh6Wj+SMhSJzUHRF1uYjiauB2rdkoz
qOYl8jrf+71UD6mYEyhqFfHOmSQ/bfMvZRxqesDKaOOnVqkSzNvOvDnZECiUGP7c
OFUqetqu6OyBtJExmyb4JuOCdGEeMHzKaCFd5pYByg3Z1psdKTV+CYSPQbH18qsj
+2tpoxTbdlXidFFnBudnh13K2HcDjmRZ+Ecj1N4fqwcyCcKS8cvXu4OHOAGEomQl
DB5SmRVGW91u64rrrQzwLFccUssVgZZqAjao8RmJAMUvVdHDdZkYQerhvg/pWJ4D
jUXP+dL+DHRqJXOwsb1suJcr6dJwxs3Q0B9PXGSPF8PFgRKxpv7bDGtMxW2nE2X3
c1k2+0dIVI6EZDvUxTBbpDH9NjZrDAWq6fgvgVtoZe4qNquqvFhd1l9QCVF7//6u
RIaC/sPBv6vV7P+fdpTCtU6Ug5R3mcRpLe689hSGfe4lkOBtC9kM0Oq/99/4cChl
pxNeKcyb0Q9AtowkSZvfREUFgERVhFrDzfH8F8HfZcIHUL8/aVTwV8eHasV7kzqh
Y7/Qe8UPSBZXPXt0oK9MmHLZJr4rt3G6FUka5fJZtYTMK09ZrboyHMaqs1mbCTHi
2VaTH/azFueViP/BRzfC44vJTVHtf7MiHAp0OLWa9nHIyS3n4r/K2LixNWHUpgO8
jtLzi15A4mn2RDnYFzB3JymDl+3cWu47nvJb2vMw0+b2YnzH6p8VJrin2aLQ3qVw
OCNsji3obu3joAUPxfcjOVOnYNYdaiCmuwNT8gqI+i1CVgPUZqpDL16wPoXAuts2
UxdHg6KtGY6OJxplCqZsdYsbc8Nr5wlHU9Gh2y2sEKsczui7G5HZodw2TBzFvbNN
3H5S1305/U2eNP6vZ4aobxetAdFxxWeu0PMHt4kIuwn7hNnw+64G2VoHoF8gS5Hv
SZgRqOpNFAPIExhTI6QqNjtekyJPjFIIfCSNJp9GKNdYY0w/mll8bVmhhfrPRXiM
hRFxONHe0sA/RBucUPm2YkIDt7vteHgu0CNG+r+k0tzziqPs1NTiIF52hoqdr7hm
Pykqf7mj8R1Q+N6BFVh++xjpkT7gpY6RScDcrOBY7FxqBb4kCA13X+G1rL1xyFEu
lXXq0BkDmFrwEkGy5JFYp8F4PfaHFPinRy1v7kYHrnBRWLaDICCrVE6HfajKJ2cz
nLGUED9H2nJQQtH4CN3qXqUoIjZY1qiNKsNHWlUJvmsEtnPUaFD+Tqzjk/LGUM5F
dq1lJskhWoAG2Ky7Wzw9kXAjzpswP/WNBrnZY1z6N1mP9YdLyg991VjWAtonNCGn
G9COsazJaFheZZBzSbqp008gKlI6H6qKfTPZ/qAOoosFnPkf0XRuqOExAdj56Exs
oOC8fIuZhVj9la8zUgWi6Py6SUHAnCt/v8/oZteeugitdj1xO/p6EwiMvRdQQs/z
Th38tK7KXkKvXJDjYjVhbTI7gOFOmeO5lcIxuLFQ8OEC4Cxs/lmJg5tbj8oj63iF
B9YvewL+FuQNVonrNqtZO4BMhqe8yCCqmgKcoWMx0R+15Gk+al/ZiHmTRgsOhnfb
1ZRFGfRNdnN3iduJqhnUf2j2I3P2uAps+my8fOnXsjW0KRK4U3puWlEw0AYHfGit
nUJMwdeCTIg58nhzFNINiSXf7BQHy0V0vn8w31fplu1P9vke9oC3gS6J/xf7MFfq
FYfqibV18AP2Pa/VX2OANccozTUU6Y0DUWguiRaaFwd6vh7ppLv6N0P1jrhWNo09
iDOdTEB27arHohhvtlAc84oKq9Xmfj3X78nsEcBOVX1t/Hqzi6k3oN8jO68AlodK
szCNC7zkUdyjWdmyOlfkByB8y6vQWzL1f7oEPYUJP+tJPJGu0EboXh3baHbvHp/E
OMugWcHtKZF/AoylT3DHL/iHm4atNyd6vUog84TBZ3MkkguFR9k+GqID3ZGEP7So
QoxV6aCE/lyb3CFQwjurWMvvLhnqYHIvyOb3LfMi6M7I+JZuq9fus5akIlCm2FeD
9qWrd6KvrZoudJFTvRg3mcWPe9YHziCiRiH2VXJe+/ZF1XAqNpwycZznbgMiYPLT
+Ahr6ohusD246GQhDAKeknv4Zb5g0nPEJYCB16H9EFYliCpsaDm8ZPoH07m4wWJ4
01vS1lSmo84zRJ6y9hCOrcci6JyVm+0GZNLnz38W661FUANQ1jycMJ8wfj6ECJ0+
ohGrV9U84oVPTOQmp/SGislC9PbNQ9/fL2TJ1SMLhgTXiHz8X8CXNtN2SNCja3z+
xesC2zh6AvEItAZVb8fu4J14EoEZJ1OqX84rzlXKlYwOzNbCICRSohUkQs+xfXnR
MqZA9Qaw3tMhi8agZ5vR6nEgZLv6PkNZ4ET2Rb2H+CSyzInR/tDZWycJ7xfFs/zx
jP94fvKTQBkSHb+BHuc+s9HInL9xNeeVlAUoer9SYBuCoKKcX2bVw8CR5AFQ+XLp
cYDlNQhJcoZxzWXpUFJYhv0AQ0jxg+G9yBEPJ8Uzi89hyMvHczWJmbb1XSwlVRL1
LanCQy82PabNVKWpaN3yHDU5ymHAXOCI4jrlf6K8PtIQXEOAmNGgWDo0C5vy5MLc
D4DQriZ4kj2/zYYz7ysgEuTb1bkdpZZIJYSgWdLjShlAjn4BubVpNvaLry7QdIql
U2lBTyCyr3RhWuDri6auRAUWAVQWF7Qt9Gv6RrUo02Siniy01+bLcGXKbdNVOzB8
LOHVI87kssDH5D4mnDknqRApYR93RFX3vsTsFKAaV3QsKLT5MItVnbIuZ21VZdzt
s09zS5G4uIJhjx5uQjxJKPECQJ/LtqazWjuTH5LJAMuytUKSDaNJNvhwyBdFmjVX
wuYlhU5PKa0bo8XP0hZ8q7BQ7h7qRXBQMn97ZtNqcsmMfvw/jquTOhlJ9tZfogB5
uMXKvt5fxqlnj2/fI6TyAE8ZlV2Wjks0lXbGWcPM2fdxzk5TpPLFh1vC9S1SKZxf
WejdIVQ24cESTgchGOIcykQsLCa6c5spEiLJsZFO8mdDCSiN/CgNlT25V9V5+D0f
9XTbLIQZCfXLObFiRO7wtj7J62GkzvMgvFPTHEU8kT/DQYmM6Cw3L+9a6e0MnAD9
RaLzbhXFKfoiyspSA9DK8E24f6KtGawBqOBmdtG4Wo95AVTFEFdrcjAdODxZxEHo
JVwCb1j9XQsb6/oO9vwkrCYfECn+E/zBF85a4RYr4tQse/cF5PbE6NWXk3yf67i0
Hik0mKA52sIQw02oYQgCIcpBqNS3E+MEqBOgRvKG7WblpMVo1LkV7moRoTwZGaQM
LoYYT/tfJocMU2opUeQUe6wSZD3hqtHRI2awe0worFudvhdazJR+fmbNBzlkeyuc
/vqXdIf5Qa6rje5yR6E54NVXar4opbSeA8CJe7hKl2tCB6HfxqbRqhRSgq86eiNJ
KMavuUkfH6ZENWF34UwY8+c8iqD1EkBoA4WRBfKH9SfGlBuwJnmHp297Jcg2RI/q
gZyAr1nr0qJbXw1U/49Pw02kdtD/lzuEbAxzBD7avl5lPrt5QXzoGVEm0olSbB4J
ExY7qypjyXhK2DXpeweRGwg/Ao0rm/iIsyQgNcVrvsvvTqxkOMC+wr08EaqNReDl
twRHPrViOmHtibFKT5gboluc9ZkD6e71j+VTALF5+RvsXmtCq2ZLPJYlumoutT6F
b6P3spoCSKWAi6PHG4cljbNUtf3Gcr11QmgVEHNhgPxQpswxa9MHXC6fVGYJy2Ez
m2v2zgl8VwIgBrBSFdCbIgEZ117T7NnXGpd55FxwKgAijCJV3YZaR7VCR5T/3CB9
Fihsua4HUbrlCaJmTzNVxScqc/7ZKGE7M/3vSer7Bbw+Kc8YwD+30KMNprWbS5gU
hRSp4kB3J63pFS47YUIeu8EXt1ewuMUJ/pFKYYVAVVUxnKnHtL6WZephSDPGTJNm
xdwgoox4lqDSCr2ioa4HZ2RNzoJnTeoVIE90Sf0Rf9EapXMYr1QocYzMW9J/34gR
enHLVnsDaW4ojbUjfAx0CSxN+joOeOF6bC+AuM5iom1WrL4fnwlpi5detAbVG+CB
bxT1rzYmWQEQ5XenObqGcqBSFr8FzC3hoD74KyhBZikp4sjVHyWRIQyhirRD5+dL
MFcOg7w5TpF9r1zRVqJvk7sd5AI03XQqdB306KnrmK68tesogy08LOdQHZXWRJN5
Fh3ZNO4wRGpyPeUjuss7KHs7tXOADcQrEeaGjcCJ416HWXXypuxuZyDf9EbLTASh
n6VpoOM4A5Sm52OUJKYy/sgL+M/WWyQSTsI/Jh2o0KgSiUv8dpsm3sSQuXnvKxfe
UN/jV5rrXYG/AkByyYM/Y2lS77OOaMXOQ7CFTjKQzf97q5y8Tu7RKsA6IfeD9DS4
ykryIeVLswI5vYY9Ps4kbJuANAJlqCT8LTM0YRr8LGb9WnCTEgljY6arKUTa8SXc
bXb9ffBXB3LKJFm0ttYl4ILGiqzo5+w1zqMslCIhVCKlHgHrrX6s2nv5gkeYwJDJ
btBcfta7JrZCxLDpy9YNF+igF7ZvkfX+kW7+LdPQuKM7czJyNe0/EETJwqKWO+fd
Wy8g3EO52KQTx1hhf7Uz1uU5U+BcB0JE3X0yqY7w2oOTqMcaAH+LTzWWxe1DDIvU
mq3Z2oNKgJkFSoBTiIaOImGSOCepnD2vLLsz/KuX3kPdhIJ8KCLJpnesfSDcwxYw
yc4qNttq9GAeLqDEBkDGsYi8BHvFpreEgnBczaAmyHHKCq8lyAj/aU5L+VLCEmJX
Pg3BKgGpOicY6+e+N5fbio7jFZWRMgNqYHxTMRvLQzu+5/6Bqf42S2ijZdBUYp9P
fAn7yY23ACJe4aBNAzzhM53QxF7Ys5vBHqM8LyMy880k/Br/JcL4kTvuzZQDXsLm
1p1RkfoM3hX1ogEZJGybN7bRYdWNGvnnSGPwuvnPyrvlA8ZGNOtG64q26N8sDNs8
j+b+BOdbBotXjusJwuu8w35dxeKDuA15H1Parv7nfIsoWD6/oto0xCSUpXiG5yjT
dx6iOYW4vGKeu2VVgzMBV3dDjjatnfsgcerznSZWT+Ex5yQNZ5D7hCUpB5/ca908
xweJZ6Bj2W0S+6ActETMnAfafALEp0e8i6pOZVE5xriTERZt0Gpv8iaximW13LNW
aBA8kGpUjCWgXzVfI3/REumM/o9lADEmhEtbNrpncFGHCpjpEuhgrlEJ+CRnAWRl
FOzBzVsAeZAZFrvsGZyWd4LpspIY6VXK3MJprTYRoxwxEbUIFYnw+cswO0x959Ps
DWAcznk0/2UcRjpPI3uGmbwPk55zLdx75YfTJT3hIAy+lEJ1WldYR+1Ho8dFk6mH
Ihc4TxzpAk2ynn3DRylCrnTHMuUDPrV3F7dn6cAX5mDb0Gk6yRNciSFnolp0TU/w
zf1EYGf7MJkxguJQ8nWM1e4sz3MdeCW0TKtKFhsXI3G1dEYlBdaqyv6OnGyjVpv1
IzdVEWoX9v0mmvN2nwZ/goCm5i1q8rF1yqfxqbpRKRMM3Q+LOR94neJRX4N7k03g
yn/cmlQos2LCVSbcmgpEDmRO9pZy3S5cePcLbQk8blSqBHr/I2gj8kJdD7uKA5tQ
bbJgt412ZrxN/vePwtxInuLVGZDE/Gdr/zEq+lx3r5m35yOgyCBb9AV6qX93ROBh
yFzCXMb13uqe9Jl5gya+8MNh8UGHhFYBkaQCNZErQb7Uq8WVQvUo0fElB170zaqN
je4Hf6je41m/h9OFGXlp/ZlLCjLnAXje9NxAzk0AbfZac4FbHynDCfhfdj2SfNKf
RnTAPsyi+V/lHeP0a3C5i1kVDYXtqMrnnd+bBF/OOMdwcOFlaUq+e6fKcNuu1IiZ
mqcsUbw8gm3IcqoB/OwQWyZNvR0CcUZ+hZfHJRi9/TQEfBVQC7vsTpNq5Lxf57EA
lGKSjT68ydRbqaOAHxS1seZkUpRCmmhH6tiWpTeFxqONv090f4wU3X/eE+GMHebV
H0m6wvttRxw/r2A9bosPkDqRtWYBJyV9ObJ5JjDJ4dfveFOIda+DzUDQpBa2pmdD
Jtfvtra8ogs67XhxqPvZhWKiuxgj2qMMA/Wa8TnRbBAOEvBEfWwH0s4M+Qqfk/iC
o4zzpKN80A5xGwWPS2LpOMpME+C1c3Ip0hkqrV1Aohyqb2FuDuJjeS7KqYFiHv8C
YNpcAchC/N98LY9PvK/ievx35jKxRqS/Hohrg25sK0uWXhsZ9Q4z+vTgxC6WWAME
sycXv35LmyqNVvxZ+7RFbLTAuJwKB4wY4RERrBanBXvItTTpCFtt5puqh5NKpz4O
cyaTaPht3Lt7boAxUsncLtofOzKL+JS3YiYiP6j/1faDT2OFl9AsRIpwmMLmaAaP
jw9y4zLOpvyLDBMn0r6QKb63DwaveMEh9h5PxXYmAA+Xp/B56jDUf1hvmUqtDJcu
Cx8gRLEqPNBc+gIoOKK+GqJt+m/eAc3C6+ONawy2rqFnDF9gJFdLSLCUjdpWS5KB
+mSfD4Jwy5E5Css7pC+p0fNGVNv7UpODpNuSFEFwVxggezvP5wTvnNjlPSDM3VQr
jmc8bmogS+dCJN2+Wwy9b8NRXWdVh7ADgB+LU1rBylpYgTduCtV/kW3c0uf/l/Mf
0hXK60hDsOY5VvFfi7q+O+MDjqpzDquSlRI7bMCDDwgX9lDJrh/oBc+Y7oWa8MNX
rWB9NzQXQqmeyN2PpEQEFlqR3ssHoNySMis2PUlwCDExxzciDOyGChb5fy8i7MXN
Nf5nFNAC4O+gc5eys7PEYm1pJwCQariUM9VfQ2pvVrUp6bcldn5YDvpoGCWxBEFk
OngRFE2EYsL7euv3AiIl8qztrsfemttnI8WP+mVL27YUkpAd4+ajShUR2bhq+88k
HFdj0ZAkcoVGuuWBAkQJ81TG0ng0FEGxCRhwlsmKhLrV5/ds369+LU4uvXAd42U3
IROTuVmhWrovYJWQksEZdnZPqm+ylb4M76UOUZ5+YZ0jm2KTpMqbecGH9U6ByIpi
sTcNAQdm/MfsQdJCLaJRv4RcD5kEB04wMTdrNcgCye2U6hRr4+ISKsRlVKZaJuD4
TUZaRahH3TXbB5k6gBb3aRwUvjBLufy4oefAh1gB9ce/KkQy2jnn4j70oVQn78ll
SHJCIONePVN711URe4vYJoCphTQE/825CkMQ0Qmm4lHnZhQxPwm5nV0ns4hhEn2+
75Szp1dksvB0yKny+SO5XyjzW9axVcaEvrUCyu9xVDFaLJsLNVg1lwaUnOQ3w2JU
m8vhoTHmUY/odFstXayJuYEWpwprgUfArUY2wgTc9j5PCkNv+NKsmNK5xcUYYAmt
hH1odo+UquLyqJAciejY3O9YWzVCFGjBsJ8hcX3vnrkwl/+JsqzRqWdtfmhcsL7U
6E9LaoTUeL4YiIAskFBoC4/9fs3AUiVEXvPjA3JDMpnm1n568uY4YgpbOgJQIOr1
Ze4KhCgv/7eINgMyiSyr1g55SF9Ll8rCB3ahNZtihl2TBV9bpvNq46CzgQ8Hf3R7
49u87IvjFo35YtAw5G/qFVm0eZD5jooYvGzRD7F/dUZS1CCnQL6mTLj5ellGpclC
GYug64Idokippge3dajQ719T6BwNrthQl5p61NfCx8F/USxs3dQkUacJQrnkET66
1Ruamg9nP/opW3+dRT6FnwzzvQgSCYAyT8HUy++AHL8HbcCL2az0pqEl8E8L+0YM
NezyricjWaOdZ2G1ZH5/SGJd0j9+xyV6iovHntvl/ZFdqSLgBbztLPmgE8+iXkSB
hjo48nShPWLNilYsMbuEp+KZwfH93tdrTcQ4ci7BUFsE61zis8iAGuVYmbmW1weC
qF2U16SGJ1xUQHQRyBJpTLbw1iERDx8YxWxk29GeEa3z72/8Z/1aqWDBGTO6ytL+
yAXzT7E8N4oWLNbQJSicoCb/+vN7xXa5wdqjJvXR5A/cIHHDmelKwpVSvUtrGew+
lxeo8nZYE1yHC9XpbVbQTHwJR0BURjIt8bS1WXErIHYaU7wkYMqmkFlnli2ZUzr9
FI4g++tIpeqlF6yGbUdXWOqNFl/Wg79H9b1A5b8XmXqDEW7as6tAmenSgYMyOq27
mOiQCYbOVMsGyKDHvv9tIYWfPYaf/JHxlYwVrioiAHpUyL3mo9RNThOXTkDEbfys
9+EBl4bEGjYuOG5kAKuJpDRK0L2pwDBgF/akAl+0DStAtqRAcJDbzUAlbHEC9IqW
I2MQX0h+vbXdC8RZk84dFhRezeCS5mhZtw6LY/4EMPsFiebgPonyEkdIbYZ4ZEve
xwizD5SYw+3/ePQDnVPI7uCLsVXMdiPuwxGRZqvYxFonHOUCdw0D2QDwt/i2qNOh
adz3m/lv6mryQAZidNLfQMvVyhH1meiAj/8u4Jj7Ty/xZm83I4oEALRzjfh5ldpi
CUUI40tYMK5svEhSs2Tp+nrJ5itLQqzWibakHt7KCYgFWjy2vPwkT0AZTJvwk70Q
PkjOP03XycvB9Rg+bAdOz+lnWNgSK7WoMgeeFGOHKLNoTuUHwCDY5B0uIZpOOfAS
RoV4efEET6mrusewJLLhS6yU0cpV6vgTSqrayjxObcJPgW/nBUCfIUvM9gnhz1tS
eSZbMTTJWgM8F5/UugX1xKR06DfEoQyGwHnSh8Ouq2kEwSqV/x5i+xgjovi7DxEe
vtIfX4MtXeKf6i/uroVNKnPaGyVUMrDPNkD8BFBa6sGgkDfzxCDqKd75clSKMpOw
/IogdaWwdVY2ksRchCgkAtK8Br7uUbAGxlXcVPas4mW1YjPDOmQEGEhd4n41SymC
7iWl18fHcGKj6qvOlFaoTEyKlsihy1PBTD06/qABC3Es30NC89CkY3M/yaEuoaFS
yAPXk74XMVCSvZasVmiDD53EoLnVB2aEfvb1YmQPU3AHof2eMS70hYBq/3WlS59f
jq3o04JsqRe+5LLn/+iE5BYBpEXhGN2f4L3M0ddj95tYE/6loOqlBMJoSPiO5sXv
drrkAJzTbsTIfghh1MyxZxTMeurnNN//zC0Anv1vx6m/re5TiF+Z2pfIgYetsxY7
Szk0S4dii023J1lYSu43Ve5G8VcJjFz+Fz0ZQfo0WGv7NLTBhAnQzqC1FpGGdO20
NJSpHZqOCyrG+VtlirkpjkSYb2DAD5nrnW2dw8DwKfQ3tHa+LERdw6XiUo0ycSbb
9/ABzxOTGpFnh4G0Im9NiTGj6KrGw3ukDXWYjI1jkac8MmNgfTaRh9mi6AIGgOTW
0INnbe0Q1Cp+WpfPkkQ1hrgHBBHmReKr3ai7RoBNxgxC/YwjJQNWNETVUVR5PCIX
UsqqV7/6Vbf30ZK+nmN2gKAw9LVbFxcXGjZ8/VlU0p1iUDYAgjcwi70ZAU2iRYeT
0yCGSuP/oZtBq1PbYzfLIOezoIbtep3RP8zyE+nblQosNRCWLVm0Ro3vCG5DHscj
cPyK5e1l6/9eg1Rz0T2RFMkKePVbGdDCNTJmSUyI2CjgYdB+/JOs6cbIPZHXpjMu
NOXzGTVV6P41ihjbW07CNnz7OB6QqPQuu5ISGoBVIdsvhh0YTsBEDTmmnIdSvwDj
uAuHOnKBU4ytRgAW5xfNjaPLDZ2gtFcEgEDJ6nCFzjBvuBtcaJAoEbQjHenOaiEk
7Mx8jMSf+2j0xBllHtLysw0WZOZGPn70xP6xDm+9U4NTaPTK/jvfFcwR/CEgO3Lk
6uLJ5FHULY46kQgCx38r11lKBqA/92rtmEE1YAjn+8+jNTVxfpiSsktIEXKJEB4a
/ik5vqj4KQxeiPF6NOXTMc9feYemUSXUnVxvRdHMWUZMpX7i+hyQtbPOwtyIoyky
y7G44sW4U6Z6Ypx2L69p3aT6nrjsUOZVqH3K4QJBYrT79ig7+K9vmMiNZl3lEklO
sZTxecKeMIjEjXbsPoPRN7OrRWEGLC76ewEJoeH08Et0J8pctH9NDgMBr/KC1jor
2rKegIyZPWECP6d3fajUjzYdfSsPYhSzIzp/uyZSAJj+SQHR5LLohA9e29jH8PCA
1BPfdV0AD5RjAPaLkwAwL4hAVGKWaZ1cOur8N3nJ7L2FSpZKfW0hU0V1ylod7JIP
txCwvWXJVtjkgMwvZ5j9iIYRzLQciCDSNX/lR0X287Jp/gGtyCd/mlNCyKWPzk3z
IpweYHex/9fyYgnVpJYxs8G4DTbkC3NBYrzUjUssH+9a0bOl4SEl0SV3LSAgRJBh
skVE1QAZPZ1t2Iiwriy5rRxZs4gG+rDLc6ngUo+44WuNuV6gZEhD374iv3n3iA/n
6DVWI/ti2ubjmpbGjlpMjFeMN48/CLK4T/XDaiSqPdu8eHa8tJ4QljE5BJZWXMgf
1wWKasvzMAuML0Gy4qZSTTCw9iJsHUXMV5F9drB56593Dwdzv/yEqB3gnbUcZDg/
2EiB3HHP/H48QgM7MAh28gLvTlTcCDfrtY1Tz9VBzqjIwmap7AMPywYnrrEVPRfh
KjVs0EFxt1XiGi0hyRDqYUhIDVCoZieFkonDT4NURsMzD/2IuG0xXWbDbaYpCU38
OPTaC8p/DtVZ1lnDuWMdRSqGeJlA4hxTnYGOwf80rTUMcGQNehFhOTLLU7ub6VGK
9vy7PAr/eqAKq6ySaptr9L0afQ926Qzgep9NrzdXC1xxBreSFD+vq+zmH8yNBbIH
zyrKR8Fl/E/MHZbYQrpmJZg5H+gg3Z5vi/gf6FrNYOIA/eVCXvPzcSv1iNfMk0u3
7/R13bfrI5sycvxE/d2Ej0sCZ9kcHA0yLRvDy5dWIt2fS2sxvbiVr1ZyXk6SjRw2
cCZ80fVCvwqPyB72iFBzQdHun/allF7N+68wTSqPLyimoSGl4xelDxFwoACAqY5U
r/XV8EeGDKq1vkFneqKY4lM1CddQHEmtCopT0Q8APHp6GRSnZai/fxRULCeXa+hJ
zX9AZ/6s0KeU1CZyfm/TIghQfV8pl4CwVUeiHWVftFkvewrm1NuvAavnQLB56Bnj
AXlMEt6KyCL+HRcESjlhsdubVq6NBXmk05ZJjyG7kz+Qb+u/fuRQ1hHtIQiLZPnc
zKgxZhnoEXQsk5II/Oshh0rHuDoyEKix2Hg2ZrxlBtvYlxw/51hYicp6ulEo8IHS
lauL4aGFDLUh1XYfWIktjsBLgeqnVLwytB7VN++Q10lO49uR07HxQJ+ZdacWZeKc
JxvuaXt28RpImszGfOl39YzMl3ZuLwcCV6wNxZSpGWn6+TbOpJoqohLXUAg3dTWu
HewoNGHULUtwQS5FV4qPp91Om34rdIX8q3+f0hh8EW0JefP6YQV/SLs0zzQi6zE+
G6OygIZUXFqmJ7W6PVM5HH1WrL5rBbCiJ5RPMfXDUcAsCS8Wx+204nQeMb+beXht
4/IN3ffR6aCriqnP2EEEGZhDKxRernHbvEYdrZQDTFUBXcqnt42EK7riyRosUcyc
x8vaa9Tv+gQ9kOD0/sClGH3iJ0KLDKf3kBB7k64k/sL2siJNt5Y3sRr2jwMi8qqP
s5tREvlgRs0y8HLonPbiSDf04V2IEn4CQcBpGgfHMBKoRrwzQr1jm4hiPbIocu9E
xi87vXp607RV+NFf8eQylqgWN3uuUH5sjjOi4gXpt+MGaTIPydi9SaknPf/1fr1Z
UePUQoTAfyuwFClnXEVvZh9YRHMsIbxuqDDL0cEvlLJTinsqZIdTwg+N+O+oCtkR
I3xrP5mCtXHviQlx35MMp1B3PmXE7uLitNdjTfvH+0/+nDoVqFS0YtNtjWQjjIvj
BEPNmV4B2Qjbm9R6ThaT2C571MBvzRFY65BAxEFtNGHHGb1s4lkI/p8JGHCMjHVe
chqb9vStXi++uuY0EQTklbtRn+za6R/g2iOCZfxDbTtNhdQ4BZNeUxqF6gqcM/Og
4SRu0TipvJacGdSUGGe2ipZCagNp3PKSI6+JSZe69NuCKcmT4wJZbLD0jSPZQCEq
T2gpggQzMbowz/ZNyqu+mKw2ABx0eDQ0bBpgtjEQg+OynlbnnGMW0oeKJyhW/Mjv
Z3tk+r/sfNgNDB1/XRHsn8NOseeT+7ZhmweTx5uQqzNG8L9NzzURYaGFwSOJlfdT
qL0NFTNlUPGdYOPWSCoveBPtZqfzapAWR6XZV7XznAQCw8mUwEHFFiyKw0alb8Dj
60zHRJQCYHruvAyL7XicbVXYiN4Kvx9zzcbxF9jJJIQUKiy42g4K4zQ5lFP/eTN6
PHam7D0xgwr+0rGtMSj2bFwDGtHneQIIeb8UmhOzBwhtBsu/V/0qd5Mult5e/xOx
u8VFmVVhJ9XW/nW+1t3eExpO7evilbEiOEY0APXd5Q82NQOA3tye8LZGrNmUrpsY
wKiV74OcmQhqBXZC7tADMVywMhYGdVpLCPl4Y6VU5s+85Rmt/XJJXfeY+bjmrZP5
wE8t6AetLEydUN7KXcO/JzOhJo76umAAIL9lAGZjjzxpnrA763mUd6dh0ZjF5evb
PztJEjBquuocbGHXudjFqLs1toXsgYwTaTbuQNFipBaoursxtuHrKyuHSilMhrQ+
j85rGs8pZFffMn6JQdiX+6rejSf5lRh+XYA4vRQjWyhaC4O8BRZOyn9ohcyiGSO4
Yz2bsuKxEVtspEipKA2AibrLLEzb4s3vGSTkVZGNNJH0nejQEbFxhQwMm/lfSD0I
fwq/+XXhwhjxyraqTRrxtgL2cz+9OFd0eCq3XEM1+rxB1cbAi2HhdCi/oJ6L22J/
wGTf2lqfUY4HQI9BGDT20Tno+nz/NkTS6B7PgpZJxypX9jCAZoM/CEPtf+Q/H3oc
YNGtpSiYgapVz6yVaJBiBzNww0gz9WSQohMWSqzTGo2rcgGj2X8LrOWUALuyUqQA
fK1R22IerAnJivIKrJo8rGijpfwxj3QWncaeg5lqCWwWerXgywjZOklq1KNQYiaN
vA2I179coJzZc27A1XQ/nG2rDMU0/R+8NrC1l0JuOgypglZdoceTTo/gnxjLHy/P
X8Oanttp821QKfn+24MPVqVkkWMN303PUuvWn2gXrM9TPo8XQdPuNXYhDr6BT3Tr
qMYXhRWem0Jim47LVznDpI2y+oGikSRKBx3DL8KEvUAA2EqxpsCmFloXB03bBNab
KrxUWnMhIDSPSt99l2nKtU/CKtBzer9XJ7K42TZipHSugtXf5BRgAGGNpR8Q8gy5
047H0I+E6Ng5uHXq/9XvFRByvBfSb8ZHXUzZ0UFbrzxRhhkc+YI2g7R2GOe/uPiE
umBhSy/R0YHBpBgxj9fDdMubO03kGihoB4AzG05uH1K6H3CHhjMRiV/IKVCMm6Lb
Q8JaQshULJy/FAAarlSlWOgR9HA7Reolu+hl95YeL2w2F9J8Ng+I1BczMZLEMdA6
rTbFAJ7m9VMwnSjjwA8X/FuDyhhatQgS62bBmnWBZLQj8SsszGRKny2xn6j8/zUI
3SPK5B9A+M1DD2bprPiou/yIo4CHfcpdMu33K28wsL4jG9eDkfc3TUNq0IJUmSSr
TH8ah+xf/THm98IqmO6e8gQoxc6AWzVsq4MLXLO2HOiDsf1a1n25KLv9KRrIdqNW
WnZfNeK9/vi+QxIn8zE7J2wQ9RoRfGHETuMDkgH0QM6S0QYRMNsU1G7ipE2mi8+3
qfRJUdpr/31LPRt11Z8dobZAvJWjcBqaWX2ibchtK6cO9WAlprMjqJfloNoH0B44
r+OwKq9e/qR9ockWBTdWH8+SuuWVuFQsRAR9z5GBWp1jfDG85NalsqcksIUS6ZV1
OqmyGi3Cw+CgIOC8zVKr6Qzvi8JYky1Kva+7Oef/+SGdIckAp+wP8jO2L9M/SNW7
/3FShxai+MtdjfTcwXuF7D3ai+CwDmqJimYec/lWaE/q5hG9NC1bCuya7A4uXgPn
8xDqnRUBhB/UFUATyuoBoDmuGUXBTzxVg9I++4XbxTW+51X2lrST9RrbXz+wVjFB
Q/hz5K1dy1f6LPMnjUT02TvIbi+94SMcRHgcwRJLFQcyUt2RZdrhInHf29jSGAHw
pxrdbL121GrEd2QvuEdVtYpcsnMH8+eKDhnRduJ8cccSmFV6XEKk8q4VLyRrsknZ
rTioKlJKyFCyQvCyKyPDR8CSXW9KDNRCGn0oTuiMXebcl2R9mPPdp/Lx/b9zRCQQ
eN/OyhE56Vuuzug/aw4UzCauxCpTqfVwzRlf4cDDRpu5OWux8mYnMVdh362s+JjU
1AuSwpB5sxMQKkBpiqZ2N+oStNSb1na+WNrAvnSKSmJ076UcRKey2AJpURGwLh2/
zer2benSbWZWDkb2+uTEgpr9yKBZSWfpyaddgujHw8Pqlb5O8xUINPLN04ditNZK
P7Z8RXrmdRyeWwMrp0Tl642xIawWZANuaVKtvfHdQBhtPHgrWip8xN83grheDuZH
qeS+lv9ZbT7Gz1UJpCt1npVUlUQdHmeYA/bKr4rN0fyhQUfa/l+iazjPdOHJNxcN
a2HYYSl8xyJnRcuxWCgF+FPG+8+jTP8z4ukItS0jxLcgLVVXjW8aI8EBVBl2hN9z
jZTPCwAXcTiTKNRZJTUwGld0rDpTZYyZLW+1e0eXf1WIXNT2j0QRdPprrRc79/bw
g7etUGBD8Z80k1pAbIWDxFX+QYf1AVxvFb0CoQ7ZjWlcnHMfqx2lrCDWoLaDgVVV
sQPk9PzdEBKghJJB4yelDTWswEpqMoutolpnU4sQWeFXH7Yw/JETecSKr0bJdhDc
calXdj+qqzuehXQkEPEBuE65Lszmx0kx+7Rb8nTI8RsPIkVdIo8Zq+kKdkcZMguG
vqdWRp/x1+jxcRl/ro75qvgzDYMd54mMMSd8WtMbWSd2rjQaOeENLdhULvV9Wqpj
9rAltvXODgYjYq8fwQQGtR+5wjFA1S1WG2raKCyETQKfMM+yzT/zihmNdnkoMBCf
4/Yqpm+xNFMS+CPxCnOeHZ7V+6QmFGtYTz0XnNRsnnblfM9ZBMQW/qsZOAWbUnK9
YDHi0v2TEyj0XIDvV9dOtX0nVkmNAEzh1i5WHY5fNVMmhr1YtMSsReSSHYia/XGg
r1mGsKbfez6G8bHOTH9BPAYRrNX/mHFfHrYeKaEPLzN42wpz/99tmaQxLBghM2Wb
YUIsziwgF+2o9t4iGhrJz9lONUilrDOOmD7Xon5FCJDn7Q5StQbQ4xKIxvZup3D0
Z7TaEZNf+CnUsI9Z4dvmMipReE8tHjH3M+oSSi5t36qDoiApgHu5MZPviR6y3KCQ
HsS5cjJHe2vZvZpzGpdYUfxWGWG0Z5g4ZurW0Ij7SUGjXqda//80iWRPNSawdiuf
lH8bSeaPzLI2jRaVLmqE+1TxJ7neaLjrsJf+UWobq89rtf7RhafYgV5yG10s0/sw
QP0hqBgLFR2lbF95hL5woO1KzVRWOzG9Tnv+dVcqKljqU4/jmn+mwp5dktjG+Wnt
8wYjFPs5wgf9DQDeV9a8wiMAMh4AFs+o8/hk2wl402ybk0K3QKBlUv2RY8SFhxnQ
jUaLUqNcbjXKtpNj1p3NwVTaVFIQarKY4xY9q6TcbruKTiIgl3izyD/j0JxbQVwn
iSA5kod8AthQiJKw01u1wZtPGaTXXoGbr0Gnhteh+PelhnIqgA0edXdgtlgH26jU
1DX9DLpdsEMC6jsldI2OSXzemrJIdKazcvL1thAIZds+SMyUenGmipL+12FsbCtH
KqoVWzgbyfvKRD1zdascSnP7RS3oDlzR0Y3xEGJ35AB6+RoPJW7HIdeSkRamuqZt
0sIb9nklsFcZ/8r8Pv/UvaGTngERYwqgXEhP7vrk40oQXEFZNbTiBo86EpyyuNNK
ctN/Tuxq+T3vwWlVMqOvy/aQK/PD8CucXmbCm4k+hLTLiwdHWk0ay6TPHk8SOWQC
LEkSv9x0mg02aV+asGjaEvVT3RLebMuSObCgKCnz7X48cEZo/+qih34GMAvGDA7v
DrO+huWPEgJQXXzB8pqMKEYFmcTDVv5PgM5YwTWpZ5xcFH7RBJG5Tx/Wf4SUzqaR
n9wHAngX8NSKnapuYquF26C3M6LyUs6OVggdMGmlt4B+Q1DsbyNJBjATPwW6B+PA
UTPj3dhRLVPzv7duYGi00/GHkZ7zmx14eOoRfpL6j58hQ8nQoiHtaZ611LdxvNPG
JQTTodjzpsDwAgJPAG9KVF61Hwd5jWCvEp5HUg2SnfOkl1jU+551o/rSUoXgjR1B
/tpeVPUqxoEBdhVF3cvgocjy9x0vGWvZPyIUmh5eXRIcWslfurtpDKMYi7oQCgrO
u47x3lzzx5Moz1Kf0wVlEoTirmn/D4sIwgJhhAm0KNxE21NY7opdBPpRH3SSfnvD
BLTldGoYNIP+BILLR5DiWa8B4yDadZ5mN9NyMu8/fPV02T8ngW1Z7Awyup5Usf4S
KezMqUlzLn8ErsKk2ARzQDGK3DFU6pq33WzhNVT/gFElS4TTo7q9YmdbgY9piHA8
Z6fIyfPjGmTDxkq1uu6mIlkkp0XTdMuGX0jd34XHsIiPLZlFDxs6i7TjLMDXj8Z9
OkyIS7H9s01Qc8fclOcWyPpjhhPA9VvV7Rur2jRL7kaqw8ldtX3VDNBVgYovW8X9
zMMTsRyt8d9gDwl/3AopFnt2Sg+/yzK2962yHjbHQNMoZ1/8J9lHIJcYwF1aJrww
X+B0EyiohFuNDSbM4DfMS958h/drIXbXVrGStza9bdn5pZ+b2R2mcUewb0/UZJB4
7EhFuSZ9gXljsDM13VUs++xpZJs6lqB1PpVZdSRyD5x3UvLPa7l71Zp0MsjL7r04
GLMXquWkBExJBo1xyMMUug3BCHzuvmmCWV6XX7CEyf68jDeKnRtH8fn4HfmyJa5w
SYnCpWkHvHIhn7xmIUrs/OAYslnOUAC7f61ZiM3Z2+c+M7Bu5PU/e97SzZUf6oeL
DpPrmCopiP7Zxwaiulps6aPH7hyLrDxL/5dWDMt5DQlx0dKktHrbIj2ezp/EJZwJ
7mPFMBUzH1UzN2k1vHe4qcb6H2inEPlyYlQ7K05wwsg1rm5kwk5nMyvNtvCR12DP
/SObOfi4OTuhvnk7bM0EtA2JAnH/Y5jqNi2EjcsFVTW64MRoCLloRFLa9sEFk9Q2
lWa8FvkMuDvOXaFt+nZKPXxzFXVXzyACtwPXqApjiqg6gyR8skCTqXm2nfwqFBqj
usN4FSG+vm6nnP2+A8rpUH0StL9IlHzLTDuX116aHeOObhzjKtw1BC6SToiiVUIY
4kMJt/DZkC928i7hIecewMV4ZVA29uxJMGgLs2akH/vitEpc7NmeQ1zTWKygF69w
3TMYKJlZccH6nPk27phxc1IfbSu2xYgA51AjPE5ISsDedOankDUgxOeWiQpo1cUy
jxO8Dss87g6eHwIS68hyiO6S6XopnA3+HErshNE7FLKon+tEO5KteXlj8CRr1Jmw
qfvFCrzOfAEJ1LR1ULxXLMRc/gWXmpA/bQuV0uBMlsEazOqBRYCvYp5QDgy5ZEqP
Nl7rDvLTRVsz1kT73RanrWbDBn7ItSFxsaqmIxyd6js/EjmVuJhAvorBHnTogg2e
iI7vOPh6geWNZh/x7nhUHfehCf4aWD8Wx70uY0lBMVU2zMjiWxbBUxq1C678eTAR
8Rb4QbgcEgMpogSONfKiHW/hIlDXFlzFPFvJEDTH/72mTXRq12O1O/8xlgHpAPgW
4dLpd4CklAItXNDau9H9AD2ZHvOcQSI1DueuZDwCJB3aHUcl+ZaC0duU2i7oWcdH
SbbHfaYMb24AXBpeNa8ot6XAM7BwV6tcEi+iMpwKCNdZCwgpMuOk6X+e7F1+2ecK
5CAuQAScvsGj9AnGTTmquIe9Tf/FT8xZs6liQptluqXJUJxt1yAqPq55NDWbHNFF
6Fi3f2yKsrhxbbqBYrxsxrtIwzy8/4v/0XVRkMl5+Pw5eYyy8gGJdABD4tSpceCC
pQbZ9ZWPs6rfw7YbalY4aE4C7z8KaxwAO6/VUmXpnwXi0xEyGFCoUM23ejIlfcrf
oXjMrz0D5ebgM9MB3uATMD1RuwxwEgKoqdcYssJjJUZ5uSKDbkQr/4v+ALxGvEI5
Rzk/GuuyLK3OWnEIKVEVr6ikmzLes/ckrfnZ+LKMK/QRLQdzBAiVaB2vXE0KaIg2
yoHYfYcROUnZ5Fnc3Ie72aW6x7hM0EIW5YAYZIhA1HXqGp5hpJEMD7yXvU1f02ZS
iYoVT1MRImdMRqem6J/E7szhE0X/SBE6Z1yCKGDYK3Zgw6aShMvLiTlF8sUIjJBI
xx/bQIYI76Fibak/ny3Ui1xa/jPlWVqFF990F4AOlTim8Gq2HFBrs7yPcqu5aKMP
Vk/1+SR9qRv8okm8O9eS5ZRyGR0Xw1jgMTfIiGqqp+zC8v+rWeConQyPmLgl8BYv
8rtSYIrnsO0QZV5yEV8MUCj8C4O6zQ4V2bkrCQPSKQ+j62KaAWOQNL1zD4lSRnme
evC6wx1Ow08WAnqPlUWr4uN15zLp2gI/oBhgzvfIBvtKsvndnCs6IZ6+uJruPQYk
sjIsuvXxw3V4uQV5Doc6g6XAmtV0QQaWTYnqjMvw5ctJy7wz6s019scfWQuR/uhU
YFYJC1Y9y/ydDIXke+iRXgoopaHYXs+AqFk+nD8D0gvWwAdy+czdQen8/SrmAczs
ycqEFh/a5O6jNGA9uTG0ZmTbkhPRe8tfdtD8H1DtujXAUmoRRWqqjyp6JZ8igNqt
k/Y3srxS50oeT0/fRSBVGOAwWlxRLf1ZY89BoRHLkFr3x9RGnbo1sFXg9XBt4nwT
N+Aut7RhqqNfz22MhsO12E4UwlJOBnj06jvRDT0fozCdwZqupL6LTctipOnBMEK2
mLObrOECmZxq21M7MaPClX4J2xzaNJmC5qVwdKNTbW4=
`pragma protect end_protected
