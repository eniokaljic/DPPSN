// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:45:30 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QppqojNO5ZPV8i0ukd+kTh5wdneckY5f5wyhnXWWnWWM1eIFwuOoCiUNsrOuUFSb
wMo3Kmg4aL/aFfDQW/Fb6qn/rTcTWnbb+ivmg9lUqDDcYk+6KAtwBD4s+pIyy+Zc
yZQ7q7z0uD07R0aphHiL/LBFNt9fIxQfnb31OwdGH+o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34720)
cG+cN1tVyY9Fa/j74+IH5T/j0zI0LUMNxGiT4udc5b8L5ismtebv1onw5VtQdx4h
8pydcMGOjpVJSQD6wa7EUl55bzWS/856DZTg0Kdm0G+/JtVcxQxKaBWswIsoI4VN
t3MCJKgki8QqByPNq80aA7qsycxuEg7orhnYz1eqqb1Vh618ClHXnO3QNwyrtqEC
cjwitTizW90e0UcAO/RIC3zjhd6wmupZJ5Pj9lDAOycYRMtIAy55q+Ypu/JadFro
ofihbUcdIKVwXAc85peewFIavYtK9nCMLp/YQqgnBdha1oquh7cLsOt2oYUUBD24
lIqgBh4xfz2UeSLlgnl9Po1RwDEcURQ1Xn7W2pVU8euBvCmtqOm/Q4DfevIu9mlW
KduzCCuZR99+XukZLJgJOJVF0gVerUiTihimF08FTsDk3PnjRlvmjmfgmBu+p/mc
KyCPpPLJCcR7+AQMhmdcpKUKh1dkNN+rrbLXeUwte3ZkiOXRZw4mrJaGsW4UNDpu
7/QLQLITIG36kFMxb3JYisofpNZXmCdfo7RnMlL0yF0eFhAl1x9PrFVAG1tao/TC
S2wRBoMjLcFdDBB7oJJ9lI2SZahtUcjbL/Am+Vj0VkHeGupSdHMf7Nfil8bAKGMQ
WHNqAEleue5U1zlZxfgO/Lk14ubwIpJR5S+OCYhOULvdyVXA/T5NtpSxfCtV+1aU
fe/BcP2U3wE3KPJRSDpt6H298ta2qY7BAaBrKXCYNBzwxdW3uqYtkXPiClVL4E5a
nf02pDpIHVNA5keodjNXuVadJBRSBGQSVPXiZq+X9p5toBlxcHGlFTyMMfZJ7lIR
YSct83FUmzyvQbLqtyJFfctoYRDvRJ/lWq00P8n8NPJ5B8RYIMYXNt73D6f4Fz8f
dfJ/1ddbHZ+qeuNtxT7TNp10R6W6c4/z6RSdpvTSrebpZ2hhUCzVaaMeLwtgogqv
TofEF84DQnb9B8PXe0iXuidRp8fvorQ7kp718SD+zrLFB6n4hM3sxP3V9306s/0Q
uXEvJlXTdYpc/5KqMmIPSUOk8+GosodN+47DFkEbhxUCvmppUlLxJI6dSz1mnrUb
39iHbFkX1U34tRUwkrbilAzCWCb4sxScB2XnNHdm0P4u/JeT897WkVDVmhySS12o
bcDe73ju1VmFhuqLRnxU5F6+NnlkgtkulWrRbeZ0GFNrP9DYifJx3DbmCTrrZUnV
bT7Ukk/EVY1ems5NSdws4b/Rfca+nZJ124UjIR7pRbR5h21D2ezYa8IEVHROV+Gl
O0tmx2vr0V28cTRr2wqhK7ysim18V8eZa32PM3Lf33287NBaB3my1U5KOt/Nbw6X
rp9AVUn45FR1tZ0tl6YzfWJdzt9Cq3wTXt/R+oceK447Vlnriv6m14iguj/ZfsgY
KM6Gs+fUJHBpUecfRGDPsf+O0FGcFY3bWKwzDRs11Rme64oXEjrfJCFblEldiWEI
AYEw7+/h3jIWkesyA77nL/6MoGYAnp9+YPuWfzK3Ue8EIsiWtmTonClzX6X5OEyT
7KRoZQnwNBoreOZvlLBlgOITnbjxIm1jYCsH348jhE10sTbm0QtjfzLlQ/esB5fs
OgP3KhFAca3eQJxUK5nDpLIRgOGLjaq/tjuIj3e+g+OkNvZuG09We1FKoj3wSCoW
b4TV9NFMEPw1ENoeOyeOgz1/3AT1eyf2+4EaTiVv8WZq6ctgcSZGwx0U/a37hVvJ
pIFQQrEdbm74kslCMdH5lTqeFDH5G65VY7Q7zInnXeSxMtwYrtWLgfE1tJf2/a1B
Ncn3uwpnBymHRudp5yIVfOsFwxfsrmmDxFH5nsWQUq9lO1Ld1Orrg98upvlDR9pH
MZx+wk/f+egua0bsgIykl5uf3F2iWr68/Kq5YDr0O+0RKD8IOe4CjyDiA4fNZQEf
A/RgjnIbO01wFm3Kt6RFRZ/QnJh2X8lG6aJ3ZYNDa6l5nN9EmtcCDxQETgzdH4y8
iIFMW3dSH8BaCKiPl6ljv015tFkSFjSLnSOnhLw+oENqmxNwHvOEbFOS6OPZP9so
/ooVX5yBQ2uvhnQl7i6SiPCpA/wPfK/M90JYqZemSPvnX1tIlJ2Q51304KSJbPu6
dQ5Pyg2xk4yr1Z65mLL3q8hNSCcLGPf2/z8USUxlfkKgOLpi9NHM+WODur7wd0xv
0b1TtJarL6dILR3gUFHMfqkGlPVGM+Aaz5/7dabdPeKcLZZuVnMZrzThHEhJ+N7u
d9IMcccS5hd5PewqfjphgNUPgAULiyGlX2bedORT8Ymj68IPPrsHnk3gO6aBiV1a
semLwPBF/tvhvOe+U8po66eLXy1Ar19cpWF2nbdDmjcbZwNO7Pj63yVe2tNZrny+
Yy2TTgWyofbGr61RojSm/byUMauZGYgeQLntpRQXxW5ovZtKXJvC9r32fPbXoFgK
E06U+xAJcBpO0Oh0pSPvW8nXeRqwNCGpH7/FT4hcsYmKyOljOGyRHF7PnWKxsdQq
SDAApjNi6DvBLCqaiDG/uVmLsjtGru2kzFm6ELV+r1udgyL2CpgNsElME4ey622E
QNES0eAHo49LMM7WEXZlj5gTaL8EENzkXyOUtf45zbbUpQi9870KyyV9E1lg3suw
l9liAlREIFaJ/uoI90Mnc7NOkTqLdV0mfyZhMAc/GRnxnjndRBVfP2qCeEirObRN
DVjMElF704HbStn+XY4nGfeBZlL1Qi391Yl198FcpfbjrgkSOpn3H5wC+cgu+ce9
UvHvqN/BaIyapXNX4lqkxhqTsGmRvEjEPl4/cM35ntEyxVVZzdeVN1fsuQc/vqN7
MpoBGoryz/salQrRk4sOAkZjTf8eR+eClMY1ar2zz0jz0wMK+VcKMoDAhnaXMhCM
3IbWYG5xjHp4kPFu0MPqTXylcBa0Vrh9KrxNG21MOsU1cN+6l8ZlcF3mKf0YXitA
xut5/98+YU93ujOqBx8fBWzUHAsObaXr/FWFxbyrnVuJcUW6wmowP3qu1guu2X1x
vKfk/KswGA/OfFqGFFjROQY7Vf4J3BLBmeHvkxuUwOrny5Va1XbYrYIJy53V+pWt
dc/IWMkCiarx9y44IliEgiJv5BjNeX4qNO99o8dOA3Q863mq/UnI59O3rlXm5VYo
3rfPYRLCml9fB66/gKlq/rzY11c6It33vtQuzpej5Mx7Ez5yTTi8zU6n3kfm0yXS
faShRhEtwSwc+QHfEtMeQ3xQ7T9JhZXE/qQOArkC0Hn6Z4LSRifvja0Gt78+Xgvi
22ig8XmnYivYpmtZFugtTk02OBzIGPuJzZJaboK61M9m4VD39h9RZPc7xjYywB8+
C8cCZQjFcGMf9N/g18OGzfN8RV5LEUfh54gq8qwpnbHJcsBDCjzMErJkJTGEOEYC
Dvq8nYuQ75oEw4bORH7Kim7rZ9wRu1qsg6ql0IJx5wnvcgxSFOKIrqKy1T26YcGW
bFCypg0yayx/uiM5OropIXAzEbrDYccA11HLh4nqoODa+dQjvroAFl3um/MlVgR0
QSdFwAafGB6G3+gVOgC3ET4D5M+OGrua/EsSu+WqcxlaqTcgj4JmdBbGnkVmxdDD
9wm0Hqk/YzIc7Yg8g2x4y0H6rrSRW4Rdi5mKtXpUS8ahi/rykNjC2l3RrkKrRSSq
k7u46lEGIcDEC7ajy8xg7E9feqPoAkWNzEeZaTqWXkTq6cCcHfApoILgQuJMUip3
Lx34x93dpaOgQ7Kv700iZ5UV57hQiMNgtiiLwQvCZfrGBrPC7nl4PoSzFa74bp9c
2EyazGG2/echNVaMrSS/zwG2nFzGEn9GGAR3S3MRQAIeskEYprcMHXyPEo3HRi/+
HQ6vzEBbbky+Lo/BQTumpHxTQDESBqNRNe5dKgkjeDItC76lKrtQTg2vOr60lm9w
+5tf27wPFpnr8JMYDkIldpMCfDjl6lHKcm2GEkCR0up1sbRkA+Ko51lU2xd/NV/A
8NK5iLe9kS84RJmGkUVHBzi3f3D2yRz5sTc6xm0VEtmScWJh5yCvVbwi305xKb8+
uf47sv0/5POjq0RdsakJzCL4wxqfwlDj4v460W93h9AaK45VetO1QL7gLSl3Bm/f
K6/ASvzFpYNLX2RrZqAMx9LFo+a/o+usHCXM7yY+wwJEYWayyxl3oLBEHp6FGTJZ
AfzC/ZmVMSn6EHHVxNSQ4rZS/VmlwdNrRyDRXQ4dMsAqnNgKWSZgFnAS7h21VlzM
0oQdkeqaEzjYm1/7JKSjKrwlHwIv1gXiVGMaB0REfKwgi+BnwdyUyXenw+gFsbL7
rAVj1CLMJZnQsudbN0IrNSWoyety7ReujjXn0d0IwzgKNRcw/Bextf+T8do+TlfR
wWZXwRkZakv2D/fhG9xg/A66R1q74uPEbp1xY57pWvENThdf7Oi8r2+XkiM6hssR
/wfTx3uRzBkSokwuJ7SpQT46sEKFKgoWoU8yHGtX+AcMZAQBDM7LSX7DWtyBZhz1
GVXNHCbN0+viZTrCuZzjt1BIVO43wkUhcWJLE3vQvMCiIBfS9mcJXnNJiAFKB8Sk
TKsMskThMXIBD7qqReQ3mCFR4yK5/07vQstK9Minatj9zzSrJ1WrSPW6t+8QeVy4
I1SewXPniyEgWfJQdToj3iYBXlHCNtRymWdVTN5aJwxmDYrUyJv7opKom1CgE8Rd
sfI76UHpD56pqqrwzRLMy97qHJmw8x7chs7Cc6TA3PknoGHrzfEKAf9qiapJC1t9
MV+pzZlU9FmRhnROayYNKmvukZ+lRGMkKaHF3BZ9SF5qaSalF82sRuPJTAgvh3FL
gpnK0UGwil2fYOiR0AZ486sbHiRBa1ymBQY6/ZRg9R0UtvqzTEXChI4NWQf+SY2m
Be9L66OOzil6MmDZv8FzpkJtZ5/Z1Z0eb+7f5ZThnXuqERcI6sAyLtlU2OCZvOhy
ajypecwUvtic+B4lsWBL8mi1YNSGd5JDJG0t5iGV8FeAWrjkQen5MQSBK7QEc8q7
hv4pxRBL7wsYCHk5+Iebj1HnWf0yhRqsmeqDarWinwbx1RnNkBBht2KBkKbGWxcF
iJL5cOd68sXq43L1ipHxN89/TnKpJdy/XDF4GU6ZzlHBAKyO0WcBfdo89A53OLQl
YSHhv8gPMBPWp+KzWbGj0HmwU19tiiAovJgV3CMVFcpTDqaUtJqNpyH+VBMReCh5
nr3MbQ/b74HPP0jI4lBLJa7uiGqiazek1yxviUxhDmaubn7NMmKvd85KtA7vviy3
BDvTQ5stbd6Kz/xUSr+EU8kjXoxbvwaPsrSQytCRhuQj5pj1+jpfgiKEy/KCF8/l
xSBAiwnGtZIf6asxW1I/wLTFuY3QmMC3gO2ICbGECj/1RcCznrxhPIlBMEAVZ7HA
F6QOG2T3yAyHcwzBAHxpZUDa+g9/GyQXYr97zJLIR2YAng8vUqa4DTej5pKjG6pT
myJ6OQqwpFRgZMHDZmb8XkSCZ9qvT9wCXdjTD102/cvEE+APk+xS23/19bmV51ra
ovkX1Y6c18xVicxj9RG/Op17dmze8lTA0QcTz5pF7cAo+iIN4wTLRaoSSCgh+z4L
1Iu0SRSMZ0sNXv61hotz9F6CWYl0Dn9C42wlVUUGrLQLuTzdVBDhlnrcs7V0uRf0
hsHWB32utEIseKVSTDU2+9He5mnHIgMPr/RKjGKyX/7begFTWjmNBudZlAiujA0o
B+938Ewe5RalBY/lFbDxuDx46CCoMqQsEw4WKF9JlpKPqT3q/Jf1lVC+Spqkx/9e
DX7XjAmz4i+KpUcCceLMhRCDpf44K9G0qVGLpOUKNcySfSTDcmTuB+MifszL0niI
ZXBClGZxW6CH8MQr584PaD3GxtegHpdvs5g9zntRz/Xak1WxDsAhXaoFhijpezzI
Hr//Ly11VGPREqm7bKJIjKqwGiLo9INTJWpZZwyTLEp9XfZVf9JdIdisec6OKtoR
5/SRlXLfuKRluxOomg2lTIkAdQZ2i2lnM0UQkU1xe+B5ycfnBH50OqU6Av5drLVs
1koqjnVmTLpMlgm3QlndR3GRlH0LlkrtIbFpmyeEyfCs7opMQ8JtqwqdCYjep7YI
33Nro4RA7vvE4DbuOGIq9CNPwykBgNYdf0WEnlAKrksgrJ0fqhSf6yVa4rMDPIrH
q8tupcUi9dbWqXpwQ66FggjMvVBB1jRGbJI38WSZTvIvgfOpe8HyRqY6wkBlAL3S
qFItb2HuBvVL6OXFCDny5Dj83LWcoQXSqElqwbukDY+JF+6rsFyHuwWZMhd0HU/6
K+SBMq1dfb3fwA8DthxNBzvP/ZmbJT6ohOOVt91YiBPjvwvI+12rkVE+n/EE9cQN
Wq2o3m9v8B4fjY5eF0r+wg9yoTPSrPoQp6ir3pj+sdC0MjNjAT2Ok2vJ4swZjv4q
swh1DdW0MRHWDEXMM/NeHAapHIDo0XIxvrFrfqhct3WnTwgt2BJH6XCyhEl4MheH
zT3njrmA/R98Vd2CfecS6npippnUQ5HP4veb/AiVmIQTn0ZjKPYpvmuxGILLLcjF
1Mgaq2O7FC1WaxKZVbFGRJ/Ju4o7q8LMfX2hCcL/QvyJDgxIscu9eDVEmFbAuac2
7leXDzEg5LsAOzBuu60KezxSIvLj3k56wKPhyLLubhZrJtkCqc6/O4eK9HekZ17h
0y8b1HP1nxhnQtJ7eZyhicrxZoRhsW1Rp2n+KNMjF0Ozzz1Zh18QHGRWIQcHBBJl
m18QKkd3wj6UrUZtTjl6Ij6IBA0Eqwa5/7q7sKn79gcPthMyrGB5oJLtpG3SPGiH
o1ZS4ANde4TLvzpav1wTXaGQcI5gIWLZuPK7Ep28JTOutEBRqK16uYZu10aIGmiW
eDA2nSv1ivJLXcaqJhDMiOBos1YfrcJi/3Dh2QW/tDF0QzKw2XNY1+IFwNXUTK2u
Y2we74Hn0B1YNL2yriwIf2nX7yKip7AWDQKH3XmCJNUhKo4Xw0C6B9gnKvPe5TlR
l7Yy+9mx1dBekxEYY2RWHCo98GpqQNQ98Nz4OQpvQgwCIIcjeVLqB7N6aeTeGZPO
EUt6U9dCQNQOlUo/mJgpvJg2AKlg/IDvhPfc/likMMRejeD0HV5dsf2Cz+WtKfBc
dx2wC6ZRvj0q4I0nnGQx/H/u61RlSa4paIZ39xOCxWzwKCfSq5B9KyX5sLXCMCn4
rpWfqVvj6A7sqm6rPvBp42FuE925vQtud+x4L045kqBSA6bU43ur/yY1qyKVXNKn
dQxHoG33OMBHldhZjINCfsRREDHRwKNysFuMcXnPjEYPTRK7+92ijT6IBToz9mLB
fOF1wjQVxUoSg4XNb91DLoUIrjbNWIQSUkAuAmyazRh49AhyFmqH+6rKQYTMlfaz
5ErmGgBPETc13bZKTtd5f4HAjW47Q+01TU/JvC5ITV6v4ye3u6iQvabxp7vjrT+T
j3pfota6jqF+aoZiqqXx31fpmA1Gx+YtbyZmSX6/Q5cQUpyt60xEF0lIwAzq+iUX
ruMp++kbvv7B8tsJJaCpqxTmJhEARrFVxFkNq8PJg7Gfbeszb5bQ+hHQEOk4rKpL
M0QmHZOq1U0KvsjuZUHIm7gLFmVC2D6oLCTJ+5UPP199qcJJItcZPAMyHHrch+q2
/kjwVR8o0ZK4HpdtP08YmKSj950ucvODNAB2Jfhy/HYbDQern0Cc85biinvHHsM3
nkH+Mm9w209dPoHZpfhSbtFZgdzzm2p9UFlFsT7nCFXveIOj2XabMODJYaWV4U4c
sobj/E/6a/f+b7OZyj57W3MhEw3Wzt+doph4wRRYZG3spGintIpMovQzdit+mYRp
e5ypYkdZT15ftKAsrttZP0J6A9plfTeTzixLuwl1zAL1MvEXRT7UgHSKFGYx9iZJ
lVKCAEv+KOdPRmMJzGaB/a/AjR1PCeo2qwlaG4eg0JHS8/l3wPXeG2fYqfTuqUPU
Xsp0MH+vfBsVIDT360NAfR9oZgcX8K/3iID1LE/Ltc+pM0SVrMCWa+iQwEmpmgmO
oIERUiCjrTK5vJv7AutlfBe7uoTdbu6XVRsyQbAPVfVbyQ1zqavgAP7SdwwyVsZv
elJejopz3PYLcWRPL6qv/xURBRecWvNFpPzGUKIfIDRAAzi5LRydGXUIyf1QxKFX
gor7Vr1gJJ5vcP1xDFXmy3Y37W8BNIYFt95kWuRICt/mYt355AewNG4LlM1yAYWo
q5Kesq2SgS/GWu8hFdZ5g3n53I3ASsq0qKr/1/8oC18L3kwiOia9NFlb8TpdRLhk
ToKwOATxI2yMZg3sNwDSTJ0gS+T3fGOEbbdxwix5D43z2xMpwcPTP5UVZT7Qh1gc
Ypuyxhj1laBgLWI2lhpXM2Mo0dLzXRBJmYY8EAMPA4VemrmkbU3pK8EbK1ALCHub
0NQ/sAYJeETcDPDGSwlCflRzmrbs6RnstjRD/Z3wGckOQOPOYlijf18OdTarqvmP
hbp+QcjqXUrQMGsIF6/0bcvIwPAPWkM3kyzpMTz0BP9CtIRIJ8v+zvAj2CJl7cip
Z9h8nLt+1mBqaV3/9DXsE6Gqdef4i55IqyyZsxjs9xMtROmYzgN0gaQ29b3CvRrw
XXw706GLew0Kq189wPL4BL8RaFhZvV1DnAE7f6mo9ucen+ZAQCHJw+vrUr6ZeArl
tDtQmcRTTjxOpQQ8yWP3TP6BotfeDMzWSyusBsgtL3CwBcEFD58SZjYFMjCo2i42
XwmZv2S0DJxUOZWlcS0ax2y4zgmHKG6/cxwD3WgTkBs9JpJ75snnKLblnOgXvy5H
khJgZPC+G9MST4YzT4kQQ3A+tELdxw9VCpdvoI6zQwQBnfuzQaNA7bt2FmPtJP9h
ErnEXYMI3HYn2fUyvilON+joRbh1tqiyvn764fKIuxWQ7RjHBhYob82CF7xWSIOm
VZynjwZJSG1VJeI/Z26/S2BI8u+5DUGPuVXDRr1gS5cpfpQO+0MPkIscUFHXxRQj
d6u4wq3LdVjeM7Xxw5kB0YR9IQfkApdeh92+Vfy2/OBhPdp1PtbUkuEJjrGtypXl
YX7WiFgOBLcoNbAXFP2G0UYnWrew9MrjQsxs/shMbf6vabbikOveL+fiVe/OQ038
EwjoYLuBAGZaAuh6lo2fvU+BKFlpJatvDGzNRrmPVlk0I7XV6ewYOwBEAi2+zHE5
6+qTVvBgHZfR0bKIWC1/m+fP5wwm7fl26Dz8JJ2locKNQ9C94Yf+1z2cd/ReIpVA
2v23c0Hmr3NQY/5QxuWKK664GOnpuOECEwDqQWt5U1iuRuj7kz9mkS29YLgeZBdL
c/Gg2y3rBX3iEqHrIKNorWWgzd3Uz4Kw6LxnB1wccGdaidQ2Nm8Qiki+2ff/eL3F
9qRnHojPmV8Cg2RSNcXPpK63Cxvh/iRXLFMxK4QspRJ3jSghJC71tp7FPqwqDXmC
bOzAktyRkZ3OKOHb2JyhcFexK1NLLslcQZLtqEfTrR8RCTYSRcSb6jnERL7LUn1H
lfz1O5ebxC46o/cTWTRCCMHw5C1G/alC7OROAv1YpLClpGJUcpzGhfz0X/eyU8AP
2ip+aY0aXXuUb11tTGf7xfdkYfTgfcejhN0IJavzzSKWuF3ASf1ehoallvTmZn+A
iXkKEgXCHA9RNFakm9YimCAT6YO0hB1UOHdF8JC8VlvkPrXC3T6JBIL6QqETPsIa
wEDNs/uVNU63kEOLZpIhO9r7Ynvv1MswRedcafdr0oWx8U76pqa1h4/RVYNcSlIB
Wp0JxikBUUiM0MyPOckrRmlDaq7Sc5XJdaU6jfOCGlNj/lwYGjJ4g+USyW2gYq0z
7FpZoKHelsLz/9nvxINuXOj69RI1UcdbOPhW7soo/sKjL9BmSaspPAziXoUG92YC
KzaKAWHRgMiBRJQlsyc3dD+j6fNBlpFFPFfiQUVY1szc6PIpuQ1HLQtw6Z5F3jll
adBTBoqIEafH14Gi6xKr8G7lMG6x29jgzIFJ05fACPv97DTgXyf+aiema08nfnFH
e4JO4H/shwoUW96gw9+o0p7rVEWDHrt62RaVFHwv8+ZhnGde76ZbMIqJgJVPeW+1
Cc1dg8NID2ru9bTRoAL3TVnEXLQuwkhW4IaDmZtb3rfwhwX9zi/KK5v52acsKLD6
bTYAcH1XCrqU+jBs7DWrpopop4KYlEe1XWsypSVrHOBew4MTLO4csh3ZRTPzK/Iv
xINdv32qhUvMgjPdQRFwxcY5iqpQXw6ARfp8nNMd80oAPKbAMKSARQjhtrqnubJX
s8aPwtPTqMOi2ctPeWa+lgyNsM4bDilHb76wuKveOfvEPApNU4jw79rvVRPTTyBR
g6BTVfPRKE57shTBFE3zKytb6RvAd7B6rDj0OHeGftqrL2ZRo7w89UCKvHNVDHw+
qz1UXYofrqqlA0fahuSROSSt6hpavZ5kcgS+jVmC94iwL9fSqVwJPkecTFDBb5lP
9oR2onQjAtmOkjZegqsFLm+f5V+5Sjfu4Ky3kXJ3iAbLAOPAMgC/dngh5HF74Ev3
xlg+h0z3HpaZu9+fACTEmKTdBRcuxf6RTfj/l0Pg8GdCS0YyFeELbeEf6+SocalI
lCNvnxZD/KSxATq7IW3rkpXGV9/kZkgM7HJNd/vs7j6uCscKHFpElw4XOAaOhWyB
vmQF+qtX59bTFi6//PrJB03K5pBL2Apws4RHS/Jr3uYctJCDA0/2spakI8YzswSJ
VRal5hipAs/WDXJ13bTub8KEXlsi/kunxDuFy5NTuEI04Ry+odfOBxGr4VUbcrRJ
GHKL+hCx3jKn27MxyUrdUnjQTe+N9uQvhPmNpk6SCVuZkJ8MyowKOhDlMMqHw3Ac
j/VOhcMgs7KFLl2Aq9QayG5JlrKWahmTFZ4chOMlB4doiCMH7k0NIYuUEuGYRXP+
2TjhqjOZMaEc3GGF5ssTYtNBsYU7bjiilWb8zHswMSSbaPb2tgeXjj6SXIkwoBU1
EJlR2ozDSlPR+MAw6BMKUwPTSToa+GyqpEiBxmeQrF3+LMSo2e43xLgU8a8gVE26
Oj+Cm2S2gZ1RzT0TbQaicQPn6TPZ30/s4yvO7Dj4AH5EvtrNRaeW6oq3gugkrKcP
tjZMLAeZgOFqmwkOmbvKdw5UFdJ3qT7Qc8PEyOPaqvZ6AJFe6xdpbQFGqKj+P6ZB
3R+9WffBKgle8hm3L9npx8vuy7NxreiWQnPNaijcxNcYQJeTBfDzvpY+SHxdN8Ur
HKAQDt4qmMrDCQcvOADNETjLC1YoFbsTFyJNUrtQSAejMl+JA3RzjcTi1F4HFWJV
WwLGiS2iYNXb1l5jTc9av576IdCibATnd1jWLjw85e+aF7QVOX6C6tFceJcWHDEf
7W+Xqpn6ugLzGYDlrGP+yL0j/wQyRKZRfNT9sWT8b+mOMcLFTdEE+TdU962R8ZtO
6BuUqL5BbDy2/kU3WrQ3H22fV7n81eKBIail2DHII2OLpqPcajya5w+YyWPa3JUz
9/MpjgjNXel7qfq/FC9QELkDlaCBJcUNxGz8p2VlxrcfTxxgHV3HGqCvvXE3GdCa
hlIXiesXpxfQzsQct+3WpGIhFoKZFiBItjB2NkpJT53c2OKAAsZ4+c5BkB7bDsBD
qZXohlnPeiGN1cMRUZiOHEcJKaeC8SOt40E535aAr2a4COzIKXsAVTawji8fwG6U
QTDSpQ0X+mg7DrR883+ENrWJUTPVJqsWh/j0p9H49DHueYDp5F2yotW4S4ePGtF1
TQ04suoOtwuOkKjzluudaNttrYJ8ZR/xweR5DVG6/aZhSjFZ0Glaxf91xkvrE4TW
+GYFoERam0VGc5MfO+AIkUnzC3He9Emy6QLkQvfRfp4X5qFSOYtNBKd8nBLqWt4p
k57BDye45N+yHIx7y01MCiSkfq2nb8T5gLlE+tz/YCqoHHVqyEouBw51PIcV2ulV
iRPuUY0fBjhw6LgTwUwt/aSGaX/fSFStwJOA7/BJ/YApevS30ugiD7qRAkcqZzM4
tR8uzlvcC80aR1yVXL1SYLChvZdUIX76toDL/qkpPWboxmKs48xPAbzIcXshQ9vL
hNeREOvdWyHjU/l56jtd0jafKPlyJC0LCHCn4IagjglIYfgZ9A5a1dfLpu6vAHi6
rX7hazmLMhsnAIhVivOlXG/1WNhZiljzl0QSaZTDOe+/w+18SPdMiR2tZCU7I974
6+L4CtDxCEBpf0cUJcONcrMDrNhPFIyJydEkoof6e8L76PCzr1VlTeRBKRc65R5Z
RzMtNkJJjDkkSiiTfYyEtd6LKLM87GcuzHLObuL2y6kj9UYjX7NkqNlvcNMW0Zfl
M9yaKXJ/gAa2nKFAvYd1fh0x+SW7qE8jnpttdNTt/qoDBrr66sp5KqLduPqhPsvK
dVZSy9OH3qBBGtQEnAc8xmtYG0DwNRgMDdvdVp8A9ouDc5ywTHrA9ouV94AHO1bI
S+W3UKifcEz4FL0yaS5GWw3O1alTy6UO7Uf7AEWw3bA1s+v5V2sYpyqYRFbWeTEz
IJRaAd7h3ZffLC1OfjOp9hGlhHZksRnllKZtjqGhjOHsnWQvxZ5KhRCoZ3A4Pwn4
4AbTNdsnREhujVEO9H/Ff48jAb+hC8r8gFe6pjuwxnsfC72OsfnG6C+Ddp/HRRMq
tL8kLBdMKAK7SQXPntwdIKgt9ydpUCDuIYT1+LuR1ikwKM5tetx+dei0D+ho/s9o
EYbDoTjPtBNhbDIbTED6iMsIzAVOxBFve769LBSYV8fNPIUgwj1wvq91mQtYME2E
7zqiM4GReEEW68xxzFVMoONTK1ht5S3ci+iBqQ0pPxiFv5HD0V3x1NMWgFvjQfd7
BuNt7Sh4LbeI+4u7gSjGC4NxLl3kn1GFKj1K2Nk4hc5h+e3G0VUiprmEm8UfFV9y
bsNhSkrUta8QfGrhIiCNoUwtOBNki7beEtlGtev3mSefe/kA+UwnA4K0jW2BjZvw
qpeDfS0tjsW6Sis1VWL9NwtNVZAPmCIN1HCgfCXDYUTn9+QMmNPPlp11mifbRxe4
eK/MVG+fSwHZrz+PeSMCc1DYyb3l1ja9mBowX402+vVBwQrdl1b30pTWiI8BvbOO
jP0tCr+KKQ3VdWjhtveug8AR7xz4sQaTHOcnwKc0MKbnEz6G5WGXwPS31qw6Fkku
SlncHYTDhz51zyL6PgeRrxhDPKJkRwzurvjI+i3qwEDFrmUrglN1N3cQA8+f0XEk
yvpAooNgl5BpbicHad8BNssCDj4if4YrGIVMmc34f93yeWspAB7Hl6smSrUN6lzK
O1mX8YFCTU44BjhZ2Zci9wHaHG340HVNhYSzGAxyUYgjXBettfqnku7pUvStUgGG
0586/pRvd+sjVUuZyCXdcu8KwQFHlodxxofEU6dyrYr705No4RXby3KPZgAzjqgn
De/Sr0aLjYAoog5C11nkeOnOTX9+2/1T/ih7bllIE45dWCeMorrJBk4LY2EGbksx
A+DmozDVnrQjEr4faChqhR/xgJUEs4rsAY5rNOTdf4uA1PGNFV24gruzstgSMBRw
87vrzilRdJS81QFdKhKqSE37/f6Za25MsbMCalofWV0e+NsMzFHcdstduyY6F/8E
6ExHIFrjMrfvWcJGa4TITNUlEIGYPj6waDQy1ct6hCTeW8WWwMxA2jucKfKePqQ3
vCoW7OqZ2Gkv5YbpsCl74dMu5s1nAPn/ajrobeDUewvUCMdOwybuXKwrbGpFkTMQ
A2RpIwNURYJfZ0y2o7yO1cv2ltuRgp2+7c8r/J+J2jNobfMPrTjVFBBllYu+GtTC
O05oicxPhxSKy24WVwhkgWXbKuEnORH/LDxV8JcrM3FIy2p+ZQqVh5LZHC2YbxYR
41kK+2YxB0zssCZtlk1FunAV46JQl5qfrXV91StnqFkqU7rbGyw1a25JC0E3ht1e
6ovVbA89QDzzAkqDKxXE58iRHqCwmkFl7lqku0EIIfiz5xBQ7lQLX8knDvac7ulS
krjP0BySe6asyyvA8DAd2XaBAj0p2n48o8aqFJtb8LEz6qGmz+xS42U5kgVSQ/Xg
pqaIcw71UQ57dZlPaG6SGOYwDgUfSAHVcSMZf1luhTJAum4iHK9HJMparQZ1h776
EjQCQ9sHd93hUmYWPYGhDFxWNBYBn4ZIc4kbZMRWYHQ3G4Bdb/sY2a39V0F9Fejd
vx9bsMg/zyHUFvV2i8cC1xg8LWpPy6D/VFCI/qk3c9pS/Ix8ujArlLIuVG232uf7
Hnoc+Mh0cX4ucfLbiqmMmfewZr7a8XJtgzGvdQWokX2ZDOCUdMXjza1fPAhAtj/G
b+UnUk6ehgPh/lgi0wbXz9MnKb0GKVEhXYwnPnllzTgOVvIZcfGtW99WRlPJqwma
OM8xJNGDEkoAfOu9jFQajQ63Ryb7OTj0oeYwsPTB27XD5ZEoKpGg2XdBnJPRG3ob
cV7rcfa5n8/EvbAAvtW1d+IqsqACYo0W4xB9dFYdy5wc5LMj37EK0lwc+iSN7zmN
y52EtC/Y/w/7JmIUOxuapZlqXzt0Hk+a36hx73EnpyHLxu2tJpaReuIv236yZkrW
cKhdBQuOXojR2hAM7jbI97NIfWkHRzRR1cB8xqqewudupnvfraLZBepPk0YzuGNr
4o2etw+JIz3IbPmcduQISHYhJczv2CA30r0dCzE3eqUPc7Eboz1LJsR8PknmvkGS
gByDzdwAWmQAxvUUk7RLfkkBiFQ1MSoh39g7MSq2YHZRow07jjh004bKWbdkT/rV
3x7M8USQ6Wx61/qe7E7J3IJEqW3GRxUI8jZfxawTMsYQc19Z0q9LpXE9IASkyBwQ
raq2b5GeMIFpbQVRd5kFGeUqogGN6ri+DsupknIwYsx5G03GdyE6Q1b6ejm2+91V
wWJ+JJv1KUspUikhNkX5rfawsMAQBhK0kuYmK0zac7MtQFqbqM6dAf9xSP8HfosE
G4QId6Eoe5l4RjZmi8bHFp9gHMlYYgJijmfJTrgvKN4bLh0Nmor0L+Rdm2zMxEXT
Ft3X42fLbo+9cNImPzLAL1ZKzlkiHxoVG+S45yBIk13zuxg1RGHpShPvq2r9fsJD
Hivt0vkd1gZvWGGqrJRRJgao8S1MwmM+xH8mclWxlIT8puEHuPBOgYCIhUYlVZTu
S49awokTqy7vKH2z8+1VLpxHED3hTnDUTT7QXOqtAf2a36OFCNrPMyTlT6+4HwFG
KO/u8D4f4v1dTF/kyOL7zep+58o+GpIxQijGPJJ4/4A/6ddvl6aG6TFNWMm4aF1P
2S63PkgdFahFJwG6bwgWjv4rV+CCAvbh1cIsUMtQMfb+5RZ1QigVF5DpKoyUC1Og
9lrQPxQ2K6NDHoEd/74P5+fTTWI2eBjWRkCGmcCySJIODqi0AJ6WTeKJI/4EIygg
2ps/+EeKGNfe7i681IinVOEbBsVT+HgfrYqApPwuLp9JgSA411IImzfhOaWmxeCg
U0bsm5BnPW5uLl71HIBtWXN+L0U5DB28j1Q/9wfcQW/firioQQnGhJDHhzyVuXhq
puU7BUDVGKquxBhuFUIA1zIuevAjZv8f+T+sVCbqK13D3fJC9A+VaGxl9lOWFCvu
N1tepIhvXbpJDRrFEebDi0fjy1qfxRyGbOP7rBOR9xL4FX0NZ/TAAqavjNHE2zcO
p7W5BLRbZ733X/vhnmX9pl8t6//RTWVb6BrChZAHdi8erSqKtt5AqZ4pnZjcpejU
YeijCFeYJIY0/4RJJAMMpf9dH6tiXhB1bKFdkhfsEIwEiXlDjnou9pLwkiYD7RZF
afmCFm4HfLH0AP77p9HzNkN1vmSKrXWR1FfxTtLmF86tl+3lT9h3Lsb8aMkkWetR
rqzDIi2ZCtoHuCj2WCWrVgerd1tgWSR7D0nsGPNN1UR8rSPuMIZsIeyEEQnqjsde
Iy6GuP6C8hAzzJVghrAo3hvpxqmqK16mw+SgDrEW9mGscAxuXVCrhBWtok6fRebS
SX33IbnTRM7THyw0RXLUM4IC+JRenxE+miaG/hdpC9slFUM2ZHYtPW3iyz6T3Bc/
XTXuvb7Br7QA3MFaBHCAMM02xUJtrH4eW8j2MOwdKmGS2YFyJxcGNKKpYAhRh826
m9StrGUbAlC6HK5MtyeSTuXh3+AfBFacjeSVHJy0RIL6rcDXDzWa4bgm8hLBfPyN
2R+H0+ahYMOUvIDn+rNY8e+KzOHporY88fBv9ZEcPc4ZYCPG3+/KznqDfhX+TMuh
yFmgzYwEjnVQfvC7ref2tR3p1SKCZX3w5eKO9TECGGTTLZ+hi/Xx78cKVBRxA0Gb
pHcwEBopuo2UX/Q+jsg/JtX0x2+vVadgxQ53xetunAFKF67sURWOHJ9sJpAe+bwB
9zxvw9ypiX4Xf4aIiniPQfGf5/Mg9XpLVEcaakx+PGReFhcsl6mdcdTjoFWuPXaQ
wPgKqK+f5+3BMe4nE+28uOnBY0JzMqdF6Qwo1n6+I+dfTcnQczIWgVJ1jly074RP
Zrn+IbS9QrrF0bcw47IPMHr1byTCLC+BZ9Z8vMvMgYGF1qU0TRdjYzsGFu+6rdKl
GoFOlRyOwM84uhOLYTYC1ubgvfIY1vWDkh3hFaHLsE03jhjrJHl7u8Wu4EPNLPbK
IbSTXrJxJiYnSVh86N7CTYGgYSqFF+KwFwJ+2SJ7W+OR7BwhHL5Dpww5xc836pA5
eO/oNVyvjQpPreXDrFQss0X3jpRNwbhuyVQMXpmpGAvgrhffCcDT3A0Au3M16Dp2
p5AdW6c9KT7Y+6DDJfnkp0qYsYkKSltGeA1IMDxfilvlwv9FKJCVeswAzdloVy5n
g7Cu5k06CF8+Zy2ymORbHxLeiyGDpHVnO1k8HUPdh7KbQYzGX6Wm4kR0jBd82+Kn
xNE9VGjR3Aqifs5eo0htPyMNEkyjliD1WE1mLvVGFJeCZbFTpfECreD5uX2Ad5rr
bpWvmrbdAQTwTCr6qKGbyKdFUuSeSIU3r+FWfuoopX9gTPooSXg6ldM/2GEBrgyH
jjVc/0X9kgEkRwHGO9NtrMfTsv5KL3LNo1rt3EfUAOZE4/jfkucecUnZhESbRoaJ
vcHNdKdn3chbRfw4GC1JdenRRm5Dz+Xk/Lyha/hjmEDrzgsmgjmdX1jgz2cZb8ED
quONL2v9Wv/ZGuLdWXBNFeB1ZRiipVYdPne6YvY/faYimdTefjnLi9+Pt87sMSOU
+K0zaiV1ZxEP/k/s+9TjFGaRhp1ZTpMc/qSiI/yzVJr9k/85U+XldloNqvDKwV/Y
qrnU87957GcVXKDL9YZpTokYollzhwtBKZ97F/wLOHW9ay5DxbrL3xNFi+d32q4s
EIWpetaA851iJtnPnIBO52xEJZhS69p3k/xxIk2wx5CxCY587eFbgksgP0HGtx8Y
rLHQfFCe7UjQZuyTyqm2tiq3PhlcDOulOCAVzIr4utp8kye2drMB9NZZ0FDhmh3A
VvZZo6Sh2cZwtnw+NWoTONgeLbO952XGSJLpNnzk77Iv3preiVOSZ4CFB0B6JJld
72lFmGwQtxm6wKvjmb++ZI9kDMNjeP4L3OwQXnS7N3/Mwt3YykkIydeeY760SOWj
jcre+ax1Nd6xuYOPldiB9eGy8V5v8D+n8t1hSHbw+7wzmNWrOUQU4lw3h1LpjRxt
7LDZJgBZA5Y3kB7MbxTB66HMQvxmG8JQvJ5novrSnqPWSMLNZxjbYAA0led550mt
tKSwR+CjBwNIv2Z5Tm+21kYAyXd76UytQpEYGzzK4ofbC3GEs80yYQV0kfnAwFz3
AQ4ozbF9dO9r3nRB2nWasJFWmvtlYsttsJvRsXFk/p1LQxEVfl/TPPgKTCs42mHC
z9OfFozJ5VXTLMkhGcTMUar7eXx+oGLksbSzdm4Tim2jkq0lfBj2Amww6WdtrUly
H3iXYZz0Bsq3nvzaMmwS5JIDo6N6MkBZt9UPF2INumr+huuqJwAgrdTBinwySXOD
Pxf9plMvqEOLgC49cTR3iCEdI5/fPO7FUyCEA/DHkwzwkiCviAPt5aMZigxfqPBx
CeREBk0t7byHZUgilHZ4b7qtnQXcMzTngUc9EgJoXlWChHPyFA0/MyCzrQ6vbUox
3KJOdaK18Wm1l0Vv+j/ge8wA5iaE5DdAGGnOUateguVpcM0yaDl1aCip2mq2NfHV
qtlRA+olBTOlfx3Rabhe24eiPcrsW7OVOB+pHaM71oQ5dRIVqU0t3eDaRmMQztvy
Doq65Kr9MFusCAIiWqxVR2rv6Nh++W2onTRYPmhJ3enrFjkhUY8vpq4heYx3PdWS
2qQjaPN7YDexr3P0spE0VPZMphAh3nO+CKhKCydWGs1JwWuGOW5OBZXYqv/UGXaw
OOxIEojlPYgm0naPxMYR0/4yhQ0Vf6TbVGt+it5EOVGx/69ZeONZ7+Gge0RmPbUL
QSrDcWOEeE7Xf/1bd6SsJEvKYgcPnlXbhblro6+YU2Q9NGbsiRX92K7fJ1XYYnfQ
Daxd3PtXMszzSDeb+kCExfydoh1yAeTxEMCWOUepURZ38fIMuD5rZSeQZ91bWM6Y
Xyn+7MYdPibfg6F178BEEmDHBC02gBl7Xa5f6O66Y6lsjKL3ppgdVtGc0swep1Uz
POKVKBwIsMuKAyBbmrvfAwOa3zTIM4112gRIiYg8Kr5lIyq/kccwju1y0DAWFyTL
uroUz24N3Svo+tGdSmvF4Sm+33wW92rckwkW9fkY9zGHdEa96SJRKEKC8pH55aY6
JrRM8qb6QVuG3+tIWHbRbuzgXEIJvwXO/mtP6E1vzxWZnECx6l/1r3fgmbfbbTkg
qSExsH/F8Q9cqO2Dk+DbO9T4y85/379mz5U0Hd7sdUk7XaVF1ma6a8ueXj8ZpXNs
eRBXzqkrZaNlnnVATcXPko4/hEUHanD+IkJkiY1GRoctAjjwvL2rxy5ZquM929lX
pYOOTziSs+ZqzzHpgNl5Z6oe1CuM8kriYNEovmMCQN5uZcaBtwv4jf3TLQw2GUDF
XOupGiZegTAcRa/uA2Uk3uYTgCG0vNkO50vgrRPM8smdFDL7vcyc93FuEgMlPQso
m6CTMGD8bYtiM/oKU97e0XfIlsZcr3eQmPh8xfwg6o6VEs0vtZB7NtXGkvg9Xelm
v9ppgPVugHFXGUKbVT0NeTmk2tmUVGpkSwRTJv969Jq4W/pnHIjyTkm+43y546Y8
QCuJeCRtunaZhbQ+kSkMQbOCiQhUXsd8O5cCPTWNUdg5Ul7zHSbV3v3iPcbwK5ea
Lj8XRG1PJ0iEmYyE7rHAsR41lI45V/QZnDTSg12LWTDO/GV6CmZ9p9zkz/Rzip5X
UW3vHzV4fnlVq4IKEP2CPEZkjCqJhJBwJ1+OR/oVqME5camyAspZxdW8iuvHWf5Z
UcAdQ/RFDibihqBdHSSUy46JsDZ6bkdHUVzn2A6CoLSnICwAdlDMzl9SzaxDsPBK
uiAo4mOdwhp3bHW/roPxd8RIdZRWL/LZDiOxuFHRx6iXfmhT36PwgLnKN2w0wz0T
KGV/ox0HUAwPS4lOlixUn7VLQDGiCFoCO4yEndlOsX+RNpz8GaW0zk6pTFeU4Id/
cLkST79vfoYM2hZCilJyM9I0GA2wEliTickNLdHznE4hmhWikvR5N3ZNhUjWKIFy
dTV6VM4eIj2Eges+pPMA4dJ4qB5MVqXNC4W5j4ii7QLQehi13wgNaJeh69iDG8dM
s+hNszXOcMhsG97pRR7ECASPPJoHpnflLzLffEB1pTPkcBq8TfbL7MWGXrSzMU/2
bzxOC8amObCdE2TMlrnGM/KifrlUKyPEO/XmBhLU8P7jm3sFesl0q7/lM3K4aQC7
pOH2Ba053kp2O20HWXWkrrfgCIOKGogGViD6AOJ3OmVzgmnPu6GXiwXJJkmuXgUS
lV7ugk9acBT0yoIGKT+9evMcsKvjgoVdekY125AuoCxs+VnwJ82lsWc7SUtWmUDY
yW4NtdMllM4m+6rIisp09vTTLLo2YkF7e6Przn5f57ZRyWM9Awwg9GQquZP3O3KZ
O7FLB16Lp0vo5tsY2Gm2dkWg/mtX85CEo8T4GjC2306qyi2yGkHbaNFd6+gfIChq
7EL1k+13l4WTKqXVTtjfftFl6ylJqUg8AoXlDUIKoRRO7b4iBqSpJtWzPhJaP4JV
kVoOso0L4mUwl2LR6aOya6V5MdBeXbs6hJSXUbSIw+Qz4Qf7pwhf80C/d8EaDLvj
ZIeQOAmhLuX24XVQugSUTxe8jIMgE7f66WwJH/CVoLVmdm5AedPvRn6uESXVlnVJ
DcsU7K0g1kBk0/gytx71lDR4bvY8EobzyzANc04h9UHZyRCxZdpQHaoiPBtXTMKa
CSeJ6JPDaL1WT5fMaBHJLheG6uprhYcyLWW1A/tmyik0ZECnAb7EMRB3fKQe8qlc
Tb/Jq07pvlxFD+13b+GM3Ztz+e7/Bt4iZf+2sMAtdr/zmYXjshIGw+SEwfeMCOaq
Ym0T3N6/V+COkeFU6bZgZ4wDH7ajSM1yPWIfcizc0lBvQWVWbCHYMOokzl9ufcx1
GLOFYefwkiYbvfAa0vuJ0zYKUd1Fi0FA8lqEz1MtaQTWsicUhaaDeCRHOu0n+3Wg
IMrIIz/UBf2+73AoaJrtc/zCNShTMrE1KkmadRB696ev6xOUhWIb7t9DGz40TzIl
Lcn3dn9C7IVaBnI1oFo051/bkUBfrI9Ehc+AsNYu2Cr7HXZOHhhI5tcp68j8cjZ5
JvIN7VFLi7rb02eH8rSNUO6El4d5btaKZ5Vgnn3Y/PJ3D0Le49bCMO/NcTxQ5ouP
w7AR5cM/g1+tdVsxgajxWt4sEdGalU+x9P/W7qDSV37YID2RUedbI5jZdK/Oq0/9
nE5eV29eBsQo+SP8z+K5GsWtTeP6lPH6D9VyOyhFLkulpaBcJK+kJUoTymOy06wd
LxEVz5ILmYEEaDKUlZts6b5/ZdBvh/QkVBMR89+wD2vOJZwvVBFrNNb6j4K1Cax7
fmERxuiyTKfqnB4uUQejCL1zZaOea6jror/jPqHDFlRSaIoiv25rfIJKSbSsLxXn
u7bZD8QoT7uunhnXlmBAaihcj2Ptk9pKVRu1VsHPxEnXvBH9Q/ZBnMUL2jVZoO9C
wMfw5M00FKgV1ZQbGeCdk5Kbs601V3RCsk/iLvZ1ANm8sFdoMObdoJWPNBlY55zF
tcOcqu22+Gh4o0xUuW22cd0hltA+M8ZLsivFdzeli0YzKpbTx8m1bpoat3d5mS0Q
cUrLh0DTl1dJnVcOphcG0KxFg+xKjjXJs0CIjVBi40j9Nkr1/HVKLEz9AsPIUYQ1
qgY+Dn9dEmPOfZ4OvTm79CgoTkBcI/f4Jq3rix+bTxInrO5q1QfHyI1fAmyFe0zP
h8F2rwsy4nvIkRj2kXe28Zd4phksy6rE6eeiWwHYphJQVurhV/aQ3CS+ZLnRf1Lr
hjDZQezXy57xpDj1pC9L99lWwks3e5SHJm5bcHJicUHaumOSd53KUMLxz4V/vV/t
+rjTB6G0MLjBhwg8L6umH7jL6SUuVHatD960UphIPPul1w3wpA3GOSHaCB40wCaH
nhFs9wLzWXkMV05ZBdqVc9MeuJJlw3SdpV6RguDDyCgjuFE0q1PNogEDw97FPQx7
Tl3y2ngJzLpxZzG7MV90+UJMiOXO8bH4Tk/7e/KWDXqQwMtB89JWhtVIe5Cw0f4q
z0hVNv6F1jo9Oe0L+KCMUvNlGoHu+r/7xMnzsFiHo9s5DCfRfGqrwtLzk4WtdbYS
59n8nnF4S1oKeyiei1nGimCqrsnFAHqaxzkzmLiMVy0Y0Lcb4PJ7pdN2/VbUggU/
ydTjcIHu4nqRVkrzg83Rh77LFNByCcGJDOb4CBgD6DMLdUqB3/dAS/pYSD9MK6Hz
0mm9xPYUcm2j8ttwtFx68F/D+zLfUjiTNDovjmFDA0UcHuyODT26Xt6wCDBz4tBo
qQSIRYuzPEySbxI6+ClWrPsZMK0Nsz+uADUeKCazp4454sOwAlz//D/HaDtarYns
5an7VxoQKBblABTNOzmJTTQ0RgEvXSKk5mZTvvGxU/X77ayvVanSptAvAT9Igt48
rw/7xvYc4gYnTum0zJpyHeGSQdaLGqtuX3STOSNVH1nDuXmUqXPgNz3BTcekVnqv
c/Ypzzgq6UVPTds3HDL02eK0GQxjfU+95qwcEJfbCi3aYxTyATfceoFR6P8m1lAE
HAjsU6GBh+NxRBNk9QVb5CqcL9Y82hMyZVnXiissqhh9Qj+jY0xCRQNRJyYaKwLV
iQ5Xdzhdfe/TaPGTJDr5i48hz+rQCs9e9i1ebNCHP3QvG5MEi6Ys1VpcNjRrDRtl
wZciX6cCw/f/SxMwxv2HPMYTgRYLDjUroTHxqOxhdbCl8uh4SC4o42nSkWgqzOo4
uBlB+/UFu8nSkACYdacs7B8KToIqclSBWqkbo8ITl4uVMwp/9BUQoUbRJBFdwyTl
p7+gO4KTmDTjAKwuPk6q/ZChES+sELUnxxkrrReTGKbD0+ZwcIe7I/oM7EbJi1cX
zpoogMrmeEI0oj+4CE7h1/ZwjDgRLCXcMlzz56yBhXOPZKVx4MBdAe10xhUFTiaw
s/EcUY5JaIrzLFRysDg1L5ppqtHRI2O+eVOko7T41b+yGM+Km/Qk7LiKmC/xCa8Q
tEmNnOq0YWGpC1xfCBIl/269eKvXJTsK7bqMYzUUKKKZ/2LM4fq6Stek64zvpw6Z
Ufg/XwUVPvW9ZwB6knUdXm2BgDy+X3ZZkxb2UlOKEuQEXo8DNsz7hBeOgrgaO7/1
DJoSEO25WOcinavtR0+B6ifW6eTXLlpWFMaAV1R5NsoW8gtV3GnPizaPSq0AjJ4X
WAvqqDNH/nZX5MEu16k17SsREW2Ptb4lQryMDh66GYfQikNx6hM2szfHlA24X1XT
Z1W+DtTzn9NH6Z1ruKx55mkcQ9eIyletVzmKFiTRhdNwPwpSfgBVbm4vdIFvPyHC
XrAgnwE1q7fb7siMi6pXD+EYj9+G6dC1QFML371Zk4psrYPlkzj0KNE7hbiixcBd
tVeCPUKu7sG2KqcPVEW0vnMhH95h/kuDCWi/yb3ZOu4uvNKAighfmdqzBxuF+leJ
mjzcvIOJpJ/LeDSK80Y9VNswIXhGOWad8AeNArg0CFuKNpK0lc6GyBMeCNCoAo0i
56thTvKZJOZQcytCm5VdXFMIas8VjPYkeGAM8xMEMKdwOvG4/6s+vguPAMjWOWw6
/RULj/l+BP73GZlU5qme7T3tIRrSzveI6Vgd4DowrnJH4z4ujQ9gnqFEU6l4PzPr
g1XLp64VESypmdHWpJsNPCYO+fknEid98YFWv96LlOQisC5dzGvHlpoYKsCk/vb1
im7SaY0DCWFlCYXhorPzPA23Rmlalub/sez/xtECc8rEExZMPtGp5SZrzga/qiGo
nwNU6c9sokE3WngsFzGShXG5JjihMsZgZhAdCjgjFhPmq0xLm2EY8AtmwXLG6yRm
Igr9A3InNaJtv/hnviKMHHXNuLGVdblMriYfX4lzswa8BJbr8HiFkGXOl1hup6lz
DG0Xr8uH8G/YZ+xG2B+SolTM5JAuu1weNKOU1dzTBHTxpVfCa3YEaAwRc20b+gGr
5XbnQgwAtIzfLEcTIvrWzCrKgGDeqnatBeW9wlJPdMhkrrIXHOYkNoRD6idvfjsH
T6qh9uC6CKc2Ash3ViWpOwaPimtJiMOcmRmXhUQPD40j+974pEhb9KJvWZorWJwf
rc5VbzeKa27Elw/9gtz6Z/MjxCZXLqssDUwaO7Hu423AHdJYvUWq92OClflgR5ol
PJcXMCvHKGhvF38FQirsibTB30tgMfLtXZmfgvnWxXjIKCgUOfMZA1vMUV8UMvN7
xOA4ZMShG2dUe4ZUMIVcyBK23+7ClP7xAwfiVXQf/Jda7mIMkZS4GAyV4q2iYE7N
PA5T0sbv1zU1i/oJDJdhiw5NmtCmddSgAsOJRpDnz0U912XuOE3GXRMk/UZqoHgE
YTgkZzg5Ite+qhIY2BHaSd/MqU/nSkkkQJOEgr0RDCnB1QEhhhDPqRpgTt8tl69I
ehwGVLb1HdXryQd70NpRN1ISsCnX9lOr8zpPA0JZF4PaKWtQB2SDtbTUCEAcuFp2
XJx/V+0+pKwevN4VOpF3fh0AwrOjqiOJIK5qiXSfOHQfgLQJXZaXAadd8qOKxrVq
HNObrl2QpUr1qJHMys2QLYqcQ6yYoa4dV/N/6iYDIhL5vnssS7IdTzKhKmaKG0in
zKfGe3pSrgCuIsMGNANY8j+C1p1UaUgq9xQmmQYedmeZVd78KT2f0dtmgFYpjnzB
IH6uy8O6MsjMC1Rj9OS8N8gUE3ydRrFnzCnG2/Hzf1SX7tb/jql1dI8Dn1jB+QfB
FH8sq6ss6z0z9f3wyxfPVawyM789EG2D0woj5q78OLjVisujbisBR/EDYRzkNRcv
ooQcOWzxHMUJynrqcfz1RDhIz6Q8oZSAujtmtn8MgbmNlUZpYZIsv0gVHLSbIIZz
TXr5YMMUmGJxszlXKMaASmeSufIn2VyJHgzMcwYrncUoQNLvtfmJZc0/2LINwBDd
eBtfDDvYJaLXzMlBiJ/4dpJRju2p0cbp3GZp0Fj7nf966uiN0EfdaugZJxR9at1G
PuVwLysVjQejfmjsZ5jPF4zVEn5mxtHfqWEdiAXJCW3uGZHknc1AXfEoz2Zh9LKd
fzbzOUUQ35+DMeTrUAwUgZWiaNhaVTMAKwPLDL5j28b4XTrwxgm8RxDZ/L0JyVOM
XTvPFRoRYj+eGm3uJo3KDK5uZjjy5FEZ21jLeA2m4mLemPUKRCG3rU0zFoQEVfM+
gj/xFIqbf2Gccx4I1Ojp0qoZgER2cTkBdCJ3ftM0KBgjf91IDwi7QnRNlJ4e0pGL
hbBTPEdoMxaIb37NTKc2Lkupx/aGIy3U96Gh8e0ru6lOqqpcFJatjPPh8IL2RRw4
MtCkPoW9x7/6C6BNVVHiglrqgHHGQTD4qZym58gKx82ngR0+rdmmFAxO6lzkZjfD
ggm+6b4pmlJVgnXVA6noK1nm4fadsE343zqkLI0Z8sppfxwSgn9rCwoG2A8Fw7Jn
H6u4ZI/uevT6vHKI8khoCQlmNFFj+e/NdR0OWDDP9grwKUM9mUFdi9nzuYnzBc3c
Vzn39UhwMXYjniOdV5avPO3HRbbL46ZVd3028aL9DL312cywXOuvXmiLFvcIOsKd
i4IHtG6LwibabY+2Iv6G/32+WZEOcqZr86vejutaKa5l+kUsMdptcOHc6MuzE/60
fCoiOyLd493dNP86eVNBtHozejIQzs5HXFHXv4IbavIhSsGfAwP3TGOlC1pCwbG3
q+yF6BU3vxQiBkL0tgiy8hwNVhU/Kyer2U1gbcFux2ICmoPDE4GcVtfdqEZxW04q
hkXqj69DmleppDngfhPrKyx0D61H8LpBp63rYUNn4LODn1BJkYKNBXqSWVpPLIcV
uiPNxWndPLz8vhDytIIiomgbY/GuGGBbe9I4Vw5KAcdHfFwrUVRYANycF9DAPid3
DQ80y8sWY+Y20WMYrJNv8ur+cKua3mGq4p2WJRnAZEO5uhVEbgkJDb/gfggXEEqm
6ONPoaP0WwqgzqXaa47hCQo0eMPXhJwJ9pn9XU/UZY+4wObj8Ns3Lh4ZO4Rdoyxh
akwD4iHMNyRNeSdVRhQsXqHREJk5oZQlbNnCeMkxKBWhXuSg5EjqQDDsfySM63vg
dGz4CaPiq6kSOjCJ+TJqgHR1hPyAXTX3/Gu/py8PZLhlwrg02RTbELw7ZweFwZI8
XOUjlZd8EbQ3MGMbGlcu4c/NyzsRFFXcFsUzWnVNHRXng+PlM/p/uk+L4pmkOnd7
8cDYU3nyvZLHgWxB2ZdLbmnDLr+CxWXYzkjhAAc2GLgCNIlputGi4XdgQOvPcPdF
T19yrl/lzjr+7RIjYevdf6WW1xSmrJh1bJTY2pUSNy+c61vyA4czqbI1kDPbEW4w
LEivIDTm0txIg58mSJYtaoKxG8MJOQBo7bEBVUIE77VY5qgorek3jKZEVoJtrUgt
nY7VaL4g3/tQ0QsdGdbIBpHQzqZu5oy4V61mFipaLIPjRnQnltPK99oRE2zMtlEe
5QtX895ZORFay2XIR5r8tRk49kxjbT7Ofh68FG/eOzTX3q38tnJ+Q5K+z96EC76g
+tU14dPIT2zJ5MThuy2jO5efbd1ctznyWffQx1K4k+VWUj6Zk/DgmvUodOj60sKU
Jkjez9aHYQZQe0fj5fWEHd/Zg7/d4YGAiBKFQ9OpwquaK0x6ZkBaQk9HYttpLfS8
CUjKEAyJWbvASAQEIsuI/KcRnhqg1KtNxWYGoqu/6V1aCB1mO5CM6Z1ZAG8UDSAu
uYrksVXsyg6hnjD3vi8Uk21E/VEMTKAkKHf/NVQc3aBEcMSkspoVmW6vXghJZ9/U
xmqdN0Z3GAHFmgorWVYWkSOaE7ZyAhBjqVRgJfSAl1LsCeCDzPArAXIis5FerXdK
qmuNy9a/AhquMSG1oH+4KQ4uh7xI+fDBkTV1XIUt6XTmP+ImtvHNFacKRkXGPCg9
l8Ml5wHnraV7qZO/EhLaMAJoja1Y9ZonFePqhXvLIFSHgaAJDyP9RrV6ilADrnl0
lMcSU9oDj08Vjij9BDsTc8dyZmfYNXY5IC6qKl04HGUkoP8xWAgydLo5yQ2WdHCJ
BPoWTwp2Wps/4ZVq7ld5pAHUQYBT/MWV4jSCDrvyJBTuxUmPNP5p9PCPNOPUZkR7
mDsv+RMAowWUuZunR0x+0HmadFY4oaysic7QTmfbsI+DYsJSa+TLSEUJql1zqUfQ
NieoS5w+mMqaHXqll4dwW2zYj8zoLf9FkoBMdgVAPZ1UhNB6u15nuZkyNNTfgVsW
5q6crfdv4/OJkpEE7cLy4nCbH/jHkCQQLXFOUqwLPeiiv2P8Xb3xNIfk3cyh9APt
dy59EzbK6ywHMKHIanJoFWnfrKuFLFu1bfq7eiOMQ1Ov8NojPzUK1Qznv2MUIMxS
qPVfuae56SKQhkzh/cyrYvjI3IbIPf0J97elYgmSZX61vRFC+2vF4O/nDaL0kbkE
Sp0p8b9LvyFPgNFU+rWMtwzViXf7OEEZG8VSuC8O4TZTKggio9VgNDx3dUqFL4DR
1X3DMLAsRQrVn+Hlv4Hb8sIpo/MkgJjtAXC0SzCpktRRQkiCJHEnAduaDGN7WwJt
P7xwWv8s0SXcwzaSL13UHd8TG0mddhWv9FTzsSrVh/4z2AZBRECsOtXOqvPUkixJ
6WJH0EFeLq9UTxFRGCOny8vUT7mlOYmWTx7oR88898V5kiEs22igVbA2eWqaAMiP
GUrAWPf/hl0IZE/mYKqNzaa1iyLQ1LM/1cSj9/N4iH1qWtgfH+p9iHxEWwYUQRef
bOi2Zrr3PdRGax8n7EGFozI+x9ZptqwkqJyYTDLAQllwUivesyZqAzRv33D75rR3
UT8qYvirpbUaD+tIm4PYNQJktsY7dSa+wvj0SyGSuf66VjIEazIoYYc3wg6RCdpr
+EPlOhrIb2u4TFMeCUWKlt+bdgRzAVeH8tlWT9bWgBTq/yKdHPzAYdX1wYNKznEl
XqFNg2nDtwivYRwBGvnln0FUjn8mD5lDP6zpe4Y6c5Tm4jV7M5JQUCwgiHv2Ne9x
+LUV4DWmPLPfF4I4pY+ezeVkMRZBN90d+bBNfIm/4UPW+iwrOq27u8xQMY/JJK21
ry9Wx2v8IIcAb2hHu94aPn+PWNEuq4G4tbdZaIcL7FGrtRX5f10yTH9wiJbNV/mB
27gFxvhEA9cXl5ZCN626+e4/OfW5F8XccUFPqESrh+pirG/fUFMrcED3VfUzlAfn
TXZI5UMWf7JMFFkOnqdyaKQXhsOLQEyFX/zqDWSyDTOsh6w4AY2cr/+iUSRGHmvi
2h8XprL/eo0zeAjeaKK99V3wSOPXN1jaMlw1AlmLLqLuJCBdjj/u/1c9t8ghE01m
StTmT7Png0DjZJFIUu7TJDCceYCNQP+lPdj0Tu7PizdilgPNVCw5ZeiJtnjyKyfE
f2ydNs9TPxkKbdpHaRg3WcimeLQuSvD3DB+jXpkoDJ227SgnXT8jnjBzzERyxprq
VCXsJ9BRgHNwyb6snwM8k2J8n/Nc+YM/ss4Cpds5sywHf5/FLKENgl5ejBe6io7G
+EcgeVAJDm0Pm0f8fEvm8U9kzuXs85il3K1w9eUcU+ZuKCs5EEUReJ7Kaui/Kpn7
VcQQgz1M3inRu2FZ8t5j3PWK+rIxQkgmlDQUcDF9joBT7TBJxcSzUVnNSMeURy0/
0BZemYE7OvSlpzIf6gAHqoJxPwUwIN9vA3VNPcQkGH2A2PaXuxqmGuo8lugnSoJQ
HpbQqcu4gs2xJ0GJkLp8F7/ZduQsoHQIoGdMGyE+QhOCjbLzWVyqp8jTSNOaemNk
jZ+u2u138YtawFjHJ0liTJBiwVEM+QkAjwqOYDnrxSjSAA/SVDj31cVX03eE38Qy
LYj6qDiFJyuG3EknouRLtcXfoKb7UOH7SsDzs349mD4JpVBxQD0GV6lAhOWhN832
+Y0Z4NOidh66PTs15/8T0dGJiPAe0dxS29MQZg4GbPNBmelgXn4vkmiLv1g32d9N
R7OatxOj+nzjYrYMnM4pwv9zsKDrejMEM450M6qcDURArcW8BRW8/dwVJ/W9JnzW
v17fa+fr0B05dW3572LcTF4ylLlfyWDnNy7DXTKQ27hbbW/lBEx7UZR7rBVujxYh
SLBMFb/XuYh+qBC6Y0zBXjLWa1cVb9azFP6zGbf98hiy2lLDMc510AG3zfISOyy2
tDJle8Lx/g0IGwTCBtusw2nG1EmGvISBEdrSYyqcmbVFhnkklJFKyAyo6It99x2f
tLpUJ+pVa5mAAbGq0fwZmodXaeKoykNAvf2ZXFef87BRlAvvyO3UZIjIb1MVgEtw
gAG49ZNJp5RgLSs3yUOwSgoT+dWHQaa01MlT1FYRH3qXLzv3eoRM3UhiI1aRyota
6xI3jtJiY90NhpsW8g6nKFjvZSr2txdnnoR7/ysc6HOy5kfJhbmhelPF/PhUyPrM
y7VEABKD6LvUNujtchTe058UHCYzqWAPXcihNFZ9K1C1PnDnOAwR73MavTvgq2XE
GJGAfvV9CPNQZ2XyLC7QPLnV4MK8pTUpWv9a3yTzzhksLy2n+4hUzLIPmjq+si4s
jAKzSZiMhDZOovFYINmqKbVk9w6UsaPOtT8kJn+2OS8Bpz3PPhAYJyyGXITqO3Pk
x2ihUSL0dMIeDHEqt2jrSJAm9G5/WnwJl/ucqBscHcSdrzUtbnJ/e+Uq/EhsN/NF
GQOK8l9ZG+pAAeKsiqJYhoz4JS5zac+NRS2H7P7F/jfh9aLk+mw2+6vQic0fC69u
ae7O/rASIrARWw6OoJkOrcbN1fuh+3XZ+SfUYDt6fZboAt1HmXmBxz9Bgjd8TTvT
lyOccnZHqj5eXbKd4AeCeLt08stNK6DYM+L/50mJW+cs+nT/aNS9g+DniZGMmt5T
PQo2WWVGKm+a1qnJUqf1d/7GRSSddtT6vlSNMc5hIsFs1/R7Otr0vXHX4O5A9tfo
O7WGxMtFauFtJ4ho4pLqtCTSKRPdCe9jftfA7DVsc1ihJiU4Qghayj3iEe9snQSa
SOwMdKSNWexS3NfMTQAo/nWbTzB7xLK571kpr5uSy2ZWK0rHNUNy1aq4UHs/DLWM
b4s9k0HR+BlZ0dYWKeihlaBG/nD7a6beW+rv2ISIUAJ5JUm1XoufpbzfGmFaPGpN
4oxEfJ+dwCNYqew+ZKIgm9R7YIJWXh3bnCecnra5gt6/A/fzNa7rvSC2MSTofAyh
F6pCqAW2eTGmw//vDOiYZZeqUJ327CPP7p0QTtoajDmeAvFXxWS798ugcXfyFZpw
rYoT9Yv4T/CNWa4PuCrulCY/2jrlBSax/cG9IPxC9jks2tYYnXwxAhDzQ3H2Uuwm
BYiuThB4D3xWEwYDg04kJA0VEn00hnx08I9umGk/h0uUstqPJwVlfByggDmp4igz
VfLih+hOAX71xsEXzPoz9ZmV2X/Xdr09CjcZptGZet4ZYc7UV779yRFH8Zi5GHSK
Gu7x+uOtVGDIzDejkuLGh9I9nO9XKyvUvau95ErPzKP7UVYZppzFCde66/+o9hA4
syEhCTpFIw/1VSCr1NKfM2RA12Mt3utCBnrdBddOlz4k8NFT28eU7tuCTn70aU8N
TpwiXGa3s4fc1q8y7Yp7zQThNidmT3EGx9bgTg1BcEU3ociIPBIVF3SCnUy/0dFf
cRTcx2eDohFoo21RSO1Stzc7QDyBt/qNLRPMG1b0Bxwxev6epLtuK6hQByps/Tgs
ZYVSznQuTRo8TxG1dmY0BnvmgGKOh6TfpNbANu6bbVX7hT1m97IIF0YfbQhUB/6h
snHN5gh17NQ55lODBE7DSCKDik1AU5lWe4q5Si7E8ALBUv0YC3ncfyAH6XgkpvrW
Pi8FGu0+nOnyGHzcP4b85t5+TjhIQc/LxPyaO4lTXbGqMRfUpI78cRY+ZkC2cnr4
MI7kxZi+QyWDuCNsGJEiqsdoY8oXJZr8MHHhjQ4TVFxIRi+/MXd2G+KThjDfvQdx
f6WkC08iheGMtU4ep+5Mbna3qfAfZRSfSaVD2/KcLrV5g+W1Tp5iwcAQAHwuFqSX
UrC6BjxuUvXz2L82PoGrFAYspLvkvkhLMHhUA1b1nh/cgKA0XsLfB5n1gJzyTmIH
i2hi2gGIe0EvFlDMNzwSkNyC3VXUL+AUEOBMl1ZLhu6OYuc9ofmHNEYDgDp54+V5
TTZB6sy8asiEP1ekwYYF6okYkNk00RAAwcyvYvaIUXXezx0hBa9Dn68vaN11TX1k
GnV//MLcZN0gQAmrwanXEbIomQ/DEEpqsdXQvTSMvG+QsI2Yj/72Ocrc5b/cJNa3
jpeya0wlswkBLzc/+6nrja9PYE6qIpOcyzwMJe1hCMlKA2tzBLEQLuxzc8jVVoai
Xmg/4QE3P7kWkzaSIdXtpZp8uoVEfQFACUl1iEjjmzj5duF1CqZ6/QseV2VHZ4ih
igZjtMJ3XmNUQbsbql+7rwyabtUnAYEBSkyoHjAzEpFBik+4LRSeuOy07JrdRWnr
02Wdg31WZWc3FLzgKu1WVZCcxmZeQZrDPeuocFqrqo/SBnnPi9lcCjwxjWKMJQ3v
/UoGDrDJsneHpFNnqt7aU3kgtfLJq+NJO0WilzkD/Fo9/ANvOrxX2rCg1JpHu4aw
qtWkxRonhLwlDpyL6mkig/LyNEbC0TuacRPaFYtmkyv2Q2wir7ss5OMib6pOBx58
ipjlWaYP6erJNg2arE9AuQ9Xbb/gSmW/+jymYdm/jNfOeXuygAKr/SnyNN8LlmRY
inzQSooTaV86IBnd1XfT03/dpqGRHVFXwSPnTHjFDIrRHWk8oNpkO1i8Tfeq4Wv3
6HkCdmBvw8NQzt7EJ5uZtxw7J8ylX+5WpAphBwmPpLVdUtURdpRNmlNGdi+J5qkO
QJsK7hxQxY82aYZ3ptYFP7cCjyxzxS/M3fw5xhSoAecCZF6bixZTCeNohtCUw5D2
wXb+iLOxa9mlAL6COhpUeJY+Upqj2yV8bXLJckig7sdNsNN1Fw77uDT1o/Qmt/r3
3d3RwBvV0vgcGK9DLo09LjQpYgFEjiwlXVL1zRBMorZcLm6CSfDSTDEJnBahDjJo
bTWvgB4Q/51/eWMqczjR8FZUziqk8dKFz3sKT8hefOByyY0/0GZg8wtXxS0fOhYF
1pMa7S9FWK5LjmFFC9q/T/HVbkiKozuTeWTsQPex7R8XSH5Hd0MOjtzQc5Q4buaQ
wPQS1ql2YppeWJdhFHTsR4XALpEJ3U0kAwdBbh8o7PbysRGFK0H+Kut0/bXyP4K9
ajnEv1Mo6LGGMT6w/JgZE3FUKBvATOvYwtv4QvPNhwtuhYSS36om+S6uET+DvXwm
yNLYF09F0kBepG07qSyAz/Kj4ia/rCwBIhHZoPL5Hmdg/Gc7ZOvDzRdBkaV5lnHT
bVjGrvpv4IHTGyqjw6UstZYz3GgRFqffmG/+yTHcJZLG8S/N5QKhNtk6Xh7NSvyY
je9DGnjtzhHygIe1NPiPLij/g4qC2NCxqi1aVk9MQ+TZoLL887IOco7Gw0pVGcNs
jwPqCXPPPhIU/tzoHcA0x8lzP+a18Y4S6Fmnseq9+FchHwh6whNFMqAaceJQaP9A
R2bKxwoG6+pxEaYh/cpLr7iDW30U/aw+IwVn2cV4nnMtDF6NWZtlFYSHSqX40Z3k
x/yeeZHJ/9NW1mSi3Tx3JfHkpV2er13k+QKtnGyDcABSO/xH1ZQHPddEGwMvCFPB
h/KD20uR0YT/NeecaH/TSWJdjXwt53IGGeqsfjAnhNWhbSBY1OsohlcmZNCzMbZO
bIwQpUE08TQbgUPOCnbKQOylL/UdJMfgMOOQdydaheZFul3l3rfpLj2LIMsyZd+y
YM9QoAz7HycDlYWPgbb56hM3PFWH6UMGOHqEbmLDDx+nbxjhCEIOFDZAYCMGKUJe
GlZEOEuZhQp6je6ixtheuPvi6wzzWiIv2Cc6pMAqa7T/ymtXoG6zWyWT+SsfgVU0
CHKMGKIKNsOD+1IbcXBbZBbatYASyoRhf0/5ihsDqaM9tvgEpFfBDawGkntmmxdp
kWPWWwWAUbTce+7a/ebpknr6upIexO29sS0PYr6oJaHcV+xpGY9u/gtWi38mRwxE
ccmv90SblKvT73xwbKgfX5wg9lNX6O8mD4+TYbNw1ffbL4Dc/jHKYyDzvGW0KAi7
3OHpeorI4za47jSXAvQzx6mKgx2owjziYxDFvcOwliwc+sQMwkmibY1xe7Rsh7vH
M0yfcV/w68+XnMl2ouoWjW8fo16t3u+Q/AZ8X675Eb0uUyersCI3JOY3vL3zZCoM
MGuOK8DQasFq8qi1i2L0gdl1LKP2ddrHMThQTKfOacjwZ3vskXO6pILMnaOUTfQu
yBBIlK21aCQbeK8MMH03oFZWudZ9YAko1VPR8HtYGnf7Ga/17WBI0tW9QTG8NZeU
qbSJgPWg1i/lmUi2YPnE2SI573B16XXrxmZ0byVXKdluFpEg4xySmNns4yPCA26b
EP6YB922Q5yJ8GteZcKY7CaRpSVYsp4vLF/TcnbifZJvw0rps7VfnoZAliG3TV0Y
QGRMOV3/538F3hyXNRmIK8tEE32PCqmbVujcOl1GUPWlM8B2mHtaLHl0uFJ07VP6
c1tZgJDqnwXvq7MJ/g9mNb+aHuANzmHfQc7XTXwFKXFGjy7rMCVTmbTmdxWofRgc
WiQ7OIWWMtYMg38FWpkBnhLNUxlcEOQ0D7bgLCLc0bqZHtvqFFlmt/4dujsbi1bD
2fDxBgkZV6dAAh9OBna0mc6wTLcXNdg70bUnKZBEA1vyivXKtAIJkcwerfkyHeMD
b9wivzg7gbW2gMh/dczyn5HLh2aCaeoRSsat8BhHmtNVoeMSXX4yQL1V1c9r7Wee
rsyddeeWwPFQDmtMK122diduwLIZ6ojvgbe21aWu2rOeGlz2iznC28wiRpZ8SdPf
Rc+wKkFVetnh4i734UxWU6iZow+lwe3QXgIDAr+CVR4L+V3CllhGbmpmHWDiNmRp
eXgrgd1jgQ/I6NBhZYpN7UYmxU9orknk4keWskJeA/MOqD1OdcKs+PENJycXoNhq
iJFA97GRcMNKPWRdbSeuwOuW3QJ5mXqqQxJYsAjl0irhugWLghKrBvN7wjmIs7I3
1tWmblsVhRYLZEXRS534SlliwZDFHZGPO07PI/3CJaEx8IT9arHV2d8CH+wIIDmu
7wbyoWZCYge2em8ildCqEfrhj3BZ+2rFhoNHNeV4H03Pl9oqzteUwXvqVh4wdkk+
I8weLeAiaLr25rStkZBnTokOCco9cEr3Duav03FB9AMAFhxejty2GyyRLTIjt6c7
KkANcoEOg8/FHCzj0Ny3bOlRhWuI9Q2eirxpVIH9SOUjDGS25y7ZpcuIwrgCmC9i
BIItBmorkFhVz2gIiZ3uW/44onE9Nypx+0O4NvJ7HttDpoBAEr5aV81nAL9Vp0dN
PucFg+MXAqwEeOHs4Zu/vQKD9c2UDCxXtEKZzOvW352sGmX70OZlx/odIrlFm0c+
yYPPi7am2IGy7dhoLagQUSe1/3e9wa1VpHJDJGxvflE7N0awz3cTZd7YdPAS4QBH
Oyna3e39l6AQY49RXhyyqvp8SZD06U7jxHIGOwjuiraH45IXXwUmWfNh6EMMGhbg
V9mcBzuyUfTwLr+febddpF2PfF/Povn7vwaEtzLR7dKiLx6hAoH/CQLwNSlSeSxy
7//feZR9Qs+Y060YjEJ0+QdYwKg9pUtoup2CHb7ufMnDWXV3b/6gcS9WjNfGxla3
BSac9a2j27dLGc6fppdL6+KJyyXjYtXXuSSKJ88SDH5YukhsaQrTqDLy6CHLc7r8
fyS9nppmsKzgbPXS7J6jg1oOOeX6S35Rql8j/YyWpLM9iNrgjvZ++FNz2dKoYne3
Dv1gUjqJk+mma8P0DY8S3fix9iwdTOvjQzet0GhGc41vED7tRuCoVspreagdmtpv
b3GJxzglJ/ZOUR0sYU0rbVHLZtCX5eQwPCRwmGnafmS0swWi8wP2/2+yVDkiQHHh
/viy14itmDGiBBeeQYZcAynT82HbnsmGJMo5RZUU0r2cMGCFQbsJmwkzDu6+c6dR
JyEFUHO8L1+sy4E31d3fk9qTFUJvrDiHNbyGS9pr4YPlglKqyu1fuY5jISbv8WhI
YUpJksJvH4RvSg2vgyczdQJ7knEKDYMXs6rD9QhYozt03kX35c+F9uxbYyLCrNfd
MVAjQFyOT70xsESRQODFKE8uYTfbSFlfFgDufGxNmf39v8ovTX1mW/rD6g5lWcUP
tkgznXaGw+7TGiC2vgt1m4tmGAJ/b0ddoKOpNRyYYSOo5TgHeFPJMHI3zOhMvFUC
/QeyEbB1wS7tCaI8QDJZRiNYGqSGoABtLLkbCcFykgGQ/HSWCm7ijz5GzAByA/d7
J7d1bOWNzXRTe8VzInMm2CVEdcaUWsun39yU4opEcXe47sPmAattRfqgxN5DrPBa
rj8Phmv/re5PgSBZXpUXzcjz29dCrSdlzkRRh5sO/MhCLkXvp8RjRI/YiSsJaEwW
+SGWZ0wohq8/k1dAcn3YYwtrNSkuOI1Dm8Z0T8m+INlZ+y8jhLbm+9xtPAfIDm1+
pUImxoG9ox2WkjqVX35w1CtDdVvUB4DxqH2zNUgPhnQw8oteefvYQ0OYtuPWpAHS
XdMABsPqM79n2lkelBE/hVRsGhLKhgq2TVZGhuJ5iA9w3slFMdktcFzVWarC7o6v
fhSv1AZ7EeVsLrTSi7JP1bkhOrnXFHGmj24pZspYovI1wt8Nctc4qbsP93My4j0e
GV3Z0UtmKICyw9NpwrVocILRuGMkQX2jfnWfll3JyMpgBarYFZrz5oLK6FTMMPA/
khKxbUjq1DrXUiNNxhZ/FmWVpa2M1FB9NvMpI/kuzl3K0FpL1zHga2X79TAoQaZx
EIkScppWHbt+H3Q3GMdPwxwRNzB97FPYV0WSuVV7HhFLqO1NlHoa6ObP4RW6A7Ir
LOaVltdJ01YnahveHKqVVSe6+71qHkx22D+yCR9bS/eZK0cRbarEfVhUD0zWzLGQ
qykqTo3z8Gs5m2PlWzCou9rzgh7RHiM/RRf7Eq+GVOA6dC4aeLk1fjQ+xxl2S8WT
xmSU+JeeurDXqN+XX2hx9Mlw6dHeehyoMdfdLoUfHZ03wR5yQkw8h9YRWppD73Rh
BRieZIGQD2T47zVtc0VDsLdnjbSPmKHHCuvawpJa7+iJyGeCnkjkKw9mRauJf3Lq
mIti5gWvwTqo710rSxkvllO3qKurbAIyrUVYs8UaXioygbsGKOydagN3vG7XZmjh
fOR5dv4SB/EfyKRZZI/67fjDceNI5QMxsYWF43L5zTdBx8TgZ9aK5sMbj0lFt/Qz
6/fRIkOjmPuN/Xb6ZrVuKTwf7aCQp6LdPWwp1LUU39wiPXkAgnN//x3l7i0PGiR3
XyFERi/NoK3e91EDa4nFT3kilQ+K459BZAa7kDL9exYDoBQuaSSJY8ErDSUqye6X
/3MMVO7DbhAVIG9wlu/snEc+JCVK/SABNLg7HH5vEiEqK7mSZNX81gETc2GCjEdf
yqHe+Lyu6EmzVBacNqQ5RZjG5GWGprAFfWYYNFxHOWz/JfHdUvXt6XqXr/n/YePc
oRzoyDQxXdoFhX3oIsecwXb1NN0nVWU3QHZjkGKgxKAZX12J6upLOk5ROClS8faG
UgXIYThccC6iDpxe7Rf/JTS053Cr55NZGHTKva8TPiPIN9f9e6AZ/slk/iZB7OJ5
z8gRe70P+36ZjQNtGeg7PsldkQjHwba+9ZqoyDDY6IPapaptjoxA44LG9aBG08Sc
wvuN1Oehz6l9ValiTOXUY53R7gGUAZhlW5up3LFTi4BJ1NDXBsHGM3dOmHpFp2IO
g0PF0U6IzrgGltZF81ldLtCnOiNsYvAALZqPudLMWuJrZFB8z7bCoUNEFGCJ8IEZ
206/ae17Umcw6sF4HKK4a6YknJot+JCIW40X+x0rd+9EtJQcizcPr3Av79AV1oZq
nfoOSKUkVcubc9Rt0Ad+9EBIyh9FcemyaZZv9C+eM+lMYVcVmo7PEV+XETgb7xVo
AaaDKGEQ+QzfnjKp7Usao4qIXDtyAZmnwPtPCC70+i52x8dwvlc54ytVBDalFlh4
2zRa2V/dxiUuOW5r8P82bRFIcZApnKYTnevILAVVQTKJ0BtII2vc0XqgWrgUvB1n
pCLtZONae4nA56TLUQzW8fbVFQecOLB1mf4iFXDhxTPz5ZNDthxcRc7VdfNkEW48
YcOXsoKMR64I2N2Ka0p1OlNphiaZ+cG29yY5QTTYkG8dzVck0ToFlKNYeccBMcMz
t9FwAi+MX8CHvyBsQd5UXSf5KdYtkXNv4W0SLkIIKI3U3vvFzyJT/D0Y6JNPFBEc
teHV0eB6C4PjFYc4sBnPbwingD9EmfeUfX0+fMp/l4AMuOXtNLL+jXyRktFPWUBV
lIO+3kmSvg0d21YejkkcYC0bzPEn5LiKTqMt3GHsAPV1FeKWAKN9a5v3qadm/9Bz
/F1jNjP8dlPCWjRY8GIFkvRWAzTgo8JtPq/pH2RLuSveYaZLMefhyTkolHH9LDV0
YyLpwWbgMUyx7GIAkh54G/8N8oroeusxUInQIa883AErvH3QzXp7L3dBBAba7ipf
VNTujIxGgifUj8NsNxL7CA+1TnGL95+EEv5moOaUtn/VTl8l0lyqB3YFeVSHp6s0
9WuvxjUae1eVld00qSVG2suVyPSEqWPXPgT1LG2RN00+FXaKu4OtbkgxB/R3qLM5
rskaYSEykVx2PxXx4GJ4G3oLknlzP8Uj+zAFpWsD5NzG+I+yU15oOo2PYHD00tZW
Okg6iz6ADG4eb/1XeVl0DysKPvhcjKPRvCTDTaCL4xbBQuwyDFsv5s5aeZW/+MMk
xPXXe/YFtrS7F6+yPjUvD1exxqF/14XI/qP4aIQIBKPcYJMtXUFalpzuDngPxxxg
DkNw4oGalbjRUfO5744GacJQXXc9KFDn/Aq/vjJAHVP7IJLdSwaEgmm8VNE25864
UuYK4FwYgrLtI2ALojHNydF5mYqlo5FgFL83p5YnIkc6Ak9vC/X/OQeTzfMlkhPP
v3IOiV7qIM9sy2hfZipbvPIJGfipq5HvTKnWKSz9A5GwLAx6JwLUdnhUCUoU5uwC
lVzqNOhqibp3+WI7xlpHvnKJQmpuO3HeWnKn8bciAHFOOCWOYwE/bCMhUlZKxpqn
MSnIf84+cmGOuMsCMhZB9w1Nf1pHCYV8uBiAzl4LN/1o2Agc4uDFN8B7aL98VHYz
qhAAdj/WyDf1ZBWzSnSMqsncigJo1dK5UGybwQH2DZd7DYYD6Nbt0hVYcM3RkJdB
jKC2U0oPK+pp95gn3ZhmNrjy2CRMNu7xqinPB1ufeu/vvRrVSb4PNQJjdQG0aHG/
2VJPuZ6WmxZoP/8WcbBALiYAjyynmV7qk5SLhIQbqJlgrVro1+hY2YDmeburv/IG
fghzkl4uPnc508yHk9kqkj/McOwzDrNc28ecxNknOF08Nztf/XYMbEUcWQGvxc7D
6ffW2euu3bzqQm03ugvpjMyxJafz7T4VSe+Shvo+GtOhpoon6oxKg0oM2H6SaKt3
L82DIHbeek/BPWRT//L1al4HRZE3HcC6YLviRobXF4dAI01c6qnvYjPqpCqtJDjC
ClDiQisjIfqlWqnLtbsNc1TwqVTKLv6ya9d+YTP8H02wlpLDH3I3b3ffIhmF6dG4
HSxcqvW0FxCzv/aZTNK7SWFClIn0bQGlnehm9HwohEpBSNd01y1YgT73JGu8KyQc
NHXrLhOW1br3y9j324iVtc3nnfbCDSh/jseTswkfGx41Hzgy7V65PDCVBiqaFUv4
Wuj+PnlqJ/6MRl4c7CC0/AdBVULCQ3Bul2CDVi+3LoxlKF80U5m7YASY+/EnLCXr
wvQseG3aZ3414zol3jqOlW3KuqUNr57xYdX7rRNtO9kjV/feCuIVlAC8jwtKuBCv
Q9UnqmckVVOku4cxWK3pPurkzzDqP8sQY+2mwOvPjhA8bOAdiHH91m30p9g6RDwb
XIxZKp80XHisqTOPEsywPyf+yKxvT8HMXha4XPBtS+JWcJxj3LHy3GDmWd6baLpM
gA9xCng14vzuIULrDORGxyD+NV2AJRlh5mrNbOBN+hAnQdth8iZOaGxZ1jlMOLPm
s1FkpFfGMOMxoKfKPk+AsjpfT4U7vBgoXZCvwKEv7PpouGPfZuh/KwNl0zrDeODS
nsNWYhvc0UKJQKP8pAWNCb05OuMQeGLAnLRq89zx/c0zaYDGj/5uAQR4kKfvVs+t
sVFy2908H0JnE3AapDvz0c3/Z9X1kVc84XlrerS2lD86fhuh7r1SM3cLVIPv9L9+
wFhUxMYaJ/bFrzDdSLKo4E30J5RXPc5+BvzVvTYYj1oKstcPd7zooIyQEvBW4KCI
mZNf7AFAhWKraBZHSuwAT45rMMaFHFX9CmDBczN9ljG8uinVbUrH8docjp9pE4lb
J3HFvExtYLa4dLtlVmI7fbrv55cF2VrbHd41FNzmvxtMvNv3bYMcnsmsHAmAZTS6
U2g++uIAtdH7jRuHglQW8Hrai9MuvBvCw5/PoY8tgBU/gdUhLgDAnGFNU4/LvyHn
0iy4i+LzibEM2tNrqi8zyFfkRTHCbNeFr8XXueW+SChfHYniVKny+24b/1wpnevn
7y3W1Snr2PrBH5CRVgLvLl/ua/eSyKZPZv9ew1jKXesjkGMWj1Kuo8Z3lGYzacXX
6tZN9TsuoEVERk9vNWGzbu59imJ4KJb8H1zCzjca7CAQuBe+PS2yQ2g5n/ug2NFk
gLlsRcYTmmSAYPxJWQEp0yGvpEpaHExwWRJMwsnqANNNKZ4WjEEkLFVMh5I62WUg
/u4ytMSkEXZ/T3mqgjzjcPXP6/tvzCdQunBWT3iUOGl2j8VfHTEdacpKFqZVA9us
O1/85h/FKKqhgwpFaVE5D3fW6xtIKOo0cGjXw5D0BKQbX4Pjd/JufelfhhT9EbOk
6DUA4Cf3LmRmDoPEjyiVZj3HbDSclsJF0nJ62ZvjGxEmS6dd8UIbHoB/T6yX6g5H
P0g8ByZN8ZFBVDOdc8cfYrJVzpz5Hc7kt5PwywCOVC/SLQ6bAWB16Li6q0qekYPl
epfdJmenzAm14bxkPi7qv05viQ8Rr5WJEw2+Wvmnc03b7jTAoufYunb2vVVumkVx
E74xXFVtafM/3C4S+YpjrCTjtyopkVNKYJR5uL5/XEgNiOTvcvd/QlWQ8YyFkGZ9
V5y/pcQl1TbSJXbdB5j0sddcj/y3qmPPzXecYoH/v/YN9DFHs3Ab1bTvBnmTVMib
01Mioqik9i5Ucq0an48idnk2Nfl9SncliwnM/tgGIdJzygHCnowgFNGSz8GfAzyf
xBqP3AZEfGQyGcgY6zKFpOI1byRWYvlNypI6sn5U4tBjHei3XMAi6NDxb560/Y2N
Il0kPn+qMm7PtPdzklye6lOgzFTGEcvtUejloBMKN1EArCFux+7zbd0Z8mQhIr7N
xM14sTd/Lvqgd/dYCwwbr89+EmhryBjSN8v2K7QAkHWlGV3LyYEi+w6to+OhSCfD
TXkVbgbRTtYtvmAsHiiaM7ZAePz9J3PwGgMgOZrGjMVyOnkMuCDPyOqMiMnokEaZ
XsL2IgdPJfIAdStEEgycueUe7MkYw5GGvmRzcZg/UEdWNeIaPxN0miQ+6tTdfR9q
O7IzATu9ZOWry234rZfM0PViyT8E4KW+++GbGw1IvN98om8rm8TqqX18kxOQ00mu
BrqrKYVV/gsJpi7ZzIGxEvXN/qRPZACjFG4OVXXEeMF3xgVDUeRo1apTqpwCsSHy
daY6ualaBVRFZuWEyvl+dyyNL9SZ7wUnCgwMWLMB2FtA13GSZybib458Jt0bgsoi
sykDqkF+qLOaeTsmU3Nk5AVXCNJP2tkpuOEI/C7Y6BfsmdE7TAolCuYXXlp49b0H
dSJNcVeiw8yfW6DE5QNYZK070B/o007iU4aYHQmoi1N+1nktyMjAPL5CYnXMtrE0
ESb6u8iRjMyFFe1J3OlcjP3/HJZUEVn8V56KGJqj8tC4zCWoAZfrbF21yi1ATdX/
PPCtW0R+SOaONoCOfav6h+QYNOc9s8Be/6AQQds21A1HQSD7e/sBu3LH2jpXo2iB
3ciMrygqiHed6FKJb2SggLFdQlqYsylhTamx0DTEg/Oi+GWFSCJuOnT7MCZCEVUC
U7HFEDrBh3sSGTMSyNAZNvRgAqR7NJlb6DPcF9SnwQgHnWMnVxgw45P6VdF74Fbt
U3ru9C1OvqX/ob/9QBTgL+uIcyEM60nlYURd/aWPBqmduh9nEOl5ma4GSH/CeoS4
Ci/PRGGXu5mVkrMhOkbtPiXXAMsymMaX9t8UBGrIpymh+wKf3xzWmmg6JNyKnvK7
/IoW4oO2Mo+JFCeTA8XyisurRVtyZ5eVU9otRrIU3X0eu4qRMnZ3qj+9Nh/PX0kN
y4OBIWdaxZTywf6mUKYZXZWpKLV9qNeSJfOwkhFF78uqWM5yt8p+5rUVGNDgkG9f
OHFL1yi5Jc5fpbO/QA+YOyrE7kfPdHsqUvoNhchmZwNlpETWjWyLn8WVpjGhpJu6
Lp5QJRl7aEWw27wC/KatAnxw1Q+Q8Pe7912tLi/8hdedn3ZMfurQiwROKuir8T7I
tgQG93wIToF7Pzlj7RgKOjIngcvSAp8yTFl6Btl2z7nSoUCokLswZddjtlHBm9R0
JHngPXcpx9S1/LgKGNh6grJVQ8dFcc6Jo82e+PaGciCbcq+Mdsb9CICvmBWxeZEN
CKXp2coordNEn7IQCNHJ+smmDN7LMkKoiZPQ3eKidK3fMM1j//SfMCGokq/CNRGs
0w1bdCuicMJyXrLOuogp9BIdovyB+IY7CQGmpADake7qP5ThuegRDcVP92XS8jHL
QcsmuLlENyBlL9zIxAuZ1xjak+W5KIBCixMOTL2ZGKpqhTin0vfxZodf3Q+AUO3n
ndxuEgoHP/F/tECNc5MXjMY7q7d4lKksrprHWAARhspOC/CP1WEldGwLPCnsY3Cr
HCxPrnyqT/xNBI2755i62v5FE2Uf1cdGJtCfiHgMJuQGFs/gcr/pEYFGwTA6++0S
sUNOKSA6vlAzdC4sM4gyorZSAUrJiKBlXdL7iTe1hotScW802Hd77kdE0ILt0MKD
SyWSu+dbqd7+rBc59ZQkpzlJnNQZj6bF72BL1Ds85/40lXHMs+T9I6ZNRoLz8U3x
b6vAbUHgY0bimYGY1jJ7nBngMkTktPbJWk2Dtn91MPD1FvCtFrLLVlO5db7U4X9L
XCuOmK5NnmHuoyrnpQKeQWmg50Na+uCPqSa+vtPguryuoh5LjmpF5+PM836guRf4
XBKS1vay8RqfGDO0866bE6wsMHcSbV2WZ9lv1vtYALhWRYV/+DAIpiN3NS2I556+
qa7E/762qSxKFP5KIoo9FxTHXjqznmpsSwwF/Wd0r8enwtgT2PL5LL/WWzRsFdfG
JKh7raOipgUmtipJCPN0rCS25bFSE0jYSqqulfelKB3Zwwd8bIXdUQNmW+MV/83F
1Wz115cll7PV4K5k9hVAyWsEPpHevFOecZ+amQXpzXHx5kOPT4N7wqL6E4WtW/Vx
uh/jF/2v3eiG/rs+a8Ik+DAzaQ7fAnBLw8ckR9DJaZnK1Razwp3FE0sQY5zCsjM5
qRsQiav1zRgeLbhr3IhOG+L/VVR848/6CNYAFsqK1wDlvy3QkNNGPyIHYDQGF5R0
H92Dc/rXoozJIO+26UM4tddh0TyGO4j/Sm2enDS9fTRWCzjFkYBplN91DM+LAPMc
OntkC+2AVgwxfDWOI1mdQ/321/DELBYk1hV+qbiFOvB72HH5gFz+j6lvht+XalTm
86DZDY5GsUBgP72UsBIor7D4knfE35MYD0GHcp/KS+DfLMLXl+wKw1LpMEtxfEWN
euA0VwyPPFwwwgEYLcg4hA+A7Bk4pkimMnO3tkEYv0m8btkW3pANlLB/5gw1Jb/u
MfHuiGQNE0w2hG1ZJjFH/iCWHXdGfdOosVSk/RJfZZG59TaagfnUhhsBRKt1miOk
jXdU3ONZRURTSxN+27kJ/Hsz7q0EOFcb01CqqOt/p2ao9IcHNpdSuCyKlqlI2nXp
KjXDOlGXlclhEk0AFnAZ7NTnpgEIulEdDvF8sUAvaAunNOs99j5XTDglBAPzs3E/
lL5IQ04YaaOrBSuUkcO+YzDuiGjw6PN2ox3CB2+5vnqsZE7aP9G7++POpIz4gvG+
moVJ8rKoQ9ptc1NvKiYAUV0hBUog6Gsrz/peoqIW7Fn1Rq3Q3iDgQEOzRj4eNWTj
LK5bQTf7orYid1TH914htQPTrHpk8aLHUXyxID/Yy8+sjWv3pJYztEOpy4FJMmn0
lWGFuP75G5i2tVhb5vw5QBUNNIudEoKmL0QZmVr2y+bWIeWMJbk81+Od5P55YDZ4
Y/bhrf7Tpa9xWrypbotthcvG9BmOVHoHR5Fnye6YjvPn4sewWLDZG2E4LIrU4Qqb
UctHFxPsZ1rs3fM3orcNXBUUNF1E9K/7+8nx9sidG6rItL30DThceAI/NU6qWDC1
6zs6peCeGjeVBCtZB/bbmBBgMGR7hyCTYTM3s3TWZI2QjrWpW5O823Ro+J2dW+v0
laOHa1Zl8VGyAH7jz8t4hRUEIaK0nyYIML7eM3Xn/bZEReNv1XAAzp/VwQ56A6kh
YWaUnLc4pB6N/jHC1tfuV10bpNiwLt9+L5f+gfJbll6a/X/HvIXLJtDzHI64vvJ7
jPTG92RI6buc4DLpxmT+bM5IClNw22d5E5Rg4yJK9h04E7WnaKIfYI3YqahlQnjm
XMK/erNT8v8WyX18eokVjonOD5klottTlZV56BD9KjDSe41zoSm5H1GqGABn5jNq
XTlpxDfVG1pv1Vt7X4JFMyWZyaKFfsWtRQT6ZExjjkonmapZdoQp9SDGmByM4gVQ
pOBaiWNpboQ9Yxe1M07I1LbWrd9gDMMOllreOU4GZK8rxVSYo6Z6N3DqHA2Q+Al/
bW0sRyNoOej7OnLVMon9Iqs1dw8qJiDhOgbGnezbiKqmLx/qO4EuIg5elORODMUi
QAFyeH7ggHD0zIgu5TBCTM7avE8uY09M56ssp4eHiojVvX6Ze2ygRK53t4FbvYyN
AL8imoAtJbO5KKkxogw5j+loT/qDSOah3b4jOwIvg75tkW2QZp6uesyhsEH+ZERH
T47zdfg+N94bRstATZIAjtmTFsSFaFEEeyz8b0IUn7mRvxsMZxClLe2MXRuh/STV
iLZrbfL4eCJHfj2JykcAsw0vUhTqV1ohV9PyOh1veaIMaybkK2sTInIkQA9T2mLl
7gHpVhFnOBrXwRirYFKcIHp8vT/Fys9uuzPK7SERRvUVBOYItallrKtIecnLQ9TA
h8DMdTMQBKZmgBIDchctIyQ0/5dZ122iP7RqTdZyrOUDQsvNy4cQQhyVQXxp5BBI
w3AghXJLw6zkvpKsvuNIJRaohJb9hXmPryw2HS/W310CdDLL+EbJjXIpAp6kOhng
fk1cLgi22mz/LVrWKhSsSfHyV0ngIQ9riSL8VpH9miML16EzKl61xal6vAweA/2Z
BIPTWY0FAETAmPe47a1uWB5XXVNSOCthN3PAfZBQQS1QxqOvhFuMnR5TvzV+OBef
FcN/kM63DJOx5x/QK6KeejVhSppq4ongzJ3RnXnJuEC9K+cSvqSFzdxnmKhYZh9R
+RlrpwoH+bjJaIqK04x6t2MRBzQbVT+wiQF/iKUpOvy2LTy0/IBGblJ7sJKnddNq
Jol0yaByzGLFZcOl97kl8pZjpjS/090oYpW46/Bl0IGFACfOvF2fJtBexf4JECe8
WzKz1d0C0KhDS1Mmjwe12J1EMF8yU63f9ryhv089APHFbM8i5vtagjFj90Dyils8
BxSWkm+YTxVZJHqoP9CK4vzSbO/BMgf3DI1AyDvp9niMuGi6e8hNdahMLIaRRbwU
jXXo3JLIGBGpi/WFD8Vbkc0D9Y7WdICPHjTaHzmKSqLTSR/a8IjaHzs1AovCSLjU
guffdo2I8tP3Rt/hBF4atqootInNvvOMdF/T4smF+6svsZ9/480LaEmL9J+QIa4/
k0B/7SwHBuSWCPLF7dZpij8EWRcFTtD7xZvn2TgEMpIuiv9oQ7ZiWHVhUwoxWPYA
AShEklgZ/aKrH5xYTBT75XchVSw/bn4ePDP7wVXi0R/HqFtSHhnXz045BDA4MmnA
1VCZwnoBWg8V34E4aoiMaLke5udNLP73oLTdiotYLfR8Ix47x3Ht+ZYqDIjsutWB
wsSBq/4BbYCGBGGyfnIsx23L6lGVn4meAkfROMmxGGZwMV+FOHMez+yQO/DxHQ0v
GrqrPWWOTTtiSgtBSu6x1HpxCtJp5c4oivTvv6qTVEr8FaMokGFxls4ub6tYu+TP
rg8DpnLDC4n9OCRD3U0tenLHxzPUcknG8Qmzez5R9P1MYSsVrh2zEwrnBXTx0PB4
SHbubNvIJl0ZiFYfWjkbsIWQ8rg2FWAAyfVXU971S0MpvPuODVvH95bIAmskiOi0
3ijCbt2jK+ZBjh0NEFiexKYQpPAKQpaP5/5uHqh1sByLNfvAOykCd0gbt6GYc8Rz
WOJwLKSwECa/F6HeRbOYnr/PCYZ2petknUNWfCuJpbD4qvV/CIvViF1F/6iFkVXb
zWmGY+hoGZj9C3//d68v0C5nJzQ6fEuQK2RjoBNWG0NPyduy1J+8Fh+02Ki7mLSd
BbYjm4u5uF6xrSZHk3Y5J3Tt1w71eH85NFHCsQwxaXZDlJZzgfj78C4cqvQWS3Pi
6jN6bBqpVGb46iSWxF8I/R5TRSed7Yd84zSBwvmmfHUzUNbyGya+xiwpk097EZt7
uhwqRbaDw2PPjbCLKnNbSMXbbypAPtyhpb6MbHF4xZDJflAonnKfWwVKgpnHSfWr
4xSo/K2VS5EfFPZJzxuFIBRnHHsBTPh0YvuI0shaN+kVRgO2sKeGJnQF8Rgna6ZO
7oZpYfoWk7GKjzOPIvft7NN8iLqZDWAH5P6Anv+tcKa/ecD/lLNlJqXUiIDWI4rv
zS5rWIS+pbMcyLj1af79UZp+qaY/MFSSJSDgWxBGhoF7K5Yy3mvQXDrfRGutlfn/
eR57rfRUKEcRaddXRPp8PyhR5BZFOzM+LHJwXRMvP6ifrafLFdb/wRjTZza3A+Ba
5v45H+w5zV4WrLbFM5fVznTvnL4D5eq1ZFWszC+CsusAabxwX8DcNlvSWFpr15gU
mEVENK+Qj+LWilV1cOjvnBbJ9O273Zn06JEvLLFQ0E8gdt65R9mkPe1cwr0f2s/s
pDuLtgY+HaDmpbXmLrY/eBvps48nmSiqWtEpMprwL86ReGmr53OL/L4EPWX/t+om
YzJNwveDt8d0hPgykRWdH6kozjpTVyxSoKDmnzKkI39sia3G61ryUNKuiwwhKikI
NBES6bl8b+W+FA5RzzdbJFgpfev7WnUWtB59EmYDySa52vEWlVk47NpeX9ukn9EH
L0GqnbPwn9+HQv3nYWnkdsSc6jcaNqGQjz9090QxywVSx1ljmnTBP95AF049ricX
zfqxllLATRo+Vfw6eya8YY14ud9a6WEFN5zXZ4AzElTl+sR5PwMormdDsFZ1yHMf
Tnw5zzYm5wL0fVb6IBrC2kTSOXDcUhiR7TPvx0/9nQkGohTm6D8Lpvo+8xACs1Ge
127RyV1Y8ogZbt6Cb74edg==
`pragma protect end_protected
