// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:45:25 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
m4H2quWLfKa5Ta6N29RqMXWsb1UqB0IAUa0Rc3b6u1vcKfHJ8coR3MXvn8djYg43
x35fYiktYtVaJEHOSIC22HbmvtbP20SgOZZ2UU4akqzyu/LsvSfF6N4gN4N2XKCP
Ep6l5+/3VtLwrqY6aZ9xrqaCLhPDLwwZdtZtbCde3J4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1488)
rrXyb18p6eS/ymxhf+/+nLHkW+A31+/zuBeFHkVag8LjWGbMviL1X/cv+xCNBlTf
C4bbgBrsBRNhZzmP3XLs9QLYCCJWprB+LtcRBmNjiDcuFLUwQaoty8l3sF2GlNwn
p/hd/BLg27PnmajCz5x2IbTyo/s/MBr6HNd9b/Lntro9Ti82AqPS8hctknSiULEE
edCeUFq/K5cSfEUqjd4mwpzt7yfBQyArqI2tH8NsOTGDL/DSSRmOaQZSXffloQRU
aOo/MG6RUbDuZJw/xDe61cBaxODf8uMowK2txfm7cW1JgaSKNTA0CgLPYwYbHuN6
MvLMQ+PfvMliMWO3wmfttW/2atoOYJbsWMaEShBTS3lUi5fXuZT4O70qJJsq6ODg
eGTVQ/3TOhql1sc/u8bKBImkqmP3IZY+AAnU67JeVHJDl+6aqKJQiMWO/K7Omy/y
3IIJT/NEFMjal577DdME3tlqB6Ns6bxzEati88OnXaCMjb9wq8VsN1qrWXtwi4LG
Yhk4TzLomwbI4hUDL1Ocnt6ijnhZgZ3qpFDyVcO4Ji5yU6PW6qIPSBMRgj/vb6ri
i6ao7zIZrWHpqGPk++epLMXUYjMYnHE3DRgRW/NY5IgAzgRECyjBYCRiRNrq1P6s
mL8ywqC2yyDiwSp6J1Va5p7tLENwA0JjY4VOPXwO0sGfQDkVHSJSS38wSmSEfedp
M7m8n7BiIkkeUe9sjDBrWcEPcE1YlOMkwA2WuEWP3bMw57vTV9eP6vd+bWJmCn7C
2KBcz30g1IBcfKdFOy4s0+gE04r4Q/VPH79MX7HwISOLdw84/G2Mo+vgcLauJwVP
P48J/XLl5NDq9eLYQgWDB/kmsuLZKPxTeiXR2QzqoVmiyQQkKo2UVioEHBz2QgIG
HLcK81DrXFibk5b9+pnmtGp6CFZQnwGzh24nHqCE3bEVIX9H/fNb9WROaM2fJJ7L
JfEK3NdHWcvje2a2RROl/GE6yZfFIVjIVPVzWXBfPjz4l/3vJQ1QkpABwLtSPpXC
QtyPf+LYvJTx1ykHuCLZrXnXL31h/i+Q/HTt71zdeRPXQ8AbgYlIbBA6WGqNPeeQ
TzhDGIAintIOsJuqPUGeYUqaVfORuWr2UjIC44mEXR18BDADKLyHuKxgV0hkUCYN
5KlQD7Z4BnwqfrhT/RUmvKaCm1PVd2NpA1oIhYxyPrulkplxJrp0B27rGT7QevLW
p+b7Ep4lw7OwY+qZWoW+T7CUUGRongbNMk6l+RSief4jsWrI+0D6oR0RhHcOq22w
45o6G+bx1wfeN5PngC5wzog7qib69Qvt97FzZJkiMhfnZR2Q8WeDIKNl65SowT0z
IPqZIKDstKbuQw9eNUfgfGy10S1OA0OuTbxe1sHlpRe+DpaPuoO5NN6uqJ14fj/m
CxJUOQouRnj0CQNEvYUftnkPi2UrXLxX5oQtU/AguvrBKsQvl7M+aluF5QqxxYGW
9IiK0yJMNTlRZCH+ERI5Czg6xzFxhtDK85Y4NfiSHA4fxg//T3hkgutzNtTJivs0
BNBYrHotEgGCVmVf4lkxaxvKm+tpyVIHrUeymdmgqeOeHe8wm02ZFsg1j9dhkfeH
D9htyVbytVnvgE8cvbhRsjhmS/NJ8GpbMVWZCvH7nV86TvowwIdAd2AYegwzZCAv
VhLdoj6/5K0PabmNh6QVPYdmTlg34s1szmoOuyHzYuzuwQt+N282yyFpqZssjFwt
jnWaRiYghK02c/jWZ22PjyxMia0LXn/tiRqNCq4+2AoJR+/0/37wqC1mKgkcz4oh
YlIx+vL8wVf+1WLl1zBJXiodhEled1bNdSz6+0evPaRTirQsrtbpIpZ94UHj2hPb
77BL4jkF7yk0r6IR6T7QIDe/YyHW40/GtuTQj3Y0iQvuOpymtndndiYfFP6+qa6/
94j+AdbaQlSoXrJ5ofiD2ZVwqm4UyYLGf2TWCm3MqKmwB6Btpz4lbN5VYeEvp0LH
`pragma protect end_protected
