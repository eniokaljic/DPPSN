// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qkiud2DgO2QagNHrtSajhvnZ4TOd8E+pRNQ8QaLT/+5gfRzjo1DadT8P+L2iHaTs
aDg+FwlP9f9IDc0gM5hdbQX81bHUPk3bfMJ3+/cZyiNLUgiePr1JJz/iT+EHWOaT
Npbsh+1/xOsBf0XmJNawO+XvvD2WIA2O2NzUvQGIc8o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 180736)
A+NqsmPsylzozmeCCNeZK4xMbMAxM3YARUMJrbbA50P8OAckPZ0u3ZTleqQUAtbs
4OjIcjdse1Yea9pJLVZfRG/0bct4M7yb2biovdKBvecvhqBrKmF3q9to/n4rpuuK
byq5cfs0b0r0b7QqAROPbVrWl2MSyZJvG1a6zsK663wmG0QT37sfvf3ApwSsnODv
wJR8IhvrIyhJNHyBn8uqa5ckEGOMNuEeuD67heGz+/DIXiuQoDysvdo4ZIzSB0LE
JdwGQk4FR5bWzTm3gDEu/uRlU96LF6m/fO6TZ8OZoLrSjDL1vpN3ZXN4OeBjmcnk
+7IwhI72RgbgNPP0K3k4xVXbAsKh7jApJv0SBo3uyYEm+zNqezXcOh/4eY2Xl1j1
7nu5MVMGNQfIqBb7dNnBgv+S75VJUDlld0ka2xcWVf69tyzIPi+AEw2o5e7RKq7O
xhvYskS/jr64d1FHpQpA0fV+EBHv5ZgVrdpvGFhMZU7sw39uxJdq7LZUiD+gy6Tq
+Axbn/smX360OFKNsAiPqYRliVYgxSBgJZzXWqlhAbLwqTQsX0oVrPyQ7JcEj1h9
8/h/W+M8SOneqNTVnUNY/Ib2foYiAKgjQ0ZTttzDSZZ/yeR3qdtpETSzCl1qQ5q5
HuShxdz5Y6Kfu9eBzVHsNHzrRTK52gAPUbK3j8bkzIwwCPnZuOpMfcc4cmwbN5MQ
kow9stxuI5twiT0DH/iB/NMfnE5PKs45//SQbFliITMQSHIvfGMmJC/ghyBYPxTH
YzRdPKxCezFH8p2qrouPZJRtjOSM1cJQcymlQP6K8JHUjPDncKseBJWusQ9Rp9GW
SxGvIL7Uv/DjilQvYrXDL0nvxbp9GqhUEqJfU1NucjBZrldi1l8WJGvbQ0+iAqVF
p12Qu4V8gYECxP+5tyEEbcxiQ3RBHahShyJUOrR1bqLGgD/OqjPwKWEy79Uo2Fml
lGFl8ygo313VMpfY8/q/A4jxMPOtTihnJB7+PHAK1zqjFMOnto40zbJDpiO3rW4w
U0ZBlT52jgj6/kJSzaNP2kaa0Gx97ZWc+UdHN4gyuY5hWnK8/OVEr0eZ4xGP/J4s
I/GN03q68c+7a6EK7HsyUNid2ryF3rCm7fEWB0p2X67cLBmRLPafdkbSlH/agyG1
pvGncIS0H2jB5/r6YCKCzjqrcNhTW8Y30Kpn9WosxRqGt/AcUPqJZZkGkcPqsZwM
rfvdHpP524c5qCmIvGDQ1fktC8ig+7q6EhaqW9shrQnSWwh0+VaHyWvL3GvP1r1I
PUCzJlxmZ69vHfEwUtkPmwTXvEUlFnB8p+OwG5JkKjbk9ocHUyny22XGGc11wwaO
3jhekIXz8U6er7DLs3dlb/qF4Dkokwvy++/0ZKtqPKYd4fgP5AnsjoKes+ju0zSU
zIALi/dsBC8aqsAxVAW9AUot+jAC9JCd9xmACcc/QP6iK+rwjiY5xz+HQsTz23eO
X8GrnZgfZ0r1hKGLxT20Pgd27yNKPzKxw25XzcG7zhGlK0IQbvxWAUEw/0MIomi9
HCiy7ev/RBzRWsNCx2U59bh5MNN5uJ9d9xKewh1c8iPVHA+wpWycgX6z4+YUsReX
jiBTmQYpK/vi846gJiQZga79hgF4M+XjHULDohH2UQ15YqcM6jJCNaxjUvNjzsab
NebbawptUQjkpmn/ZI3DxzAtxpjwNjbrorlKqllw5gRvjtycEKIJKXlLCYw76rPv
EgF9PBs+JiKoPJx3VM47Bgn9z81a8epSXCphjDrI1jdXSRjxJBTLMGfXDQoY/8fQ
DS0Ii3vXpT0YswzmK/0xLQCqS1EyX+f86zkjEoVyNXLDb2JjVxWDcPOJDmEdZ9ts
bqgkcUNYT25FetEGoHe09PUrYYLkosGMCJ1QRc5dTJ7mnKUKiUnBBV11+ph8fJUf
ZpSqLBzs1ZV9Z3eitWurKag1dN8zBizNus0qUG/kFiz7+ZDnhsDbiJ0wObplTYoj
XtYcEXp+v/d82AQgadYp/gR2LDbQLs45WJhXqom1Rk5aC6RnhUIInYJUEwaHCjIJ
pYj+QR+s9SgDmG9V3R8eTn6VlkxeL7a+wBMDKN5zO2oxcOv7bRgU5/j4PNfjZ3OV
Su9wpUUagyX26Bx5JT9wyufu8mcnkJ0YHGX4p5t+zNlvSArMbgUxQV2yhWgPz5dZ
DQaY4MxedEZoyu/Qv1c34EyeR15hDuJdKN7uiNcZjspXze1Of+DtxL7lqAqbaoo8
kDLI63mhgQeI34TdRVDMzOXMtIqHMf+u/xyhJXgZenaSvydjSf3jJGihb2sNWdYS
dZ8Y40acdOIdcQ2TSN1JnNOwH7yDV+N56DufN92hRmm6maN/DCk01dU04fsMcUv9
AN4p2eyLkZyQv595ehETZcu+BsKaWVNX6U4yD+xJUIp1SIxABhQbweFywyt1XuAo
lt7Z5MS5YgVyIRc3CURQZLsfIXyn9d6f8XJQObMiBrMrzd4CgW1lbYLitegcuai3
E+EmC3nWy/kLjlVN9gpuj9jzfoqttupd3UTHL6KcS8Q3j0VNEWeJPQ/KzGwUWRDH
dsoKxBLL6BG0UYb8dTtqEPMb4G23k1nIJQZd0Xi+MHt0nIKLvgdguSEf3AKkis9V
dcFDmVqIqOcuL6VdLLBnA0W5DJYNz1ghXVHhYV9rfgT8ugi+wVQWRczyeaefgSvQ
dUMTF3Grx/LGW5KxydiVatO8HGYEDZTK29B3ujtUBtphY0V7k+lEPpYyatqfeqvC
KdmBhm9oGEm4HscIfGM4iwdzFqDVHubRkvt0f6rXX0NVJCinq2KOu2VObn41eMVc
X0+gqYsO5/1GB1NhGEFkGfaqGTVIIFP8AhYX6VmtZ1u3Qs2Z6yDLdfF+MGe2KZi0
QtSiE1fjRH+oQbGeVxBHjKvmww4QQrZJvpDw5qp4LzpZHFgv7HSZswwefZXGv8Y7
VzcUyP0LOzAZZVAJbI52fxzb4FQg0zyhLuPaiEujlczPeLY8xqCcie2onj3eWUG0
OB+1RN9JMu2JayyNs1lqDN558OgYKXeJ8sQ7h8SIuDf0tZwIVJj28bwC226L3NMl
MBp+MutSIP5Y+ef8XhLZ+dZDgocz0zUwJ340AVZq3s+r5WRjTAb9FzRIBR5Qc4IE
5+HFT9ZQbpe1lezwJHRZylFbLuXXBOHrY5HuloPIZrWfSQpm1okOH/Ibu7bStZX7
Z98pudLs5EkV7KwVkfnm+U53Ahojv1rEziE+tagCWO5je6Sk8vHgJF0Lnl5zoMCX
xNUWp8izoHE5zq+MVuLCvlYQA8Y9sbR6CWMv6aYbySXXAxcjF0BoqoSZJgBkVWvn
lUYuXzHb3CH21/LDycQdL2VpNAPaTHxBS5sIidTPP/qyAKtadIXQdc4WGWGOq57l
nDJ3/XNHGTTuVldq3dWOuCVrOLUPYebwBBBdfFHh2wFeArIKRGcUIaiKwAuF2hZ6
keyPaJzGvWqXGAiXFonA08ZA8/QMLHTOMxZhot4EU3h+GHNTmjbz9CiEwfFq9wu9
RJWd0ZQfORiH4pFmp0KmkxEns3QLSCLMSCzk/5k8iWc5KoU2n6AQn/+ZFjlpH9SN
UqU1q1Us118Zc86nc3MKMBLlH4zoSnndhF1eRpVG6BFPdAIW9yBXDjBMbILwmn1Q
2JrsjUaS9zogounKLxI2/QxeagNqDvnLZXSrO38pBR12avj2RMoN1SjI8YVDEn0b
unkM+sT9P3eAj6cO2/pUdTxFsnn2ksj4XenzOSIER7dl87A8+U/jaYEALIF+/dXH
h6vl+7acBZd36mz31z605GWCR31ow4XVeAo8mjVKkAN2i8isX4tkZF51NjU08QmN
7aSW81iPG1FNhQc/pb9pC5UpM+PgsYluyYBgJ+JRxQtjSR5V+GtE8eBj8JpAlp5I
fyLZmYSavppQmhMSuoweloBxHnEvk6t5VctXFkvB0o0ITFMXaLZvofE02FlGtikx
3SzJCAqZIBR7e/rLk3EjZxAYnumIACzC3kVDKCna3W4oMGrGRNwLdZ1jOHVupNji
6q9X6Y50XGkkcsfCocHaSIHEMMw8/pR0Y3ywbUhrJBqCrV10NNvXYR6Ji24VxQ0R
qOhQRwmxgflMdDfDEvKI2TBb03VQXpP5998XScoOJ3U3S1E8WGUcwA5SckavOfyu
YrrFnhXoDs6KIc4TztIh1CSybadlhXhDJvXMB1hi3nPOI7Pw0uXgqnQpKiw2Do+K
D95BBxw5haJf/f2nqpVquiFLC+0wHCSLeUz4JHlWHL0RcbnEfsgCCy+CzYelB7v7
7gFcAeQi+wzHA95dexJBruUVNr5BfNebAtQd0melApZAZB3TMQXg5EIYS+BchksM
o9gD32ugjDVTEJ6c81ZIuOjgr8Iy/tnB2AQ9FDpXZfRBqHj1H7TaL0fyQNOr6Pfv
0Y3fKwf5e/urTQ3AUIIokAK45IIHwO/frdkOUf94lKU0BYgeYJjyDPqzb4eFPfbo
I6ZSqA+nkiWrXFqLE2f7TQde1w6E9J1BDi+/pDQ+Kl+PHfI7xc/uLyT9Cqie8g33
EtJLVKigCt37KjrT/ZMmTX05Kmh+gTonXQ211CcpA8zhS71QTxkbKWg75Xqjg31z
dokGL4pQ6rwg0IYzaaN/qdx7WzKbfKDG+V5s9x+wWbu9w4hhRS4bcxVyUg9rAG0s
mfKoqyDgl+JFP+yMIPUbg7LkCdIkiYfoKVfUWalsdXFMorsNs+TQ1uqGmiwDKCtY
SF1DHk9dnlhewE2lX/IgS9ZCPZWdwpUDadrP4C5C3uMPhJUQXwy/Hu63BRKe5leq
NrHeVWJrX2ZCtQwBN6ojDGM5xONLQd/Tbtjxh9nOMKk/cXV/dOODWIxNJR7ZiZyj
77yVEMUJoiULg0UPe+61edNs3JHTNefw0Y5/S3S5igmUzs0SQewKvQI56dTAx5WV
xvID4PPIfGnSRlZLx2jL/CT0mBn0IVq/SFOu8QJjxU88pUV0qBfJaKxUGAGv7xG2
QpHqQn7S57covVXCmm7RL6XZ3hVpdOCwmH2W/n0bSCAvPjt4Lr0xKmwrcNUI7z39
szE+2axcQzfv4eRbq5ExNXDnTGUcnlHF5fVfG3OMLf2p2/IkpovRBK1ycpNoNzJp
PDu4jxWQIMKe2TcXBt6wvcLNMqQa/LdAqjh8Pg5Yz3dnUwUvjW0Mk6VJMmFJfIeJ
kmgitKJrTVVrBnCIBwHYJt3K881hJNpvcgnV6bpz9RAhJZVuEQeMCOPww1cVmi3v
BKRbHnzdQYfS2StgFYs034sKp06paqyvEXzVSrSbJhvgie+r1UJXSoNp4zm4rOrn
5xGbPjmHLBi14lGOb0xtBDYyiqUqbTmlr4ej+9uAOO4mftumz6rY2QCL9mAQtQy9
BfiLJJku4K8NqbTIwzOXW1YHIZbXElDZImXLx9DwzMLXPI8iT13LaelmX7ux0F/z
xX2iXeNAnGXWjNUMeKcZOGN1vBY+FT3ZfssEDcHi2Xr4Auya3VuP7r5wkQY4Ph3V
b6w7uoxOkh4G7O6n4VXUU9UYDNeaGRJxGUfPzsqi03GZGmTQlleS5iwJlQU4/lFM
+UyBl5IpjVDaa/9KKtsWjPaKASF++fen6hI801yDgMYSRfvvXUrfJE+4CkZYic/z
7D+cIiHlQIyAPimYgWKQU3Biy1QVHI1P3w6APesHhvu3Jv0MxBZ53H8qOG3iAOaP
daJsDcrh5QNnuuav3dk6wcI33azOLVoXFU05OJw9CiPMxvJ6ERYvzFCpvkG9pslh
7eULA2Q6SYDWcCDIh5sBcVN7uw+IACh3CNwlxxODzG/z2QUdlDUTqeVHUFy4xAuO
Jc2fTXGDc09MMmwHknPfMTLhTtbaWLrSLq+22haSfy3ejITT7eZLYp1x/cLAIRLK
uySLSaaNQdnLF+9D5eoLSo683zTtvHFeHa0Tjrpyxr8RKnvGxSejkBthR9th8u0/
MDVVJbFTExmRHZtFnchQqbbyWRUR5Q2WFV8ZRlF8KKXNNZ2ypd14FXmuvJ0uPk6d
P0pX855EUfKlZD6kyoBM1Z/xQVmm4VuR7laJu00B+DrNTPKPAsdDJavoNN8WQ3BE
Ms0O3KjtwdRDK3v8ES++FnHOl014wtjjF1bgggO0KUPBR4NmxkQfMdoea7uhtHgz
RR0yT29P8lwpr4SKkNM7nOWxuCWTbpW2MhHtJUoPtoTzw4LLisXKrWDRAHipWTCi
VUGZ249vg0XpP4zHla+q9Puw4FLobHUyvPuj2c5C0c9faKk1gr23kM50fyPbOz/j
wDUV9j6wwF7alU9dhXzFhx4aYDITeMocKiNJiyZKdm/62lRkKnUJItEKAQ701dnA
0sE0hJZ99rVMifgXr4JJngVB34nnJqFeXbUju58hTNEUWmP1/53i/KxHu/HInwKB
LqIQLY7f9+b+kfiNKQcXNdrHiQQ7hoUx2CL7Wc04tB6XtFlzu56rhS/b6inXtvDz
R4FYOSz/m3uwH7JoOAy4egbIGkjmKG3Eyldb3DWy7c6Axwgn5Yn/AJJDk9YdrAZV
ms4KbGqO9Y3nVdcX9pt8PFvxZzkGP9SH/5HjYlvKzm6k29D6bZ23T1bkwJL2TFzh
oa9pF4agR6SqCj8fepBz8uYoIterma+eRUb1CmoMN12g7Fk/bq/wrPMEh8XXDFyK
tX/cbbnWV2hcZUzXJwY6432R/OUW0jS1vLCC0LvDDBBbwYDOOukJEox48wXrJuzP
nYnYfF7FdPFIkKp/cPu/5uWhbHbk1VxTfsgeBRl2DHIvw2oFeVPKf5gcvN7CBrSc
T20eJZIPhi893Apbm0wjacGDV7S0vPW+gupsduWIJC9dyo79OJ6BlN1Bl8x4W0dA
6q3gNtq4A1H6tzTZl/l2QxVQbNrizVppj1tzvU0HciUjNAAHywR4DIpA4FACZF+I
pr/1LYZi3dQd3xmA6fiDj1tMa/w4ZZrAFvKDyg+EcrJ9iF5dVXRsgxVuWrsWNFP3
Eq5oPND5ZOu6Aq3/Bmw0X+SD81z0GTUWBNfWjknRvnZZUg3tN1afn2iiymH4+Ach
znZW+1SSn/Q/xAnzcMbCiZ/P/KhclocugM2uqQ09IAYW5QcI/AGAwa4MNJ+xlJxp
WWY1aMOzhc4T8+FAR23I4nRx1qjj4hXzHQRoe/xDa8YT50T/OFrtDnAX5Wr8XX43
0pmgNpZIHx7BXRcmJ1VQQe2fEiqoLqJmizlxCXt44ykHxo88OcKekcuHY6GqDwrR
VJtroM0vPaxUp3xMrVsxX6TVLmik2eSSZspfAWgLEuHjRAtSrgFZU1Acos843UbA
Kgk1Eji+Csm99oDoVDfRttmrtmYCCNoNwwfhNS50/8c+0aCXRIgIxdRJTzs9nl2G
ZfFMg7ztyEXCbxzywZejCuw8cd1GJEPCz70CbCbWY/QpFP1niKgyWuMzIzXJOmFB
HpPFNdOnCDqbW+pDW+KlbNecqYazNxxn5uAziABtD5c5l2stYQgjimTLfTkXJJz9
cDvkEFMVVFgCpaFMlApi0pSh8tuXUkYz0Tsn7SzeEXHW3VqEQ6RLYfNryWRNhoHk
34oDa6VNQbHpelvqgD/FLFiS1J+dqvHSAP/L6bH8shI0tY+3j5j84xWxl+c4YnIb
l4c+twWSM60cA5R6/MCg3UQGxrab25SQ3sF5Qgf2bPdFO9lIuc4+JI4XUPM72L03
0DfmGRBnDjDcRBsAEd/4gLjVtQg7AL5bhLhZuJdM/MGUO/FtkWOGuzNyVnJZTOCu
bEC1ERhMUso9gBNAfxKLaeI6i4X5YgOsRXZSBtqzXJsD+onrGHojdBzZ36u6p5bk
6TlwioyM4JBy1YutrAbp/z+H7aGS1DVyUUO8lsXIcxrp2hAAzJgOfL5s71TXTzah
N69Nlk81UKOeFiUzlaYOb9xhchmmRFcVYDW5uU0e5DC78mrpiUjuQ2KG20rBa6xW
ek5u2285rba2i0qRMinx8sfuMS8F7KcksKOkmkAGBptqJqpTdBX9QYvTevRqyUff
/SMl21eV6hGOQIt+f87uUsvPlFiqK7wiu2HQUUijTvcmEm6hK+fxfEeLJZEi4dz3
AwTfSdkg3l4NsyegJOnq6GzFKPeK5kfGRUuyU6TrQbkIaRN8IR8uGMRgwYR9Jbvg
2bWfZF4Yf/OJEloe+N9rXDEZsnzgBLA/S7ICWjqQDacVI9iaBwbS2J5YxkY3SrNB
YnBbZp2NIRTEubkhRwQywY/s3ZDI7azVq2NWcoGbLwCmLDJqhosIvfY6xV5HimeZ
/9+JtstKo64yOSF+ycYcAEC9yNDkcTu8++O9rSZo2IcWXWzxisBSK8Zaws0kw5Ir
VxTIDf3YikmIFhclZlD3bxxMcy9kIm9oI6vhxEWLcWx0QFdemRd2SjrzRm/+0Qia
al4fYsIGOPGqZyVuIGQiPn0mc4KLT5uD+QgeH3DinplwsDuiRIox58W3On0Qa2e+
cQf5I9fkqb7FI4nai9tbFbi/x7B2d5XTH5VMQMoTdq1efrYU21tJB33vwsJU0lik
H3v3vvYkZQxjqlicuPF+VbAI1Sv5Haw6fj1CknkJQU3pNA2PaJpdQrDzWknchkQ4
A+9J68MD/iNKhf3SDdPZTZcIzmy9xsw1CiQ9/Fd97G5trb8oTnDv4l/WqnSkHxLx
3rsYThrHRDEkXz7Fpv8ZZr66t9+cPXrSNNpGmTHDbrr8HuQHTGUzBTJ63zjajQsL
iR88q9d6QbD8dL/J+ihUoLOZ2TC/fYV5l/jef+iMQpPGnhMZfQAmu+ZB4Dj+6Xk9
6J8eUibPSqbgbEHlQiNq9NMqzV4OxQMszOno72jOzbo+NWYLPTZCFItjDIXmIjsY
MYIz+GPXyMi/zSio6NMPkH9m+gXikYjEFzfPLhfsgsOFtk/YxyuUi1eknnenObm0
ffAJ2FX3AuUVGx5dy6ax+OszQtzKRT6zV7UZ5ppWTBqZc4qkTTGuxBpim6OM+YAB
7iLpVs+BWsOGn+lqOAaXiqLbw4s6QYpHRsdSXU5MfR2oiuBc0iqEQM4R1FXawpUg
nyghI38/KSbHWIZePSRykJSIDrULkgOrmFLHPCxiUVb5oiketKR5kr82lizlqiXF
pQ1csN5Uf/9VSK+JE0JTRceSTgZOlTLBQd8oph19oaz0zl2sOg+tau+dtklftDg6
pEdcy08w7hiN9sgaKzut+pEKEz3u7orrC8PHqWf3iqGRhSocuSgWuiy2rAR0fohC
NHhtahdw2EIe9P1fsWnFNIfBeE6K2HjoCWfi+jp4+e+r7iyGvQgOlJqG9WNXIyDo
Crx7m/umCBEwpeD+AzBRWmhX9Yp1NmTYNyoNYLCWl3GEEB0jXioKuKmazuuNIbkC
YpE+jHOk/JaEUlAnKs2QAX6dzhO8vyZQP6Jp5NKGJsEBEi/csPlIOf389PbWLiCh
Jg5tGp67OsJH9yqELUKvoPXgAd9ubNWPxUhOWZBbW75MgRtsKwuaeSPrDjQMeSy5
CpbKQPVKMXVLdhyAR4TGI85k4gM9R54uoKshjegGaMFhu7PsWc9UHi+L/VUud2LE
in2OXLR92ykTfzCKKF2f11sSo20Ca8d6/Qsu0cvNnrQ/t4Z3PHSMiQrDvM7n8T5R
YC7STH0JpueZ5pnVlUXw0w3/UO48puiP94PVO96V7txddp5hvw95oPbv9SUxbBVE
KVA04dlVumMTlovF5I2YozImEbr3QkpL69Bi+0jwikwkWj8X6pKRODfF9k8Xhj6u
pYj6z+qNghsDeBAQIx1DKpdIBmIs5PV8SWhEPBieCqQjl621mxir3aQa8RyT8t6F
HS3d1WDLi7KYUitzEsz1xa+jTtarOGMauA757ISfmxG+bp18AR7URn3ziu8GUOFQ
b8JrQAXWExFOfQYmi4iCDgxSYsuBWb939kaerfu8pznKZP5v1MASVtnUujUB0w5U
/UrnvRbgtonv4gLrgDvStWiiSYJZxTp3nJI4R/dUcOrq2BUqkTBW7r5xTWRTrcwj
lESAJ54hONmZY6ABwTR1a1zdcvU9wbuzzTkc7pkKadvv3T4KJgcLL5f12TIOBL/T
tJ9naj8xJ0XHPL5XpyNEOYECbQ5s7jbdSQHWfd2XszgGVfstj19D1e8FX7SiV0rf
Ap4/wlKG7WSWavimV/C0mIznsE9+EVP70asVP+jdZ6NoAiXHt7eVVuN1NvX5Nuav
MAQ9BemL8rKPEIdqoKttFdUPXgkybKnCBGIg21XTXpj8JhDCP0WqeN0ez2FUth0h
1GR2OegUn0/g5dH66hgEgaSlubWRteHejPXloQixrR9WRB2g6LRFAw7PZWJI992c
P87irKl/8ey4dKC6PfgVYtzuUIzxADcyg43BcZgHYKv+3qh5DCxEU+WG8qegEYoo
G0WQPxgUwOltp1jiO0O2LXTL+Szs2/w3pYvZg1LROE/xU0DaHqR/L7w6ikoMxMDv
TJ79G0bCMelxq8HjrNyPGf1X70YNQzUirqp25AqPsbvBL/U+95YC9exU22bwSvQ6
/sldH/lJWVZr1GUyn1zNtLXgorerElkGaMNCiCeuLCpBJozjS7EmMBJuRuO2TPjS
BdaJ1fHU3KaviNMsjRlAzo0FFD9IHOuZtgFdq0tB+oplFTEroU3/jt42Y/o3rcAB
PxrAZdCI+gKMcZCR+gJAkjUuBkbpa7Hj81JxAh15ugOqDSD37VV9ZdQYWCCkIr2/
8jqfI9KTCiAWNp5CInuiO/LZ24KS3bc1E4fwDC29SqCr3xpeiFYV2DqPxwOSwAni
5yedI0yXJV+lxkO6R2gK5wvgSQX0YlJovf/L0ytN21zrXbN54DkyP2Usx9SntjXu
6fI3aE/1gjXtJ2pzhd0KZcATmyGlj/6/KG0T63w8/m7OHDBBGURLWfHmQT1decsd
6rw6XDC9NuC8rjxEv4CNEKH0fT4PqfZMeEy6UmCZvaWY1+Pip+ETBzZST3D38u/4
gOithHX8eJo5vspe7OC3h562hmS7BexdhbLXqztakkN0QJm1celeT6G9iPIfSAO7
jN1ENQBsG5qHOWL67mglQlHu9TPX10n0OTjMPc2GO6y3Bj05W1wCbealsPAnt+9V
uSOLMbOMCrqZyXqwXg0bllXCrE6oxJTkiliVThmUgvv5r4tvILtzXhongLlzkyuC
lELNGA2LHZjEkLpkIPloiJfpdsYwaiQrslTeZT6vAU/v/4TDi67qsPmJJvuNhX86
ZH5nqjCUuSrvwmc756YcLjEoRLGyOrLlVmqS4AYS5anojGHvFBMky0sx4GrpZEK2
ChQGIawUE61Xw9flgNgpzJT5XijdjkMNYLiwEL7+AydDE1qKVxGLX/I6C/2lGars
ZQD4kUvf4kAY2X4UMRpdcZJR7pHMcQC4Phig/QeTMg0Eh3OH2jPW/UM14CcE2KFH
5cz7LIVr249JSCRCWeOGjh496QvTHO2KdhVj64H/VX27NDHv48TMMO+VriQiRf6X
DCowNSpMWeHB/h/2GXdtM+K6Wy/GgMkFJOoJWn/jaqciG1YxRIRrDsh2klrFNcvx
1ggO1Vav9WJXnh8JAMsmuYtujrHVHPtS18Pfe/aX5d7/NQgdfj+4KNJd0tP/8EUv
lZwxzv822TqLz6EB4mGl7Zk1Dt496Nmcn6UiKhAazuEAUtTLZSPmxw1G4IJb8/eR
fu3ep2aruN2N5iDl2Nn9naD+6ckUBs+e2yBP88/x9N7+J8HcFPbeBXTCChZXlr1G
ln6I7w6qhk1y/iDzWaAjpX27uINaktnwCLAAL5ZqZRCDertIxZx3JRXBjDLrPHYE
KpNHdifhnppwTbDaGTF7uBb0++1royRtykJRg7TeudtCMspaYyKatNVvPL0JKg8L
RXwoSW7EmsaoWTK8wC8lN//0GZ2K1mZqz3CWK+WUSb1QFCCT1SHUNaPQ99uYjgaM
pe4AChzhkfOkXENGn4oNBoEPaRr5B0KriP4anEjScZfMsWGB1BD8SaL1BLpehI1c
KqhYwhghVC4D7CceMtH1/0zQB9vVA33NCToTbAkS5gZcDGP+wN1shldh4k2lewXk
kDRnk7nO07k0It31b+J4fO+4fb0qcTTYGsYV6nHXk5oYT42NBEI2/CtG2UmSrkss
aLdedS3M9cS6bCMH6lHmR6bFDcoXJiHuSU5EgnwrV/6yxwckpNWo7I3OqabkDPeM
UicLfojAOhH4q1ZbdOcMe0nuGpRX0dLgcl4fxEQSjrC2CqNSI7PlLF1QmkkW+fYM
AIS5+SjSCqt3r1Wwfq4kZv9s5Ha+aCN3LR9tuVOxv9VVDOhSz9PdQKhy6WDOTM3Y
ye0gjGU2th47yRhoTHi8T7KmjQZC0vrP5pkEYACPmMHmucVquvyrdD+AcZpvQiu5
KzJQa1AUa1zT5zRJHIC8h0o0zL/HaVnUZk2k8kU5W6+lCsjHJNdfNg+DBVQsy21a
Gb91UhWSnBCIOl+E1YflWO3DNmTi4xHA1ZjGd/RIdFpD5WtfIAnNH4YYh6TpB5SG
angCgLVDvmzMFGmqP9FxjpoIsHhK6zwcMmoZzA2td5rvVHuCVe9hox4AgV2uDgMd
hdS3HYXIQEKkrO+B0H2gwDk2ZcrwvXmVx1JMyag6IfNxg2W4VCNgNKXw4hyx7R0g
jSsNo9rc2nZfroiKeFCBp7GEFbPC4bKWwB21GgBx46lmTe8auOdJxWmMiMlm68zu
vJv7/DYbBKT+hlR0Tr76DW0RTm0uIZbMbeGEC/IfXj3g09clA62BCTmk4OmjK1kL
kB6pFrYr+LtI7tba4vZPkgMnNbyti33YB7DC9aZBRT0csoN+F87ern6s/IQ7psvK
JTtsLw6wAIUwYwF0hrwwVoRwoB1TXBoEHh/gPd201FrNw0dVcBkVDqNTMWCz8jWj
4Nd347fRJZIUekTEEgbG13vxLXsHcVN5PffS/RbHOwoWM+K2b6gl4a7m1afAwkhV
GQbmAdev+Bt8TarxLbQ0T/t7xCpQK9Ktilp2F94Jz0Fu9+s1DLcFKCbzJI9R0lxM
pBHRZNmzkhxu+ZqF4HuFB7F4r03sNs94zXf6bx9NCUUvqucoDz8oQ1forXEaX1vG
Bt6ziqNRlmYobqpiNI3TNvFXYgfqP08hK4C2Hm8q6J1SrHlVJeEsh15e7aLkm+O2
5g8lYBDOx1BBpGXWafu44DhwKM2dFDb3Py0RVxGR+mNAEDjMtBDEy5IgW6NRNmBH
nTX2Kzjk7ibLsJsOgQhRXoVAOuvoOAhBOmACRHdR1mQ1r38SdxXhAc8ORC7AYw9b
26eX/dOLHkeAoqQMZrKdLl1n6iKMKRd57iSA8ecYVKqoBd6u4I94LZxFSik4u8k9
xGYvqfvO7u92qk0Kd4OeyyUZl0zT0LwcC2jPCJPTeymmQMqMRP6sUQzZ3ikn5ixB
dkSITtlWXNaZjuQU3xzGpfsmfPmhbIx/AmpxHSIoU7CwBw+pwg7h8CqMS36Wl4oO
Vlwm08n24fUs20sau22Ob4VNBKrUncDAJsxWAw7Ksf8uKnIamAO0QNQKrcn7bfSn
51u4JmIoHPWkyeoh8bhYhh3dCD9QgYNXfh7dTrhGISXaliy3svYdKbL/YG0k8xWe
5SBgzEBSGpFUrXbHCHAOmpa/tqDD4Shb6+YZeYczZQXsRaJmkBIeopt4fGqA+m5c
K2kfUHA7PdeMVz8tFbr2pbaDazdyUMbkehsTKqJJxGLk2psZ2YVywr2VNCYeyB0f
A167Sij7fDR+phUGvf63pnq6/hVAZV9b9nhvZhTOhk62jeYCNW6ZXcO/grrWAlzx
M34eDTw6MD4OdkSQZ0yLFXDYtdNOtPHRQK2riBN4SkRnj+HkVtZLF4lWk5YOSjKJ
zaRYW0OO0XvJuZPWSCXZ93N8hgavbaCnLszqeXiXdG5LDxv0ZtKWpgiOcYhmHACu
TWN65E8d07OR27mZo8Y1gBJkmdK3sqge4NSPjpALu3shRqBtYj6HmuhNYaL/EG4e
cB12HgUImhgWflf/AQCaDLtRxYHzUCdaXJ14vky4V+hGenDJVhdkgD+i2QDhr+sx
OyU5TE0v7YgudA/HXTnW8fzgoQP1btGq022y3Irn0zqVosOFZAx8gyT23n173g2p
aQu1E6OqFtL4wYT05TdlWVAc5zgHI1ZtSmgvWDUtxBCYrfkBgsH7zajyk9FcVFOn
W23Vc0I99KddiMh6Pgt5ZdICveqEty1nHvc919B7mZfpUzXbli9bfpdk3yQgVh8D
2/u6O+lHYOgtIyugWUgJj3mEW7DVPjYLXoj02pC8bzc6tF4Pz0WzkDqoTuN0QnVs
4gKR5TkHw25YGpJU28ZoZO4iO7qhzja4Fv/2bu7PPyZRmp+HExPOaXCX++XqodX/
mfqm1CTbhLz5lmyPxPtFv3tDmiobwPsfGMvydNUamXQS9ZtsTPrAVuY6lDWQd0hi
l95p7/2GylezPTAQQQWwaTLi+OEthhyv36pik7U2QxRAoXjIvtC02MSXs5e3uo05
lL05P7YjU9gjJaZeciE6U33W7s8Vm/Q3dRl9vqdUNKdg5zmtLL6HhzfFbud9CJJB
MJeaMJkUppNUurM03xzeFd4WWJM1fugV43XRwCZL3YdDVnQpu9cXQ5Hs74wGygWn
kqw3msKYTVkdVst2PmFJrGvo3RgCvSm5UL430cqovtvcYZ4GslaDOPhDLvhM15aE
s/nRYbRaMGU9MmUOkjOGBpl7XeWwAEVBcNFi8ziGA/VpS+w/bL29IuGhh2R/7XF8
rxfhVEbdPNRmnw+hY/eRLBI0O5PLbEZ+WmDa4fNYnu+CI4FvuJk2M8l+DnUGYzqB
S6RVEFtG8QsZaSp5PEFYk/VSVBAI4CtZGUmOlGYKo6tfLKBJ2gm6O4sOM3wHC8Pd
4lEbyhUAZ00KmGfCrVFH0zvcfyVzoUi2S8e033oEc17RX+HaVobNm3vuRoGhiAjD
KyAz1HLL4nCRJpF+aDCcs4xUoEZLtwe/wseLkFNPEKmmDn2Wqm2kUW060wTeUYUc
PKxK/YMxoXN5T1I8cHggRa51FJb0A+rdMXeaDEP+xjvbQEmGTuo6m2Isa4ja3y1p
CQhsBdhkxESweb41lyctoFLtNJS5U/47LfWNxXPs3VkjYCswF5emfGbdJhHgFnjE
uEco1cnqH1Jxtdlj18Q8P4HWj1kEa3y26S4JFvaQhI/nhTBX5P62LRa+vBfTsFOE
GwZLKuKpFFQbAr+1Tcu8wZtLpk7Zydkmg++C+9IV1hsUesW5ArNCb9+/+jstX9qV
gJX5qVFjAZV0eG1KOTtvKT17aqTmDWn3An4h92Tyg5EfQ7dti7a+waxRLStf8EuP
5kfjR+Jbcxs8p2CkYl87Y6Y3kW1uwEsn3ZahUCbfRczoxbzRawWFMFtIiWu/dAKb
KsSppWzWv1kAhnze4S+58HYQUoVwh4VCC0JVWruP+rIG3vw54F0CP/kmpB7ZLlAi
blNmdVkzHMRJE8FxaYFHvOz6XjKNZtdHprpvaYBkmcUzu9t5TI6NXPoGPamHvq5N
HUkExqjEwctccWk2L1vcpgtof+2GYzbKjBm5pQV6R/zk2McQsfbNvhQwTLLWoM9f
SEBCD4slhF6vM1hFFNd6xb/ykatVdQnOv+y6Q2pShFY12aUGk7Ezv85uzx7OkCQW
cdawSdUOOreKw2gR6IrOpdSw44+DqauhVfppmPewm8mWJSkiLtIGbMUEPodpg9y+
1bW/t7rU3i1uxv9trZpNhnZN0Hyq4E53I/UnIenNPePzJFS6sYJfO4sPw/uyJm5h
eDrhk9BjsOHvogoctkgU0SOtM+ZxG//59gxY/2JQQZPyZAeM8yb6qIpn3bp/29jd
hcVrd3SFxDgtwQ+XmRadG1xBlvmfRk1lb7vf+VJXDtEZmCB4mWGMhshmDDmG+LhK
irY+itZXIGQnyVrK5Ulyj5XEa84FWzSc1TRbM8ZZPMV4c4Gb32H9+h/YbT/453B2
6cgeT3i8Oc25qxOCiJPJYj2JvAd5L+o1M18MSlqGD4qD8uLEqBJ0+wJP9ZbJFHnN
e3sZaz/OiFk/ejMmjbzOQc0eiiYWDnjRcHMPdB3rJH+Hvy6m/W5xejn5tQytGEb8
51F8O0MqDgcKoOB0/P+es8zJprv8PO3K/wXTIJMaigJydvn3xsSGZVSyrE+lJqR4
5FpbPsk5CINYbLOyu9V8GkQONfIQx6OqTAqQ3IuhDJYPp71ja6PDSxbUJEDjc9Rb
1SAABEaRyvn/bqgLP0driF0luk1k6SrH1LVD8sNk5Xe+1aF17QaqjkaaiQGX3pZU
el4Yrh9qng6uit0umCVuZlmw8egMIvB1aArz/E/7CKOne/gDf6Pf3MYSwFYsKPa/
4D9575AHEdIWr+AkHJn3PCfNN081dV6rmqt1ha2Kw8M1aZWADxvbQujuiK34BfRr
rkb3zTXvUtOe2wZyEOb4ftErQla/0wtDSAdTdpooxiqazrAF2aunnMTnb5OOCP4Y
WTOc8T7cPVjmroldWbQAlNbTdTDXVp0dXWL1/S7kfyXraloOU0nhwrcECKM/hFMp
H0PM/GdplBZW9PJ3wgXA293mvX7byyknmTfcjHepSbwrKQ0DDQ0L14OOuhByrOCU
pKIubcW0Vzgs4eitRHffsjuS5NFTuEvWxcvL3YP+MlTOwTkGzURjloSgGDUyzNUi
pIreAWhwlZxtDBaEntMbq9dF/f80V3im41IqVpKJxsZRsVmPN7CCnH+KZGjog0C5
q2QwMe34Vyl7NcpBZduOYyEIvhqCTgVANvOyPL1j+ZQSYbDu1EAPR0mUUtvUMWY5
6px37RC0Vw13+ceirYKM8oNDvE/PwZvOB+JEOmfO1a6ZKwiySbnlHTBBezSL1q1u
77XQTE3GW12FOp6y9/8va0HThOSVl3CegNZip26yBAV8LB4uyQcWZXms//Q8x0fD
TGuGVPiJYKypYgCRIKW2QUx3/0qXzuUxLbnT+mghZy/LgX/DiY+7GbKEuV6S6K9R
DZvOLHJk2WL2aEb8cBCVV/2onji8EGmB1r6Y+alA+dsT7dFJpYjCuYK4Pqyw5Y+e
9gsyiIgo2HdSwmiuLUK/YNXyUqVI/lqsZmAagP9mshY+UqIDIwmO8LcADJIOXaxo
Hs9akRiu5Qled13BsXNHSwLpe/Sfn190jQjel4joDIvWfXmgAx+9OugV4AFK/cz2
ljsA/46el/72EEcQKgchQMg5Oz0xe47G4X0h8xLdvCKwBpfM4ntLAsuIsXvsQdti
8lkVmy59vlojbCQn7xKUQukbY7K6Fj6NTTT9afH/zTAAmFUKIZTJ0yTxXUyFR9ha
GK+nRrK3ZRMUaHQbMfvkUUGfKIvuSne2mvqld9bh9DHp3DRWWzyvmvEdA3Uh8Tet
oT4c4aDkETmj00aDEq7LuuX9YwIQXhymBpNoPJXtl5LbaplawC2ucdYctBruSBdI
2VJkiV+W0WCxcBBecJQ6tav58CaDtyodNb0lQSaS3ZbGc4ME8L8O14pJzE0hshgN
kMMoY1lvxsODsE1Fkwv/NX2vTxY+7F8uS7ho/sftSRiLvqhGDqyecVwsbybFQqIC
DiJaIdP/x72ha70e/32E8RriIQ0K8XCSfAIdyBAegaOGGcNx0BJJY1Y0gt4CkW2x
led4zjoUIvBckSbaBWnoD55OrxSYJn64qFkC7mCggn9E11Nglkk8+XihuyNZk54L
PqVJ3rFeJIdmgZ0IwIJYnzgi1IICs09mTxmzrU20Le4Az3KAXpNXDGLon+crNWPM
ht4YT8l+fRfwUDbTmJ6KJJQQzg0yvMT25pnp40OJqiWQhXJbUYi1buArxUaj25Ed
22bOXB+AGub7ZJgVHv5Lhdj7xf2Oz3qn1ZRbUnHCcs1XHmpBk1cusjHV/bBsxaS5
hJLflXAzVChjHXC0JEtIs2Rdm//gE97vI2WoUjUIMy3OZBD7YKO220r1nCasESI+
Canv4v3q4rBfS1gA9KqwF2vF2GgCyp0wnXtG4etVkaAiVd1esnRaEPPOokG8MfNh
yejS+x3RqPJMaklccj12kfvbNODlBRvRTkhAsT391MuMyV7LdcNK1kHiDrIR7j4Q
YeLuboLkYx/p1YJFYAPRfsu4dv7udDAiHb3HLYTyi6foj134sw6Buoj80MawGLeN
DV7U4rKDiaXXRIK/+BMIQiinXHrFacVHbV7UZJ9MWYoB0u6Ro3OoGQ3jMGNbqO8E
i9jNK3sZM9ptooaKNE5cKAazIyPte8poCshlmxHvTZ2qas2UPP/wvy1lvtr99bYc
fUy4hbLhWSLiVZidjIbrfXUs/gww6fet4cD9AL6DJ+XE2ltyOLPJfrYM4Z0zPijh
h8d/fB+BqziBqffPBIzLIkk2eL2h/HVTn2gSSDC7/24qRC6X5+qWUQ11yWQ6iwTo
qW5LXmCMtcG+FDXX/PRXApvQZvqKcCjZHVErbXpf/Uoms51+HbfeySY8NKGI0r60
CTXBEYfUBHswsayWJsk2Xb/J/E22v9XM4PvRBURRtdvZl+o7J3O84vgmvJ4LaaMx
/aUizT7qkvpjb1WkCEX+wVi9fdPoNv236aGttlzwfLzAIYfgRgB6QjE+ISouirX+
iP1+0EZbH9dR3WRKHMO3aDVHK0KCyG3LhhhSFu9akrLesaotm+mMCQfolT6ywUh0
adE2cBJ9xLGgVxftBO5C0VTvcIF15u4Fx/RNDRrgQxDzHR0N+xu3sosmwDHZqzTa
JEChWdtdZdg1mRoVVufEPbz8P+NaZWPmhAFVzJ0aQZQaQ3PyicK1esE/uOLcfhWF
hwUD88cFbTMm3PVRifKvts9D20X2O+ZzYTTUT6+7rTvgkifTZy0s5W8OXcdk3jaA
VB8y+klhH5EfGpkqgeEErP0wYuIsa9/tbEPADePS9XaJuEnt/yCZ2zty23KmtLrC
vFFjnHITlRjv+3Us2y1aN2CSLU5Pt/YQyVtS4oxE3qrhHgqaCnvttwANAho6bBI0
WWw/tH5/KZvwOisStUx76CbiJUtRfli3BfIWqEIdlmRJ2sk4rgk4w4wZxtvnAWbI
ABN6TtqFRwlZPkeqNzmyMVvArSvDnudr6CGcRFlnaz6JHX2YH7MxtB6mP3bbDn6n
8lTPdTLNqwcHWZv6ICZ3PBUTRwrNLoV/+4FQUQ7A8Vg4fpejI0/WINJ327azqyJE
vtMake2JDcZQCHmPHNmlJf1Ryg5X+WxSs4Df9vCowG62GrmdH57DP3f3KRQnurwz
hQdgUcRAKiaE5EROUQDOHMGlU8DApEXUSYECniF2txHqo7TBxb/TEq5xImv08okv
V6duN+4PNGiPCW5AItnsQ2L2QNXrWXbRIbhqgjAIGyMOkiGUi21d9iHXFeucMmSM
C2PaaDTuDxff3xrIASogZ10x5wFab0wNHN64jKegGLsqTjzoHcxjaFWpLx7wV5Oy
cfyl8tazcbcfBw5MrWXXwy8vHkEvo+8V+NU8ZyQY34rR6JXq3WF83cwiSu5iIQCD
C/LQT+6s3TX9h+/yIrYWPZjU9r4yZj2dZYDgw1vrxEbpN7Un0t/zkDJuWFVkBsu/
g868f9s4qg3oUsoATXl+BT8vPo5n+lPWBa60/+vFlUHiCLWwiybkN1aLkPKK2t9t
FLXVXLr4+KrEZUipB+o75LaCsu1qhXo2JDPJ+5RRJA5iP9Ybas6HTui/xmZKc3oc
M27Tnjc/iuDqoOV4LX+qbLGJ5bksyYCXy+bWU8460FysHbCqiTpbaguCrGP6QI9e
W9ZWKyQamZcLv32RH7WdCBH7SqBRhWY/AOx8HsWUv45g+kXKSAV23uJH5ESz7oA5
xs7YI/Ja3RVQvbAY7yVqEMN3wa3Pl6V23+cKd75NN0XzOjLF6DiEgd3KmF+jS78i
gxkQ/Yj94aN4GfwF25oIgqxAeEv6eWSttXBMKGx26bCVJsKWklFCZW3+Bw+Ibq81
6FsPoAOkQIAIjl6Q9wt6B199YFD1lrui45SNzjrLIEfb5PXMKxZw/9Oxv6x+N+P7
19+/dzdN1tBlEb8/SU7kGouC7V5OF8/6aBis18sCYHs4/N8NGpdNmp3bVGN3usGl
yOeLo29I29YeTRHT7UNdqY5tAy/WpVYWIJNZdPAdYJd9Icdh2OR7sstTJ6i1XGpv
dN9p8GvZtP5Znt3yuBmLrHAsiCFYzUqL1sZ2qJyEVD5j9T42hky7Q8htc24hHg6K
vp0JfPukCMOlX41YfiDOkaNARONojz1v5eG6fBz8E4R5jETVUXUMFeDhTHsVVoDP
zXkaeIyDAgIJAjniGoG8nHAIpfx9FLDMsU9cTMaNp9l14c3CM7QOsq3a4nMn9Y7r
m9qJUDSbSZr+7/2dGVRUmEPb+ecW3eqq6nxg7jtPgyxAI/84kEhbw4nittBovmC1
17Te756L7aydTJRUrx/8LplMvLPPDYgt8c4w5IHYCGmhEV4jlvWqVQraPQ+ZTJkd
ATLL76uXW1NRVAPay6fRS7M70Ae2oOgZO1Nh0IIlJuVFCxg6bS98YEuEzfSB817g
y/XdqytQR0aWG1qF+VqM5/Kdi0FOy1JCrzN3MEJ4GlYPkuJOm7TxJE/i7wgdiVNx
a8x/4bSAyTX2ARCr4WU9gEziSif5kmJV5+wzDFhkfctBVMSF79rSniLqFft33ule
g5z7dupqELlhAZ35V/HdABsdyx0GlY//zBHHD/0gHpceTdEFJtcI4klSIlkNfTzp
ilzPJ1k+XORz+/kOFU59U+nSslRmC+UOOlj2R61KATmM3gZ0z466WkdpTQSZVWc3
zYjI6Z0KdlfYdxWl1cy+lhnuL8mjRzmyoF4dmBX7zG0pMljPkXts6qDCN185oXJz
EranNEHQlT5pwBr+241ijb+JTeKXLOfGQDfRvyM6fgs8NdZVzjB0uiG37/rWaZLl
wNV0c99cLLe3CdVGsRhriC0VBOuqOHRl9S1DfVCQHBVukY1NDV8cN6glzdHg6zu1
ZSIWcpFghFHWKZxn/y04YN9lugzuw3eEneQ9aqm5mDOW2GrmnLEvLwcpmKDa0+S8
BdW15KV3U6okLvZk7DfzOGvglISMsiVGWa1lIjG2O9VkAG6ssR3XTbs131wIAqiQ
mse8TOKQKTQCOG+VAyk/ZzxCRF6NjVwkcn7zHOpqdMgULamrYCVH/AVv7rtEcuuW
CMWTyyBlY9UaN2uhL86U0oMghcn1Nf2dYv4D/BTfLhndBi9Yqtzb0G7VYVairVHC
WwMqDb7Z9AXpqx2GnrFwzYhg4qtOWH7S/FnBsf0NHhX5PhwZhk7Woy4K5bYCO9Cc
KfXCJjxlLlm8+flhrllXwfzqlMOm7Nw4807qqzLz8DUki9hAkrjZBNbxUFW7PRHZ
cagoHgh7Rs5BGdgsKbxYe6UC+0v5S4g4xTRHrxAkiayuGwyradK6fSBXgFh2nztX
Up5B3B2Cf+GbFdpWY6WiB0l25tEwvCn2DtIaQrMTLmiTldG9DehRwgZbtFz7hzSC
ZKIaCzWvCi3NfjSYqITyQeROeo5oveo8e59l5IyTVHaQMJdmFZqmvuV2BJU6fAB+
e0xHtkuZTeK3LdBR5vCuGFIko8jeBtXpyNt71TeTSzOsBfwtaMi/iw6f+ssIDPnP
mV6NUR/XgIU/840+FQo+NFZ8mBxtWTPIIU0LwwnEcyozaiv3iVeFhAvaaKXCmRqp
xPc0Tw8xZ3oqtAezkDJqEEzLku3//AafXVR8LjEgTDCsQ2BWAjDAIZKoU+0lxjIr
AEbqExPN8ttYN+ruTKhTKMtS2LH1f/8yoFJPgcZ8Gu0vAf0uDVkfqB0ImTObw6jn
rnGE2SQLp/5hRv0e1xqqLMh0uR1hSAnh5ZmrJwGGL1qK292kNEJNgZiLAOcoaFZ5
MVG4dxJqEE2IyEErQo/NhFuwFwcYAweEzYStFjbzYSeQdzhDjLUZam47zE5dnTEl
Qa6ymHYs7Fs1KOSwTtrDDj3WvXNX7t0Oz6/xPY7m5SqVjAtttoFTmd6xyaMGTpFx
9TLI0kJXxjL0/NUMmenbAlhdDOycu2vrKq9OxApEAfWACkeKg+sxtUPmF2c9rszG
fOjl5qqoAN2UzQ6ZDjxlA8ISFvrO5vjGHcY/y61IYgyhTw5sI8YyQgylWWTmCHPq
NP/bRL55JTV6LrJaXNMMofTiU888qwoMSighrrEjp2xk/pjfDte5hbCUy4doFkKx
rjOPgmY4KJe1a2Og45Nm4RTKtllMmWSEo8AdR1DIa8S56QjkeTX6gvfweHpdCXpG
fi+pR/Etkd1miMuYUr55bIOgN1oKo7fsDWBV3qiHP1gj7vIliVfBQC6RcFwEL5TC
PjfDJt/odNw5tlRWOJGp++iZkiixFXQ5A2HBMbID4klL0h46AmxoL68CcFR0FL9D
mx0RYxBNpMJg3eH/zgYbrSC4pEBGwklZvKOXnW8Lpo4sB+TlanrVxB1KpzrqGkoq
sKnBwS20RepY3mlC+AEuvnOVZMaARiLq1dCLXsI1Q8rHoTcsQlde2bTTaSZlLLtF
eVst9mOULP2Fh/UhwN+6U6i1R4LVMKvufXz8BV1IrkxY40ZszGLdGXujY5aalVS9
lIYbmcJmLzvvH+Xnl4vbEmvQNDW1ctU9e+r4eI52dJBfll01Siw8TD9eHsh7d83a
IYF1GD1qQ8iQz6v0L8UMnkM25wMImMSRloyEcHQxJ6t3ZbOcZvevYQRhtNWOp/r8
Va9x7paA6I4zjPVDD8L1Ql4hGkil/xJmoW7hAquOwbxi/7kFNxqG0OmDiqJ+cHS5
d6lAJYZ+D4b2g/11s+AYZb4DhBAjOjRnmWU8OZx2Sky6s1VliX0s2Ybvf/+N2i39
HX4R2wRn2LqfVpcPxUR8E+Ov1cyzTpLwhtviwDVxSSHZWsG5vYZF3SBbg/vSskWB
Lc1UaUEqx+WelNSBu5D3UG23fLQAhvSI4VkHeWwz0jWmCeWEVvrWVqd890meR93F
YWXy2zZvL0CE4jmnsfXi4GO9cbI+hu1g+yMqCYcIxVBSN8qUzMmxeXhjfG1CvrLg
mtPNF89JdYIMqW+F2iv3ujmXrLAAbn+CkUb2RgkuW/Nzb5/bY0OaAovY90Yu4eig
9QNOGVHDwlyElMqE6lHBM4DZl0SjrmUoZn1kOF8jp8AmODVl+1nQVADL2C2GgOh0
P6mq9VL0N+g2en+wHSDoSrxpPlTNU3ZOAwlUiSU3ZdMhktjkVPLsBIRB/j6aZTtZ
mljTmIJPCzR1dQ03n10ISL0GsIZsyNSPHZSESnqntdMTVSXRfMRrm3gORoF486Op
Ldhd/KW3ozH65FfkqlPbZoTQlKGdSPmm/5r8WV5+efKZzlMRGzsKELkBgwJeBFL/
LmzzSSyxE/e7k+jdin3/pzCmKKP4r7AyLsT2iIiuKrgv+u1OSy1Rz9oCDU//0IMj
1/YSzYOqumNw8TiTB+nF7b5HGtPXQ7ytfdEptyiYx8vWZAZJhmjp+goMvD3oQHTg
U4mmqjwmbTtAxRq/L0I6aorInHtbtPmGjGMS54+CL8vHSoG60C6UWu+XtGq5U/WN
Fw0cf732SYQO2h+Xu0+mU/dknZrnJxsmT+dyZufERxUgv9N4nvIBCbY+a3YHvEVq
EVcP2cTVrWIGopcU/51v5goXl9JAg+ENjhdm4yPt4pCFUTicEVZTCh0lXzxuIX+Z
Yz0yxfzfZYPKyMilkhSChIbfw3l8o1Vb9KPx7WmviXgf+chyvyPWXDGyCF1hAYqx
wnRcDSmbQq/Y7xQ9OWQbq+dCyIZsJfxNmh2toncoNMsvMrY1Xb8jnJ+FxpwAI5hY
0AmF+YzO6/GHcaP9JsNAfaw9ATJhuNfGVO11k3XU4yjzpIihQfx9mhIYWAOfNfUN
l37qSuhfefLAXzSQDbCD/uxG+wF8I/FpBb3LP5hXF7faUDyC7Aghqgyx5GYOrLsw
Kz3hv/McKD1LwwzKHcA8TSGJ28jo8bmzXzIxNLbwrTGYi4EQODX4VEveAd3wWWgb
rO32KXEkXJ9quyOBZaeWGEEcHeFGHTojBxqAvfb0VaIem4aAITKKNPM/tx/U3spG
oZotQSKTS0MQ5M7dHY9an4TMX9cIMl7WVHpizQfIqySn21CXbWiif5NuiaPYLIpV
wlXyp430d1IwwWg/mrSUXjqvZg+2eedznfN38cixrptkrDTHJL/xAP5Z7l4BhIWK
hCztUuqucXOuQYPnix0gESXkeQsmvP5lpTYhTivPoQbc6BN69GEVtJf+2tShUsw4
ZOd3lL+Ci8lBekQ0tqY3TOMgnkYX2WT4ateBuj94FmGUrnAh6oBHPYwkvDGvPzrw
Yaiav67M5Rtbvy2+T1I3aBk1HK6p+EVghOzq+tzxzzBDaqLxRRPcZAM/CBKY0lBE
D+nWpCsZ5bqLcF3+hPaeBSYO6TRFqIUq1+WH89glQhwMPjqxsl4nr27WTjfVALhv
AgqMqcPnV/VUh+eX3i0pENIgjUygxBjXdUoUAqjVSZOScuO7ZiCgeKs7EZb2NRvp
vxbyMMujOfXWJA792Ka/y1xK7B2UFBNCXvIlCMY+cuy5z9g6r62TXyuhx0xQHm4i
CdCgcqLUjn82LRF6eKgGcqzoJ9jPJKPqMaOEVAWuUGtE5HoGd2nfxIjFKL4Md3v5
WZj+WtGoQwvufZQqE9z6VOEpTvU1QrY7/g6PQPSuc5zWrmzc2PapP/5X707Rch6p
T3QBM8ntb6wl1uf97hzTuC2dqcgSSYu6Qr9NtqKCsjsiplN476FsEFEEKgsFv/xu
WH6rPkrZ3hmDwsRrAAZtZfjbkzvnnL+LueiS+qwEX59fROEvzk0ACaSOUmWctyFL
9okoaLLaFvEsGKx4m1gsnkH932Cz8+xxBm1NuSVofLCI5HBliGbtW88fsnMiiG5W
uLmcoZCBPX3HegQkeBVwF2sLX8IuELpiStVI+L/iZt/MDOxQCOSAmpd9c+DOxvIo
AVoQkdqYF/SqJFICR1PEH79VwnMegRCXVl8xuqilcgxLgkh++fWkeWvxwoYYV8SJ
vdtJADeAqEqoY66PGfHv50IVnsI5a6JlZn/aMnu/JnTUrYFcRlJ5r0uAhWhdzfl/
USnQ4gxGN/iAAvLr3r7hsxGOcHbaNdpL1SkprUPA2Z07nO/S5MfE6lT0v7NMWLob
OdfvXcV1QrIoptGuhbdOtnRzaGRCxvlvWeIzevR+EtRrYd8hBZpxTUKauymQROfV
qQDDOjIx1FDOFYOXWqhG55HVB+UnCCHy198Ys2qQ0SF4EBcy53bBNKU0vOYhh6k0
cW87YOufzu6CkofyOrc5mdzgtRPiK4KkUfR19ZsJwYxtwSGkDHf8HC3JGplL0HEe
y5rJ/XgEXkbAlw4VpHkUe+KILqIk+oug5zUXKmk59Ip69wxKwISlh4/TsdBLdbs1
lipvwZ46fDF7p01kLzI5wA5prQLE2bQGoLnxDur+8r2jrakDetpSVe1auKLQiEMQ
ybspOyItUWmV5NGhau/WnUSjPAt7izpNdmJdwWA/iMwHXTrkhCZFqdSFs43a2/B3
1VGGGnzaPhCWaomT8z2LlnU4A1na+dfGati1xY6RkPERYUfQ2jVq6hjKcoBsXYyn
NOuUzcRYJMxr1y9qJkdJn1gQ7j3tYbttg/ThUvsRDA1juhtIZmUBjVoyyl0SZStp
oi5bplkDkmHT8nlJ1Xi2sfwDUo9fphfv4eYFiQyPWzXYMGaf4WVr1OnBBUzyOoaH
75reHUqtHGVG4hnmMn142r2RsRXE/cOZ8ScfTO2uvqvc6aIWKcNm+VFuAQIhrQan
Heh/JRdUjOIpt1hQsLbxuR3bVvRFtggpjCy+hAN25X9TDc1+zJZEIq/xZmyAAitL
As3sV0iDbALeAV1KYN81d1/ZRohJfR5bjdqNT0YTfFuyAgibIKPzeWN8mxTUAaSm
wqkzJETHCE4CDw44UYfCMXYcB58irKYwx5Qk/mtskAdyvhnKlY/Brbr9wBLGsNoB
0PDo7E2m1AGtGdKRlDmFaeTmkraANJVO9RqxdXNVQJHbaLRfoDDRWTuMjBQcv01z
rjijR3PvYPLYm4ED1fEdAv7UloawOvsTFCE7v/q4xtWteku1eUOFeNIzQ6A7j3Qf
pa2ow4NttGoTzgV/SHPcRbDPJ7lAiRnX9PwkB5BfpAJWtxNtQEIolcQqqQ4HfBUh
3lcI87X59/9vvSurprpDWP8TlhtyYDlI+V3ZZVUZre9GhNr47obhzR3zoYDpw7sb
+HfoljCzP6M4BKP30N7FApt+wE+cxG7U7f9cB/jKd+/l3lhYDqp3dz6lO5LDqeK+
ZWYf2u5kSDXXpYgyC9JKVTsHvQmHT9cc9TTcN28KZSeeU5+4iX3j/7uNljfqRQPr
BPJFb/ThvU7IzKNcFmRR3H/MUSWFUBhPv9U4gZ+5uT5RuJuOrf1DdppDkmAEZjeW
ODxp73DVPI8IyA2Ketl+Fuhaq3KV2d5zvkWWv+tLrpRdB4kpEECEUyQgeWp28jrV
G1kaBdkBkyOVrY59oeEPqYr4mLt8ErPjBXm+0CWmxppgC2N1pG8dCj0gWhNk7wuR
+YuVrG8B5xcd0zSHAtbH5aBonPBNyie8ZdCWEK1dUM7aCxasN0CJGvm7+yh3ptJT
Q1k/DRvralzDcOJ/JrD4DHVpeq15nVruYyZYJKrDmvS620DronwluJBT+8wgGEgA
JwzlTrWRG0YBuu31l+xrO0xQlMWZJykQzV7lVcOHTV1DhSMi0/L/zW8CHJyd1Dce
TBDZIRmSBCADg/qPo67K7JA62j2Ud6CzT9GNyeABKmL4jVhv9WEY9V+0ou/LSMk8
Dmr/kvLYtvV63wUSpoJ2etxr5i3WyiAYBO/58Dlczp158Y0HGLS4JL7I5C5WmC62
tqccoUzhOBFKNak6DsHEyunhNRbP6No1N/iNSUfdaf5JyFO1VYslJGCIumbN5UnH
/GMT3McuwB9HeKXg3SZ+4e+bMKOevclKhkXGJT9+pzKr76eMjfhI+asgksJKT/8q
3LU+cCc7+/67Ii+22dr10jExtnYgOqKBYmn3lp4Txo5lk3ea78gxBbzcMmgWtcmn
hZkh3BTI8+eBnP6LhW+YK3VYOPZvu85v4wHQQ1UyvJGEkRJc8DkHuBqEQWNy+iiZ
RozQ5fRRRrqrUAdAswZjhd8WstZU2cp2W3CaEJI9f0Nck0eq4Ih1PBigI6jnuw2T
4q7UwsW9nLC3S9SBf+TbNlCPZMEcNojZ9sQ3YftQIlXk/WWgQhlnwyB8QM6WPibE
G/0ZE/F0gsp6f7sgQp7k4El/aEn+X50m7teUY+MMBf8SlHaR2hrh6vX4lhp5NzzD
3qpI3As1PbHgwHmLn1XpU7Ma6/WcQ+pjwhZaWLWImo8ABYl9INnpmauWVisaOjs0
7xomw5QACoFzkXY3MuNEMDki7AiQv6+i96k2/QYJcx1yPXu5TG13RA17jWwsfxHy
4L/qFSBzEIRv6NLF3OJOhjetQeJPnetMh7g7kH+50WWbpLbTg/n7ca/b2aCn9vKe
Kh/AsDwY2DxdZboyR6J+xdYRczLdmC3k8WsPniZslIPG7WFKWu1VhzJZAzcKjFiL
xPmNU5fLiVRfSu/cH0Lq16g753aHt1Tjp0w3d30IqdKTweIDR9tUTfnu9raL5cPm
j+JyzCP5ZTNKwZesjhn9aGdio9jUZ6g5NXLgSL2F1Ai1L90GYBph8ii1L9KQ8XX1
WsZjPhfZYNi3jOBN8CyUL/GYJQx89U7F+xi+xD5uCyhI4tZ8U8XNR7zMnItjujzL
IbI8S6pWXulg9EaID93icNRlklz3mbphTMCR5bhrY5hdaMzxmu2oguCMH/nWEgah
DQW8AQHPUFFEsKTpZ1HFQALQ8VRbqnX4JG2bu2h0lefyJ5icNBBNQqrE2VNzuiDj
/H/U2+v+hOaOzwqK1eb4MNJq2qyipvQX+lpqJhWdkBhBMqcTknHg+hlAzoOzFFbz
cEY+niUzrhlGUOvL5oVxDglTSiwqDKv1yM1+rR8TfCKWCqwY1hbVKnAdVxaBYMfQ
oJNy5UEYd18n0Zp+TJHqR+2hQOcq79xLJlRy5p0mIr6nmqR+Vv1ZKgBBHG7YPzht
sOZTJPzb9oUQvOdXFVeTPcqEflkDFHBqUfOAbCp0Wh1JNC4QwqUPt/DYl7DTda2l
xjr9Dlg7ecWuUlqFzU7XbaZEUptgJyDO4cPdoOUR/LiBqVSHjzMuekFlE7DJGUVL
FKc1G3l1eTL9CqLJ2IXhThcJ4H+yjqzpMsPVc/o6C54qxglIJ2IiQOZS9cXoPwwP
9A/fNs01VzEaViE8sVO+s3+7YYWhARMn+v2U1Vydb30FaFM6vRs/aGfNBwAsyCC4
3TzLvbSRCvccebe9DulfJ6gBwJJfIa6f9swPKWfZkptsHwvTRGy9v+xtR2EUC0V/
9NlVXL56P6lvQYR6uWOLxpgVxUlD4Cpj4W7Bb4vfx11MEAQ+q4Lt01VGV4c+rFGl
udaljSQH4irEEr/2PsHUiPuPsX2CwshKPpxWusm6AHR8411wgrM06y5sCUjf3TDl
WlYRP1nSr8RCyJSqjhNxYVRPBLZdMf4sNYcK7Iun4OfyaP0iJO9Di5Z4iSxkQw5s
NDsndlLa5J92Sg+JnChwKPezA8dmHyQ1bIVJ3wkyVHHZy6QiwUJ0kKMc+B6wrbSv
9KcLm/rzJzJYApbL7OSDwRq4kveROydmw6d0/2NJh8hXiWPj0uo1/JkUdsStlRKc
h7sY89g5MKR2YI51hY5nyRiHspmI/I47AxMSCKAm8oAkh8okAW7ptfO0dB6jlJ4S
u0pcCkvFHSgQt6/FecJpYvjQa/dyKTv1UwEjA74WtlGq9rd9Wzb7l31SL6qfsULj
hu69XqMx/HLAvQJU2nceJTSC50l7zYqsuIhCX3nzliXT5loTX0nZgBvdIKABA3gM
lZqiqlL9WmzNwit54smeJw8IsKv4mcjctlPy5K15Y2sexB84Y4U0yhXwH2oGlkm5
hdi7bC2ykLsia323ygRmPzbLMcj7eeuf0GHEgD+sk+xQh5//VDeCj7YWkskv3/nh
eWRJ7KCBRCxdmZOOBGmJ2nvgbOBM8XbVN/2KURQlT2Bu/9sJynQuwgckJFfr/Xb5
cfrmEBOJyMS8lWUjcwc8ocVvFCCqDdSIv6iycHS1BPE0A0J3KYNAU+GgPuroVSSz
AqSC81+4oLDlRERN4s0E+RJv7z5uBugjZVfxO4PcrRyl2foh2iYzkR2ZH25BnCGz
xiYFE8B8eJUdXFSx1eGybSoRNlHPv7LwdBhuaUWxLct+bvN3u4PDeMR6AENwrg2E
bI2N1CsXPvRR2n4FCVujSpaFVvu82bWI3jEbRG/wVsy9dm5sy64VLPcaaN+Uc7O4
Qh5Ip0ZTYWXlQpEAE1AdaI7P7IMsc0xqsBVdWL0ZCinbBaDtJsVB8cYb/eftkFIN
BABzOOISyxWxpqPbHQJ2eEdKoQzSEPK2iwQyHVV4DDfh5Vu7b9dQta8BvkIQMj5r
PlbyTztrLUuPcjVP0e4s+O3cTCivbYktwBALL19VXuHy0rKQrOoH3fr2TzDo32HU
3dTh5NizBUvZk8h6f8EHD3Z/uF15kFT+iQzU9lP9yJDifPmlBNZc67oXZhRlr4gG
91Eirm5Ceyi1R8XMjfgk+V4LJBYsUfgIOgkHn/Mq2gE+wAbccF3y1/Q9fZjwqhNO
efnNT6CZeEXGgUTe64uVtRsZezOEU/wmVMSRB8/suJGpyqGqk4bDShRjFIdu7hvW
qoUKYUqhpV2m9+QKCTHHqzwsO/a265wL4QwlQBBvHnb7/sUWLoAaemIh0yM6sd7+
2Iv8eX3QBcjNat/MtrFUbP0SKCJ5Io1opVImR/eOkQbUgiFRamVEV5GxBxk4Wc6S
vdBtFu6MzFd21d/dONKSQtsYcNjOyhidzdYOgB75IuVWw7b56Y671GEDc1qiGsoF
9WuXrHpjrd2HudjC0b8laLpMrCbCQWRawH1WQq3miaouYsIaBgwarJ3aBISLOmFp
ioQ3xKu0o/PM6h7XfxiMCiHykVzyJmyngPCodT5h9/pD5JG8z1Akp4jgK+3H9p7x
ClBYFSgFAjeRcjvrHEwAdUryCVmZm1z6NWJIRIeoA9smmJqrNzQKbNL7P5B0d7QV
5kWPz7O9N1Mi2f7OYQAwe1kqi8n7XMufAcX/4v/t678NRkNn95LRt3yM90LBzgoB
NLEZ87meNB8e6sXv8RTxn3M+mxvl7q6xJBJICDjXo79VJGeAawxaPK7uqXJ3Z9Y6
xxtX4X2y9Y8nyTDgZ4DYQLWkJosY5CUut7OWrfVqNIBEckb6+UqEdI/LHElzeUkO
slK6ThtTatUwIPAOv1xYpc6RNG8DZGuZ+X/waabvuKfvGha5ffXnFCiuwCNVRw1M
ik3tF8ehIri5LUw3LIagYejY4n1hsDT7dkw0hK3HKm3l/90iaANZ+mjUEpgnF7mp
JBPvQtkgipvY/GEteRPZtZJh1f30V6zN+yfchW4sU9qdN+U85UqUdodw1SG8Y77O
kIm+xsoyXEuNUCaBGLaADgUc+cTxkQXxNzKJ7WzyYSxZUMQyPEdRulPhuK+X8JXB
BinsiVDXC4uOmsmfdUMgFyNrOrpAKwB7ToYzBulDDM5cxrgeCXVt3qypsKKlMZdU
7v8QY0Dz9X8gWdRVgk0R2twGkpXGrwOSA1cIBfByarP94kxN/RuI0XmbuDSQZAcx
BUWCrV7ObhTAALsUJE2MfH72yAp7GOegbQ/w6R+s7o/YsTbiA4nGCW7/cADHerKN
PaCSegWDOrJ954uz6vduv/23EmlThKuN77iujT9uBGadB0/Kw6MtaD0F78A2YaBc
ROwUa3n9gpFs0F3p7kTVBRQgkh7q+kMP7pMQTrmyLPyo8wcJUq7GbDf65tYBiRUh
iq15m8uw9COA/C3C++p97czx0yZrEBJAvZMcximG9rk3lUCr3qV1FVQSsHKQYXTp
ADnn/FFnH/m7OtXYbZm9ikJynTOYYAccZkIc6Y5ZvxRM+C2yLrlZ5useu9I8LBBl
XLVdNYh13WAKAn+yE78LDXnE7ertx6fNsp0FT01ZYCzzVBcYcWi3laMGUnrUon5i
LKRnPaM1hPW7aDqK4tA+6GK8pmIonvHkXsD13cU0lp1M9v/oArCAAfRkUF/7ZSKX
prWYYxab/ilI8ZpGeToF7FZ1tKvOL61AEMB//+RZINaH1q0ydMCRl1AUgwXA7j4R
EcygWE6tedEaOvhJJY/8PQjsE30lYVVsJjSQ3gjregVx0uJx2mjvWDKcEqnvJ/CB
tF1N09qC/2i3QI4k05Pw25VJdZfCNO8b3DNSGxQezqC7g/a2OdwmaXMq9eLpHHAv
dS/aPTR3h6x7k6TP38EOXfkNwfKARbZ5zU+Ttv2NILz0O0eqQxHQNnD1np2eMUP3
YEQQZ1Iys94MyOyrP0VX56cahTf5J0wJA/G+CaP/UR+4ZBcQQSROH4yd59ZrWtzI
x9BUGHVjQKQbNn44AW07gtSKtC+xBTYVdOgZXWt28XaHy4ryUMXayhz5W/Q46G6f
0cjYAG+UwS46p5MNiag4Q7dGfYMft8HHmFPoCDhuMgbz0NggatDjiXaYzZy+s3BW
OdbWRcakgT5KVxLa55sMA01LVx/l2VqXztZ9EMPtScqvA3Pdb4PTVNmJS3X2y0Q4
trWc2xby6TDQHZduiuQLRByu3zj0fVg5YlmL7kNpmDhrfMV0nSMcXP5qzjQoflFf
C/p+ZTIq6sktvLvc+MVqy76OKgY+FBXJDN3L3SYZblTDyk/9JcZCv34krEEi2KWk
ZS7TKpsZHmgEbz7L6Q9t7QjpWzdoTh4ChBhgakK+qnjTEOPP7Avgc2gxGwvbFS4O
GGUJOelDaZgdwDUtlYI61byMVF2Zb99EITU/GNQYxfOVDKTQi5TPWeAjDfA+5qHt
GZofBarv2SjOTVUJfkK4i82yl4A9HTbGd4wU45WgcnnqtEo2nNJOVvJbJqnwXmQK
L7qTw+KGjcrFpmATp2v4L8oPz041AmNR+qirWtzA54oFnXdmBA0jnfwDPUXJq9dE
ra6Q/1FbhnVuHU5RZYtzkiwBBdPDkkOXT7dGzurpqZQEIiGXGBpdwQk1tvM6+TpK
FseVyKdJW3L40DMfCL0UWYYXkr/7UypiUWgHBvic9qI8hZXStljU5qPjET9rc1ZM
yPg94vgxFtDZEHhZ52MPoVN44caTsupq3D+Onxnd96Gupm5/adM1u/ZDeD/B/MSz
/P3dAiHhqPIx1KWDwBkDJfY3ZfijAoIUufqfM5StuWoUBqYOvIuh1bht2YmTS7Dn
EvU1PACdYg++YW0wDICEqkWg68+Fh67RJWfGQ4cBqYTdvTP1Q5SI5Yiz2IarmKyR
EMZAl8w+BnUqMQKxFvfmjIXTUQiCYIMfme1Z02X2SCaApLgfIX8n5qrei98wNxPV
gX23u2dM0QdjuugM7X+jmPJbmyJaz0T4s7wF6MT9QwDFQcmIi49Ma/gkL34CVfz/
5TmlF35XvC0BHKSH6jwzX7Z9xUWvfsvAGWLQZHv8lmuhUFGXPSVzaeshx/EkLHyH
uPI46zxwVGdumOuIOVHKgwPlp3EKaZvmIO91LXcQBbuCi3/iJ65ycBKbJxjKAdKb
8ThB7/c9E/6VPx+2r8QPmfB0DWCbe8EV11r+4EepGUigaNQNU0Xwlqz5kudsFYhO
R1Spz6ZRuq8BiUGhmx2cRzLuIVNYYvfXi/EfBvVVYZOj2KCnzjlrEVn1snl7I6Cs
JQFDbHjHSM8QidGd14N05yybn3yrUfWXBbR4vjJ5l4zfyxfYuuVViVSXQuNBKg84
bsCCp3iPOAvw2pwRYQXlo6ujG1teMaTsT8skjJLu2eQtuKt0n9uxnZYvuUzueIHM
IPOO45e4Cu6vU+uzZXoKG2ibfBdedwYl3dhauO1E2F3SmKR9FKPfXk9KiNLCUFYD
pATookTkcwjmDyQGhU8SKd1QjezB5bt+C0wEVAwhDiFfwl2oI7XoOiV0D7Luuapl
r6ESaVAf2q+D7WRuO2kMPmzTR6d5KqOKHwOrffPJ7saMIlxU/I+x2jjdiE4KfG1k
WB0fi/6cjIdRF7xP/HpWVFZg6ayNevhaph2fyBNP/5TPfFeAqaSJMRrF1mPiUzLX
+EOXKN1YY2msPZmhndtRpVpibwhvZotgG5MzsrXKoND+rbckTo9lp3DdPif7ftwq
n9o91rcmyvuhRlN16ABCtf56NPEBbquEl4DTwEHKGgdx7kw6nxDi+XKBj0itZ5T8
qf/5BwC7YSuPVSEFlkXLSZbkCAC2CcLgFfEVxbWCUiw5O7agOedrwXcQOxh3R2j5
+VzXsRMP9X3hIQ2QWqZU7HldghPUwuA92djSZWSJuJqq3F37Mpn16AgFycL9hDe9
VXm02TKgnnqXAMH9SCCEXKRpoDzgI2pl+rBZ0s+lCwa7Cw5NJIP0r5uM+IcXvdG7
59R2drymCvh447wG9985fc1pen/w80wvfpWOoMCLhXF02zHRCB7Tkd/F/FC3QdPO
Na1cYUFgrLEbaBE/2e9bQpm90xS4KOdl6v7FITIU3ohlf4TcY07oucHUcm5rYr7R
g7bkabNbWMr5C9o2g+fN/AIF9Gc66BcnB3GfcnlI7TiD3HTGSpPRdTjlssY/hHLX
AFpTPjARCaU9kTySDtzx4mZ899OwUYPqDTWrYhMeMP/JWnSvCkhHDLGeysQ7N8+I
lPqxfuOm8oRmsfsTsIM/cr+KKp+yPor8w6sCBtwGocb9XtN50Kh9G81+St+oJztr
Fx67YLAr7IVp6hTd1MFknBxWhcWjSThkXYT+66LS09yISlmQVsA1hv9XkEN0Qwjt
GwP+FRs0dJP+trXNyKasTDJysAl7sH8NZejzNUwl0QUsfgge3QAeKw+WI9cKDnji
juQGJISq6jNFDrBNT8VEHj0bYwlEhZFREfhhfiQVnjFk4Q4S6JZY4nRgUOsjW1fq
vxae4sP6e22ZN8qzSZ5OBZFj4uYCY6MBxw8mzkftMywyKT75DQwPnSc78r1EibWB
KP0EsUABgr5owTCZXlDWetEHT87MQF30Jx+dfm1ce7vKD5srHtuaOxXFcgmSz+ni
l28mUhUR7Iw/khmyzxt8k7LDh9BDGF99Hj7pEuhQ0F8vIfh/lnPuKYVujsh5PaFf
eZqkRKdfE+cIpZdHl4Tj5kfl9BxdO32quWdLXb1OHS6vXYLes/eLiVO/rpRcB+cW
Xc9Q4bmZU8xUiaYMe1fNjkV8YbJpv9vdnpFJLI/H548rABh+dgQIUzPaMVeYJIqo
sr8ET9KO05nEiZx7+1vo8vclthE7j+Qvnb4tIFCQS6nhDoVHWt66ofrpukwJBM6m
lQsVjzW+tN2QmXh1YXM5QiBTQuy080UxzWTSrIdxx4G9Z2wycgmQVgnCQFEJc1ku
KcGfV4jE/ZJBgvuN21aN9/p4u+iZpXRuZt4E27miv4RxZu5HcIDnlCGvuOzRAIIS
pKK4ZKVreurYBctYdRFmMpfQjVWMpnKq4+bQf9cjDsyKm3BKIOz4FW7dHMGLK89U
bzzJlBmmyPA/zYdBzz3bzxUv5l/dmd1bRoDeEMhok7x3IIcfjRP6pmi/7xy9h4Eg
RaVMhsV5YfHV7wOtPmm16qcB1PuNMLmIAOurz1ieNH7bpq84wTDzQoU8iuMlhJmo
66lsW3x7s+gU4J5mop9+keFIT+wi6Wq/nrAWvakvJ3UQT8r2+5XCqRZxCzXMU+hG
Q/Q+Ul1oj8TPwDCM6i8xxZCklkMtDB6bXIaeNs4layb3KDsK2d5sG2B4HpRJ2tOj
lJIYSWjOWkynfV8vZrHifUW6fR3k7cAHMfUhjRklapGds362w1nvUS+kp3lK9gUJ
LnjYJ9RB+wVwAavBX+AIDpSLjqur5Mcwtk8XExZX+rDUTFiKRauhxvnhQrlcfMx0
qgKBDWj0jd8k+03KbTOiLJ1vuCkxOgtyfU4rfYfwSJy9WIfRQfVuQQUaceKVhCfq
14Ri/H3wb1QHuj2N1aHbiqiOQDHZCGXeaIGAUTGsmgZ0urh4EXKkhGxkfNAmrHkx
21G/+enELaNVyd7KqUEjaFTHGHpEP0mTucn59qyXzR7qYxGWymZp5A7VQDQigr1w
b8sqDZQidFbNyAMRXETf425z6NeAAtaHBNrpEx7ka75/1QlNBfeIwRYj1l3Hsa9L
XGFMMJiJ/7yyllx5LwE5nn+LelsFr2YXLLU5Mowb/YFMGN+qbw7ORJAJgeXeNhsG
ll5sm7RrDf5nHroz+cslkjInf4POWwMEzHeo6LdTC6P6LDfkFZNJpcMEW1YZcYPd
eoqxO0K0Vf1n/+4kqy5FOf9N0X5W+DhzgQ5pSkKpeikE/509eeVauis7x+yRQZoe
Wg/D6O9dihKRjly8n7jVglf3wZzC3Gt/KwEZwyZx9+Qwf6WIhYSG8JdQShaPwMri
1OeUcYbYAXmrZuhQyKauXxbIJbhRb9VQM3/qayHOlIQ1qQTu6KSOe/mvMJKzR+75
eJ1vT4OTo4hvVmYhW2TX/PBiOSIPNAoaArrHdkG1kEc7TP6a8wYTYF8oMRogzNb3
U919+q73fbbGrSPp925zjBJxAtx80IHbShnCTjGWEAeYmApG2h2zMkxwPmPYN7bP
65Md0OTkX7eRR9tSxow+s29GHzXHHTzdsd1rIssnWsmGXb20+Fj2LEkH2+Y6Byo7
eFU+YEEhAG2Nl+T1Hb1BpdOlDVjIVJoUm3U2P3nP7bid5kbakkJ1v5FH/gYo7bN2
VsQoucWetjTO+q1/ztdSSqXEhQHpt17hzoEl+TmElo9nFXCFJ1Ip0hJInCxFJ0Hy
XxfULcdaELQVtoioisICHP0cs1FrGVHZr72yawVZWTAyhzTwyBOXt+ckWRo5Oead
d9A5q8iZgL3s7D7e5Ps0WvnbBud4CoNah6G4xK7QcioB3i1CDNzi69/o5wkvvJy4
/cIzJeeRB2CbiVLWEebb1BcLer5ZXW0rTjHdOtlIbCTW4631wGjP4081U8Q5hFlH
I87X0q15xdb7aFkIgH9SrixjK5cDahkstK5ZqltVGA5O6uz0yQxStnlux2t7Y2gW
gWx2RjmhhDyTWEpNQzM42laU1eSPwO8hKZ7mkObhhAG3K+yUBo4roO92FUrKAWjU
a96G9Ix1KHDojxaEUFsnSQo4EKaG98MTyceMdRnVUVpxfmL7xFzgzawS0ccT3Xk5
SFUhNlj0W1kQ9R/4CkmiZ0xWoV5SnBkInw9KMygFANwcpgxFyXAqnSknnHdLEb9J
uWMDyjPnSasFQOi+jFH1r3FAdPQpu11q9xDnut2tQE4bRi0Qn/qtn9hoDWgPewKp
Iehov+kmxLpU5LG2dY5n1uuYoffZLAea8MqzsiWkvrsw8kIXTkXXQEW8wHY9ibTD
sMe5RtcJkBnzX/tnyNzgrsnieSp5iobZU+Lrcb+xMbXUu7cvM/0AkWWM6OSHumDp
bhmARYHZ4j/6aVrPr+eGeADuDSUyjkRXHQDjn0b0E81bN2UGmL9VDmW9who6uAGd
Jf4moXaO6frT+QODYEiEq4DjAWqwdtI9LfV/zU7hTkh4SFrVceWJtc0H9Z9VfP6w
ts4IKB5+3bhoggM3Xf6D3v8sBR2ehAXNqv6uYTFSrjRv3ekvaf5S0wFS4b6tmKde
gwW2OAfnK363gajTFeOd0t86xhi4sTVoowtPLRSX9BvvHFED9cenHDjcrLw4eYlO
5lefSlI1Dj9W1ENAJAPgvF5WAZvzliLuKEWgq555jiVUPWEGgAAe7+q0ytiMK3+m
iPwZ8IweZlYuetdxe1AU/YRGW/UXWxt4scyCmnh8/lGtt7uJ3o2JbOAJ61B28eMi
kJxIjuEllSRKh/W3SQR0w6uA5Fe5UrDPql6B0HE7GsOFOY4fdy1IPPzAzazjij3C
EaKyU0uRSbh6YPUjELN3dLcJDRY0SkIuA+eFPHB+a4wNjgGrdJw6Xa5KsQlV6YSi
3BvYimXRyvFyDNIJYZwckWXXj7h0VsM5O4VmE/micPPkybbKSlZU/K3p8F5744yU
P9nbnbXPzgUTfqAbDZyIj6plzVXmT0tHA5yeyFmHUSDuisIamjo9IAFAWboAqm73
dDfTyeSXiVaGHGjaDf339PyK2NbJG5rFA71lt8ugNoJRpNUWuzTzJ9QssSr9uD4b
m3/AYssqgQowKE3nwN2eX7O7kbNAelv9+B8KoIPxMEEx1L1Dy2OoIGO/I16esx1O
ybNWt4n6lF+COFB/t9ReetJFVYXz0ZoLe8MGBpLVXqD+YW/vXtFDAiknpT1Cilil
AYA3BbUGV+hNzKmMIYbJpYqH04ZqjQs87ne8r4D0F9rQMPTM/9aR3RdwILllSqSi
Db424GaWL27YcCvYqh5yl98Q1zi726nvnv4i+LoiM0sFeq0jbAvNf+H8uYnJq53o
zbpQGmtq+p8P8qgjaK5nnApb0Ov/2fpBEDU698JH5Wuyo7QRvfSsMwafegKYuhNU
v9RWqjwodwkqjOz/AC8bif0SPjVsnWM+yDsiLkMv81opwDumNoIS/XNF/vQXpk91
N5CRgtCbm1QkPLtx3B+uZwLqyfYvwxEM70HOTPZ14n5LOFp+gNYjZAqjmex4/o01
Jz0IC1JsaX+WU9qwvTrH9ASBxrYwyy9ANSSJz/bocqSHrM3pE0eYsB+v6H4nmkal
pZotIFc1BEb6L+kePG9h1dwfdJBgKuxmPZKbDy29D4qdqTs/mgYFgDIdVp0v2G6x
GBtR9keAF6qLwstl7Qq3WE1YtxzdukOQTryuELapPiS1zTvLJCz3gXlzK9gv71tS
5BVCiHFPNNLDbSzFVYGoJTaVLUwIJq0/DGnL+xC49vzYrYqOQybyZ9Go6s4pjMF4
BeFhhVXGJ6HX4fsOi9oIc5hotsqALl1ERaQBwHqU0eWNn1dFhrVCg5rDdUvN5h6V
gfHevl0esIFcAasT/uO2JxmevkbD0KDS5o69HlRX7toyvDXiYPdiNWRYFf7yYvB4
wDR7rzy9bXQwXi+y4LJvGAvY9N1+FFXhxKdbN07dR7IvObyiz+jSEpQ8UIA7XXpR
VnQshISK4a6Cu9D6u0/qDpg1/+j9t7dtUmjMqktUvsfsydQvblCROR/6HosaQNfB
s9wazAt3IL23QXzczYUcJO2CJBe3RWIWNLXdYx6iYG8/1iL/Inol/+Iu+/zOtAIu
Y0nFO7sSKR7cIdoiu5jfUuYsNqPwJRkaPmctn5JWGLfhHDlhqd3fkmAF/oiNAh0K
/Gx/WtD61Kgfkrc45wa5BHcygDZWXIpTgz/CFEPEQWRR8M/Iue/WLLbredH9e9W3
ZRxawFa8RrolS6+lyjtYcTErPzw26D+xs0AItdhaA5p3kk9SkECZIscvCJo+C+vI
bHgDfcLaP4FePflU7/tpcWwK8OIVxVwK5ksoDWFAyEWV6FotY02yyU9Qc7G7oSx6
BXtV/rr+SY9LeYoO4LV7wb7o2k2JUHzxW9XTbn1YkKgTXeBACGwZ+Xv2ziPImA7+
++4qJPaXf2XDjHSohpJpgfhuIjQowR/u8lZbmIBBXppPhodhGo6NeWHRl9GIcFmT
BzYl/7Knrm4V0TjeoHIriP84tsOs7DGaIS5dgsj/SHdh7MymZoxzmZiX4mQcU1I8
NlNjYJJbiKMf9HDZqkbhKbNhs78l2icYZsZf5lyrBH9FlrlIRoEse1W+dWKTLZzw
7Unq3S1v4Hint8kkwxlQpcwUxV6kJfTCEwoFu9tkGqozBZ8BOgp6W3wwkj6kTthJ
NsZ/PPySf5frCBCnn1ETqmN5mZH87wjsU626HNDzID3uFieW/OBZauU7Ni02nslU
/hcTBJzMZGFLS+kQPYtBf8xtPTld3Az/k4bM8rB0BqvxGJuQq0K9UXbQX8S4fT/E
7LSBgPgWo/z4Ly6BrdHMX4CNPzA9XowHP6lM2P6Ih9U4uDGV/Bvt6y1qEFN5vnSF
83Kd9qVh07TxYpzn9dEFaAmaySmjeL/1XvRfnjOQ9gHhxfR3FgaxtCsN4UhXMWLz
2x/eqPZtoqgPnl3bhACSPX35oyHP/2/L/3ive7Q1N7x2IVtp6t+jRbVl336ILvNL
Kn36wyVFvY35q4cbbeN67EU3En/ZbPq6yQysr5TGAAKozGtaWXus3TWXM+mzydV8
39/br0UISHxhO+8QFDxwBg9bVfVvdlFvjMLZbq8fOadQdOToVIbMXD7jlpQZUaMn
3Q2OsO1jBhKgvab5C5rIdSiM6Z0oyj1OqfHETmTgfg99HG2Fh6qe2ynPh4WyB0U/
8ab+NcJTdpYzEt9OikUOt39H/gYx/jD/LWpnyr9Y3rQTU+kxixKmRFW3Q2RkSezK
9Uxwo1yVA64Q/3HkWKnJckCwI3QfFpyOrqo9eQPsAY/GYSq4UWdNGa3NOGUPC0Fc
QdV9Id20IDWF5nszdmMBsbkKJBKdA3tLYrDdjjQA3uOYFgxpxJRwe0zwsuxHN8Cp
ounRZ9IyQn3o+IgV0W8bvNJcKfyERXN+sjwBattfJ1gRnogIS944w5d/ZE+DCxS0
m8BrS9z2lM0sPZP4qD6eeFJ4aLinBzNEJzD+qzSnkto2WDP10PhJTQDbGMgrXr9u
wlmvqBUekL30jqqpl7+om1ITA6D5v52yenyvAKHtPCf3ugxrW8a3N4XvsuszLAA6
2ZQbSwLDli4HqXQynbScQNpK5M8RgmtJebK9oqS6eyYBxwhU1XHSIRwx7PA8eaMM
y2nxxkunlAyDwnE12MJ4APTqMmV+vJmTdFuFxSyDDZ564t2knyIkZ6Xr7H/UJ2aM
96umRSofm4CzVRVGXn+i07/HRxlv7ixda2zsM/AegU2ui/zV7l5uBRtC3WZxYO49
nBvGf5QevPJeI3ad6OVKD22D8xH7YRGDG6Otq9a/cwiepq+PwBS/pajz7Ol5QM5a
PMYRwk5tqFqb/cF+oQCUSMRX85tUMBaIgBi1SRHTMGGD4azkw97Nrvow9L2WN7+Z
XPBe7DOt9dscxmRJn0yJom5d/P4QBPlBQMQN1/pI8QfClxrN3bw0vo4eKCaY81UA
FdmRMKpwIA1jw5oMvhj0Au97+Yq2QBrw/z99S3vDRPotU87ncrtjclrdK/+3L5wK
pjl+BZPoHrzi9s2mW77xCe25B6aU2LYvQjfN8bCbCktdUVmlmExf7krrlzQD/KWc
BpW9RsnVuwZhKWxf9EReLydLpCJttdNaBRbU9MjoZBGrPaGiNLuc7WdP0KCB5FfR
VikS/2FbfxiMiIqE2XPdrO0FNCz7SJzNBB9hhHoTbkkEvI1IVywJ3gKljYtAiXpx
PRBXMuE7Yu+yfFoxi64PaDkIImJ6eWURobS7J2Q0ax5ZkcMUgkgZcNqPJCGTdYDw
b1sf/cKTll4ChmmR26uOz1cPyGqoHXeO+QFWWP1JReCPtyKgkhYlFIWk/xp5RBC8
JwrQMjQ1d0ivppn+eilJgOsOIs/j+WADu65U3oA83y0KuveNlcA7iWKY9/NHGrXs
1WAHmbfgGCwyKlIh/D7gORHDKOoWp3IHp3BZV0j8PGJFyspBRkmgWZ5z4yGf4/2Y
6JcChTgGD3DMsHw+7oEbf/JiQLKMkY/rwSyS1baSN4p9f4CKYKO4ZpSUChZDCxMn
Y1S9ErWipAveUxjsuDRkmLVYzwzVGXWUC1HSHUTYUtxUp423RZXFiKZ3zktWXdx8
2kaW1rUwwp8ySzVlpVKpTJMWkrib/IP6rP5MM0oMPbBMfY1ZV1GthlHdJn4elIom
sCLtOca+U39wBChfYcUGbYuxXsid16WzOyq+NTD5n/zvjglpUkeLg9nnl5+iIZf7
U3beQZL1xnsBewn0/mDIlVk3Y5NY2XWUUVv3Ke+kaB5VYCDfry6WtNZ74ndNmJyk
/yEuYFrAdwloWzFtXCw7Bvmdlg3pGDzYzO0Dw79Lg96qcA6h8H83W7yk0gaJjU5v
LWn0y9IVQchXpt5z91FdXmdKuY2z9/HZXlUSpRX8qqLhtIPMEoO31Bz13ZtdEGLh
zr1fiHJ5MPBI9grvFTuqKKnQBEwWeDYYK3yoRKademmyGi9sarhDOkikrZuUNf9r
eWCenr7yO3QGBJzHKA0P/YJ6Z5vZeTLPxtH6sC/esNSi82Z0gvEsLSbnmEU1F5j2
w4ilcgG2RXENqheELJ+Lu7yA8BTkdt1jlcE0ov83ZK1JM7Gycpl/EubQnxF71PoC
1VkfTLy1SGvJISqoHPgrVgZotY8g+7++OF3uwenYjU89+m8Lv6xJbywANDqVtGsI
HRLmnhprjnOkOwH9NScs+47u9bGcxmTiD7jqGZDhBQ8U7UjS2mx2FUIPVSfjweLF
Xow38Fr5SvkldtciM4Bl4oVi45VR3+WLdxpJ1zzmsj6Xprg6YoqTDgTV1qbmvksr
40MSTqAH5eBkfgRixbJcOIxKibk7qPXeLra5rlFArpKa++qWukJ+7434TrOgOGPS
of+DFAO1i/a5VV5uJd7edvY3w9IYhHrswfecKKnk/OnmVVsNgYxN0ugIhBCufgmp
JKI39NwAggAhnn9vvZSsAn/VQ0o/RPrCzPADMEEFUVSQ00p7DaWJncDCBS+18YgX
UwiMkjPH0qxO5dtLT0obcKoSgItbBjQ7rJJm8fhYf/PyRkbL6qXge8UlAHj53cnS
dpYQSJbW84wXODOZdQRWGrUUEYSXvadBEH6Aw6NNV8j8VtJWw/lsc96LpZzp4Hpq
X6uxkk2GDWmalrKm6bn3Z4GLBbGQGcn+DafHKuCqk4ogdtme4hmEbxoI2dBCbeGA
rkLE1kn852KPVVo+cGCr9Ia5jaE60FEzyWzbbv3XLOru8AqL4Cc1VR33UZE5NFzw
AW2GktvwhQPT1rYuWKWKl+NyjwdHCnCSw076IgN1MmGgc+8TSYPowhFl+pGzHkOw
NCmpTUusi3kqCZ1G3cetonjDM1q4fuxwqMFxNWONcL8twObDVvZRxCO8zVAQ9P2r
MuNk0UWaBAshK+ZqfIYtqReAllsNj4svoae9zLsuch/xDQL1+WgrO9+FFkNdHQuI
zbojHvKEG1aWdku2U7pLuEngcfzQha9/rNAIlRW3VquS++hZD9Ah03kopNjLxtOT
agjuSNcJ/pe9NrsQX7kvD62j24vNpl3oFJxMfchHf3s0gytQlv4Nn7EqHPUcF1kZ
zbKMsHmRb+lmu2NZsvf1XCDHRqyaq3LAORaxizPFCBkX7bGc+U7jsrhmGR6JSy+I
A6YiRuxXLaIpIdBArZIyNT3Ngwwp6Y6LmFIVpHbiOw1ExBiRFIip+jnWBXDK3BV5
d7UvmaaYRWDesVmphBxvRKRzz6Qh3hRuQGmQr00voLpDHIcZB0W5vfVHn9b4bqIr
j9gI2JGKH2tuz3TgOLAkjg+MxjW4wDg2+ZKnSm1xwMih6WE4riTiFmjSN6nm7X6g
yt7x3mDM+OOXKeXVd/aLaa/fJ7wV6tYhhOu0xMd6vZRLHVhoLY1BFpyMy2XuIivx
8tZikGxXqkIVUNwUZuk1kf5RY5jWnX5ibQmonOrNT1lCfPkn0jQFaEIt3agX5UMn
uo74HANR0cRusVMoEXfivqmpRFDsrCqqaDUeDpowJLWEG40bLh67stwsxmiVKdj7
T4QKJksL0GEO9diFLr/QTg/ZXbxdn/857c4N03Mqygo57gfKi1bH8lw2iJZEytkf
3jeslsXomig9j3TxPwpLv3+LYayxLCPo7tKbwaFFG5PBuxcnFcTRAiDwxOtorB/U
bhNr3Si9Rqfq1l/swhCvMF8CAeNwfi4W/CTS4PXy4qUul2vik46KiZ7iUBalUlSE
EIUDF03+DHmG5Ck+a1wpGL+iyyB88uDSUmdTqItuLf1wR3ULB+AyXFLHos/837UW
z154TsBKxg5Br8oNEaq0hsSSIdJGTO0YvUxTiUApFnDXA1gnyVDiOGEPWqu++p9S
1UUvhKFMtVx/Z8gUjg2cCnr9Kk74h86kX9PiwslJIWA+vsRtrGclIgLfYGwyLmbh
c4kVJa4MJeADd4wAviBtFWfbFXRTKbzvGby4WnuBF30++02t1GhxrBsX6VHJ3wpz
L1xkmFYjNR9/qWYbHXRWj1Ht6OGsA8+DrF8COjq9gSzyP4eKSz07VzTsWO2qUIQ/
chkPh8GAMeMSO00w+RRgcUfc3HGWM6k1ui3GvAgbvLHcdjAsocbiYrh0+hY89lNt
DsTIWo+9YtDD2pPlAeg85yq+rKC59pIJhLfRwe126DBaKDObe7/weacjS6tqfE48
VfHSqYJVKG+1aH0wpreBtz67BGz+ebHxBhPctqs60HnqEeRrjZO6K9RGJ+/wyg20
wvRHsYSd1qspZJhVtotpSp9jR4ULP/8hD6VG82xJ5GD6qu05ucnT3s3ydKC3ZFUF
a73xN+XTLsoQjHJPhyb8mdJ+YVnx5fRUeWIOKQj2KxYLlcbnTneuUl9ECJKSFIg1
sDWceGg0uv3v5UX5KryKidsUhUfedRYYaP90O2Tl4o7E2GGDAGpMBdYDMDwQqeVJ
nOisHlGqSnV2fxqhN32wNx3bkv2k+aCBMVWrPxSbNVyOnMiRsf4BelocFvXrgUc9
oWAmeAVpGYgZZ9IugBGm56lOISaOT8LUvSBDCW0n89YAxfAXRGasuGyeCHNeb0se
o4+ip9upFE3vhdnpHNocqk2G3/1JgYLUaX3YveTZNCjxQZ1iCXRqt86xcwHmXNCd
AbcTOCtJMoGeSbyvt7XwaA4zuuYlfTsWoUAY88/pqKD+Lxu17kyyEu0A1wl2p9be
qbAnAM9jY1Qqw9ljvfxJck7xCfKCM+y7Ls5PAuMsK+iM8uh/KE6qmN4s7ce4jWhT
XO2nR3cZP2EVj85t27xRkJSzqtYPZe/CjHdFhuJU5D9bqd0NvEbx11JsGkFLQ88d
baxrM9Y/75H/o50tN7HGhvrjXQHVW52K0HivnXq+bynOoDi9m8WsEaRl/3PSt5+s
DOUsPeUWhCX6JT9ByFMdt7dpa7l5m+YWJsUH/ekw1xwh7tU+iyi7ZEtp7iAHC+hf
VxKoJTpDfrLZxfejaoRjkdXmxi+3D52IlGm631E9PIAVd//dpkJhaCy8Wm1bUBml
brCAbeNqf4qR5KxF7dWtT3rxGt1aufPYzjtEkZEflUWYMeeqDvKVQqPd7fGnLQvg
CW4LpfMkQtMunICnTo2vGYBBNBZFLqsiGVqJ4wi68pFkWIpcLv/WBRe2sksPiH50
X2yFTqVSHHHlcW80f7JU8ja+5ZjQ+XB+p6n7u5LJf0IXQVR2/tGTfUFh/OIur+8P
olPL3Gxye7mAyy4qe8JQ2Uzw6nRcA3tMxhCunhGQnzeyeH+jYT7RjQeiUcQq5Mnz
uOiDJwwL6DERYWJjtwwrGuVkYu7rL2tmK5iIHJcuvPD6FPzzReDqtv/4K4LmoXlw
6Jo9YGNReETWiREvUF/SotEnhVkG18Xh/t5k0qGXqR6iT05UOHtYYAn3y1uSKfp6
ylkoAr3r6saFUDP/JWiie/IiPChJJP7pkZBbJMPdZ1L3ciYx0474nLYE1Lyxo5gx
5IQ5ye6frYqHqEyl/0xL8Is1iLq+h8LmNNNublDC5BTK+tCVmocqHQ3wfxabnfzo
r4GHsKxLLWMu0p4pDxei3B93ITZFvoyNE9k5f7P623C9bsTtm5tTLVAIltS+nfOd
/ClHoMTwJfm8dNNvmiuwL3l5tiko/JcLdiDCnQEt05P9GCGC1U508h96HhC8BKRF
xZOPp7x4MBUcCpRpJZYMr255pdlOI0M28fZ8Y+Au8Wkqa68y7LoWivDJ5VErs1dI
h+lq4m33lJ6ctCDJfLcT9IS0UqohpfbO2ZlsswlhX9eM7jHJ6FDJejODxCWk0N2I
99RjqgXexueUg7aks2ledRFOMMQdv0BVjfRMpr5CMljeX+9mzuL6AgeJFvzoCEbz
RvA9lveJKgtnZnfMy8U7dLVrzjPZ/B6xDFbz96LoPtZ62ftlBncEH0BbuOj8JjDw
IlWNo9QiIosmnytXfs4pQecNrZQklPnU2Gwpz2y5kSQIRT486cdsyL519e50/xpL
aoFcAjDps2n7utTGaRMtvMyUWDLvTg9CETAT0N3cI+PnbdmYIzCnYKLT+G7xFj49
BSxYOGfbWqFZKLEgehlLixu+SQ0LiSAqKj0TF6r2TELhJtNNuhtenOjmUnneiBEA
WWXvbrhT+H1NjZuYV06YtiN5D3IsfvwASz8nKbgvht8bjzFutnmX/aPEkLHKfRDY
dEDqtPrY5HBFqK8dAiBw7YZ78cShqQe8bu9O8/7eb9UC5cwRUHCwTQ2ljLJqM1mV
JaTUe1P2eYX8QtjCx793ERcsLSRWvtlfh+XcapBvx0l1tog9clAE5WfUgHlp84Uu
2oG/onlmDA+HV5G7dS9P1nomoMUtX9L3d6cR7Yy7759a1ZL+gYno2vSRBY3RrPPQ
WXyoLGVlPrUUVcea6ezDvx+QxJ8dbaiqOlQKyd1ZPaMyML7Mn6rtDBX5S+4t9Ooh
XBG3Espi4Q6+oCWQdBAkrKutuRtRFibaGpG9H8HIJ0mYWStyLh0GW8g4KgLu+v6g
U2DVrVfupyX0GgdGm4krjsMS9QD1bW8OJ6vYvdTDRuwbjaIX/Hoj7V16yafWQA8Z
i05xNQInVzSljF1onwxsmX8Yn3j3WdgRMkcJc/h2WJyfxM6upSFLkrgViI+sMYcY
7fG9yBd74i7o4dG4F9j7OXy/t7Y3MlMfiA6HDLloOO39SkmUA17vu/7xzOB+ZG2V
msAmKClD8I11AfMAbBdTRIyr2xeGNHbDBy1MhnvdFS/2ValZkCizNLWIv7aoQ9WS
6LJGFuDThmaalgMQUGNSS1xCyg/iaAjpPFGPVxMbkRgIf3JZrkMlCiAKI28s9/KB
/KGu/v8mFTE4MD0kbTbyQ3tYKAxekmDQcskaR9niNQw8c/gULGnkBqb6jHlO9tO1
93lBi/fAaH1h6ukqcJsKFTWcQ4b64+6w2iPAWvjadq3LUcHyRdW1ReDLGATMmIO5
yYNbsxIBUlhWeSH87Z2m3Smbj7QSyhPQqnOGM7M9kF6Ujnf/2ViL3l+E68KTLi3A
jzzcP9qmdWbjnh7/q7PY4gmPeMzBRlEGVyAXgej0mq49051z6S0o95+lo3NhmxeG
FSO/jbXwioN4K1DiDjH/zoA06lJBlMnMQVUTpJzmhX1AnH2NMVzET4dTbzEOBMLT
QaPR6azjAgO55lncWaAMPIOMzg58HIFB2ZzFSDtloZNl9lQSYgVjP0tyv5YQFSJa
qsif4Ug4zyCJOroCLaUmKy8Yz2GCVwMfhIa95qHiPPLIAvqCe2xrFV0GTTb0OMmp
e7VuuHIZc+7i7gvg+k83894Rm4qvsL7XwqNMBG7lIdKJuLxSHHj3RrsHRd/mfCEV
cVtcuk3grTeZ3J7uUy8hjIyO9d+5N1hGIU/ZK9mLiJFocvBJsndq6mF9F3FrJDhD
iA+aeDw0FNVavGUjKY/lntTb2qWhCMgRjPtoQBpWWN2+PjlSwE112vqAZfam+onP
cQpOHniyqsEBbktvBo7NccudYBW0PrZyi07rWvpnQqBC41lV4u3ufsMJ0zOFt3Qg
anw2jyDi3f8OfBUC9cD8sxF6ryM3m+KEF6IGtogoRAsuq8mdS3J+BD7WDzpP0Lr0
uUvmaSx9dAwhRgOG2fNHVxGKt5sxRsGOynnOAYOz0qHgUnQdj7Dv9vURDP+K+VF3
Ra7bTj02v1GUxT3nwd8rwEmyI4H+uVyKPkFYFG9lUPIICrTwZD3ZhJr/GsXqr3c0
PGOEdcwOYYpvb0m4H/Pd1ysi4KdhSA5h8yG4AAWkS5Hff/VA67EcDMKul+evHOMt
QMlWUe77mVJOnRZn/697uLAZx1Z3xib6fywCsDcvcZ/tPhnpJnFA5VX+j0m4nQAk
g/d1EojLJmvgjpjUZlj/zM4MLR0akwtMITEDzJ+2mTJjNS13Tq5knoPKZ0ibIHb3
C1G50DbOyXeTUddYDKYciA+P3l1e8d93FfAFQXcpJhvm12/PI4f/I5znliKc5g+V
op22vFHq/fQYXZJmhq/fdBNVcBv8XnTEafkT+30SwZeG45DVteh+5U57Ciq/vWsT
JNYf7ps5nHbcXvaBfJrf7NZhhpyVORjAawygTOuvi9A6S2FAched2WTOvewkGBIG
68EdDwa6f9iL3mDRcvI8UnwTdijgbVzAPDIWcjVVmtof3kF2gbehEbbQSlVFUAIC
U2bAkTYES4KSV5iLG7RMJoYtDfQ4IUsV9kQtCNBnWbnQ+OBv5i64IH/W16DVMOx6
EBtKOqlcOmxfTPgebsOZDYaInBj3HCiTt9JKJ86NiBeCKwNsBavjBGEX/mA7igvS
wv5y8KYtevgj9cpeMLg5SLecrGmrWCg5cK8P5LHhxvzd6Swtftd8GN5yGZRX5nzL
Fl/PtwE/6GkfsoJVqxYGgqRXFF179xMOX/39sYCH3iCG3v5YtJgki5RwBezVKaGS
F+QOSkpFi5AZmvFxBckc0OrEwVjfLqGWu1NJff8W2RWbYsSyeTLMO7PP27ASOx0G
tzOrnkevmcnspDLbYUHT7EchC146hcFfpxfv+r3mjYV4AmR76aU3p6nuP5V1rak5
4q17i8LS2oDMzQGgYjQIpnjMxiGOSpIpDFVMKexXbXHsp9tbPHM7JznoZzfmzBHc
zO2IEmnryWizYjmu2sCcmaT9zEkIJGMkUJV1x9wkvLZdZVWE8ZcYhyqaAlVWLJ2W
FZJDpeOJ2SBkzckLU2dM1kSyd30hTJzW+6Rt8NEsKZPXPOolvRmCVjESRNr9cI3E
g4mpk7aTVu+UQ+79IfaduxSqik9SkK8l/QIerT8o3X5biRbIxdijvwE9n3TH2HUp
S2Q4Rx6nb7QPTIhi9gTMeZUV6qH8WKe7jKqlEPhMvjIEvGJWBZ6Md+KTAN3qs0Ft
CcCzi7T0eFg2kFhlTOaoyNBdXQrVGYjp08IhMoQLHoL+9wYxErxdAyb1/5TY8AsK
A7WI392SkvLcBRJUHw5qsm+Z54RBCXnRCs80Q187up95Ys7VWzeyAsdP+wEEBgX5
fXfBlHAnc7e0E7SfphBKF97B8FDcA0A3bLUS0ogG+tY00OlBTy3EGGCHVpLWlwpE
1wA2fi2f0jqbJ3S8JnL8Hc5okqUJP2DDRBMPT9MWyN+4JHRrmHpZ9RiiKcmzPIo4
QZ1cgD5x7ijG8QH9OO0VEhm+crjbMTgQ86ep0kJ+fQzUCUMCluMAeKO4iIeam9G5
GXQWf0TDjEJG/sLYtzs15y8wkhaBIXqAdFsiRR8+0H6n1M2MIMmgmd44k9OBpjxe
9TGhnRP8tFFx4FSTS9DFo91PKdQHqOh1g9E7tqQxA2VuUkJwvh4uwxLpD6paV5bS
C1Uj8d6vpH0vWK/4LifzrbrDvH4/ABlvWUK6gVvyAD26wJLq0zIxYysu9JXl9pKj
//wGNcSmb/Gnd5msMJ8XoNhvLvNi4en2VdPK8xMOeNOYfnyde1wIsk9uNed5t5Uq
97XTUs2/qONflXZ8OKHPb1vqs3xU2WA892vnNLjPIacFA6ujA1yxWU+wi4nSENre
lFuTaV/W+l67P3YMrWe7rw/Itm5QjlYVeMVXDNL3R+DOpBzW//4GzASxo8XF2UxR
zfNBwRm4oSkm0SNga547XnbyGz8ddSKLsieD07wTheO2PHDWk5Rivv6ipKFaMmwd
pHux8e3wOHhdfrxnt+TF0UDj2awbtwyG4/nLHtpQ9o4Wg+mLR7YfmHiWPQrxufIa
6R8XMt+a3VHt8jwGUt1++apaARHw9aBGX8iRi5T3FeN/U+SjgZQ9/Fpsb42Xl11Z
mwvSMkb/FLQ0EwQKlOEOu38LwxV3EunQZfzNnKG0Gxb0zZGdednFUd2H02jUcwZA
NW73NT8N77mivx0rgskfz5jbgu6HPnVDM5JedST8+HXbLIWPD7yUH3coeq/tX96Z
/caTJnKTIPBlmFiK3osD3tpGrG79Ny7JABe+04poiHK006jOjB7AdYc6cf8KQSBG
jWEAdXYFVH7Xz2uTgeNsUaY5OyrPlrnqBUH7jpSMPhtlGEopLHYokIEHCOfEMtIJ
V1DbewGeBN9gQJN8sgdFztpSPQL3PtN1qGtnGOdHns6xywXL4wXYB8w6zBONyLSm
c3t+P7RBdjx0vcRGxu5bNZXN9LphRbwTYIAj91+Y2hwLJxZNblxDiOBjTMdLcqOv
6TOIF9xfpOV9Jsb7FJSA4EKrmMBHtSo7Re5iNt84oducDRlnu9bJku1z48cRtbL5
XR0hHgjh1Vv+AmY6HQrIWzASka5e6NYHEn+wFNjxMjwH88iz0UQqDvnVpwIWmyiY
Z3WeEd4/r6bGN2nIH6RYCxKaPLCxoVRzhzGePlkda6qR02nyJQHoWpj2PXD9KX+l
YEgiIQDvPSYrL98b23ncw4qCgTRYgyDrPCoBGUwmqsC+C0EGFSuaG3Erzp5UxlPA
2/Lh2Imklkrr+kUonA/V+EvkEcrQEjVz/A2v9p8jhdgw6y6EJ2nFh8LzRyiag7DV
1oanizf4IZfBr35mI2LdT5/JylByCYqxrUVeNDMntnjUMYetXo8SMOEkFCbDxQeZ
VzWgQJ7fQ5/zkv7ysiwWvXr1ja7dMHsfM27mZN2doEN0nsCXNgOQ9xyuaV1mmSMV
u0o7zolQFjAplrdAwa7eoa62zg9smaU6GBTi0taUt/AWJImduKrQtjD6SRSSqP0u
/AFtN/bmgrefbNljT62Dgn5T1oxb39fEUNpiB5ruMRoAFfAlpYk58PY+UAfCL2a0
vgx0gk2P5pbA9WAOkxs3/IUzhBaNx63o7c02HrrNODwElPRsAFlcwyTb+QTKMpwq
yenc7BdHkd0b9uLJgTX3gOrwiaMagh9QQnQbSCm3Qw/wl5N/7M+2CffRXa83WnH/
3w48kD/IIy1k1gx97D1/vLAIzJ7W7Dx487KX/mDx4zBXZHmlnf0TUVIhMugmO+b7
kZU5sPqFnZSWFl2SaqZtrVI6izOA4GAAo7kIBkiL5aXBzrw7xR/32DK4v+cNaR+i
Kk+wDI5HiF3tBxQ7j/cqHsIPKD/IhqViagZdYkPZ4D7BUXj6aqWrzi3Qc2zMH6Iv
dtUJ9Hbb+fX6BjSTkLY3CSNrgjZE+i6I988J88Tc+ls9HKmJICMXv5Jx/0QDBJiZ
0DU5xsqKRm7Ytq1yvWoO39v3J/n1+mwX418Q2UpRLjFUZvEYmx0bxlB5TAmoBoEm
oPtRMmR9Cduoh3yRmT39BQjtC3DbkEFRhmTUeaWmphaRIrh33fdWD27YYnJ42FIb
OIRVKGtd5jP+XgXwruoPkVSL235Xfjhfl+sdo8DIjdgtWiXgksCfR71eJ9U0pN9I
ZsxLK4WxmbTY3PqYSPa4XEjAUpoP3AZcqopJ3xWAZ3oUgPYjwzBVxhkcMUcUmxwg
KwpasMQObvstyWycVSMwp4TorANmKaKeWTMdCABoj3ZOKDyZy6hy7KwXEXNiZu36
uSEidkt4qGD8FQvJEgLNLS68lGbeZqEhoItCmIIAjI4HIzsFnNvEEyM04FlrYOGn
6hAtpkaktF0pOYTf+lNbiidUJApsNCGqPTVn3atYFk75Pe5WQ4L06m6GHIqddIDS
qc7msvS1OaXtfAuLIq1EJunsKAgnoYuED9FXcUcTmGdwZNVeFvEwqMmV0DywuojF
MJ0ff1ahuVOgo8FT3ZM6z91kK6YwhOjPWUAjJLoZobJRwqhb46IA7FFsle+epa/4
jrxcku27lTXq5ENRgLGyEllyDASvogNl3nj73N/D4kBKhbF17gmKKbQlDsU3Yw/s
4BLDqXXliHKEaNMTBwy3ad+1eo7YvCKuv50VpDnkNnxW0mSk7m/u1mWU2zbAF5Kb
ehfLFPsu82iHXLbCLJ96n2A8/gij76VcYgWm8wVkUoeiKXYy5NTrR7qqrJxs9koA
nwktKVy8mP3PIGY3XQP/xzAkEToq09W+laM884QQCs42lRq30Jz0N9752Xp3wyDb
HWRFKZqIPGX8frWNmKo+bitQiLBXyc1L7g9+oeGHnfZzNcaiWVo8xZjRjYeQPGAe
LvCYKf902HUDLrzeUWAGjJti2oC6vEUU2+si6aCQ2BlVOZvi+GvIYVtOOBDT8jD4
S1NnpFiSxZmSjxd5FK9fnB5eyerQV5LCWnH4s/TuYoFFo8hiLEYaFb6TKcYtQNWp
03qDHvpUvkuc2cjErQGok3/QlE2CSpRf4FZ/4OSFc0KGOBhCVx37jTX24ZEi9nmy
TUvndXEu6GFsN0e3lJJFrrEinC3zS6khW6+b4A6NupTsjTeUlQd9YNV8xjHKuybB
1DcSwbsL0tBXa6U81BnBupetzGrPITEJaNPydOkdvJe0WBDruW7D18CXc/9cGM7N
AxXcAJpK0mbzXNEMnoWpqJnFL1pcSbll7ulrDkX5pTZGx+WpLhR6x39mZ2bbNaGD
eEE2xky/VmH/xwNiNp+bFd39TIqTQRI5c4aEPGnBCWQ8QzFPxB+viB+fVkTchU6A
qE2pQm20KIZUieFugh3TFCWG/YvBiPaTM7jyj5sMVTSugdAq/oXkPRY0UE3KEaxJ
iBHBAOOisq8uD7Xh1AmLoIpTRjLJSqj6fQYK1BXM1Coc2La/+BRnNlSM2Tl3xOuL
boLw9LsLiZ7rN/Fzywg3AfWAQEUOVmmYwwaC6MzbqY8gTtPZQKwFn1mZPXdaENqP
mJzEle5FpGDSXtPAgRllBJH/c1N30MvSybQQzn3kgDe5FwkkFnrcgwA0zNLO99tO
pJ3g/fkpKJD1NsH0DHuFRFvYl7IYD7FSInJVFIlBMwO/AawMVLb97R+7qyttDkZe
3Y3/5a0vdv8qoPTC3Yw4uxuD4c6q/YRTLuPmw4XC5Fj21UbBLdgtiI4LLy8p+ss+
VeTc/cVpY8GoNOejirrdwR+U9Nl5SuiJtrF8nuBFNXcNn3zYpLj3ixfCzu24q4sz
4myaoJmQvaabixHpa8k2IVxZW0xj3g0nbPfDvXR08zbM2Yg6QD5hHI26Wtz9ehoq
Cs7y0v8UG77AmxCvIIMMuKkvJw4othMTHho9A6V50hjNq55UxKO64tzg9PasN4DX
lxLmiHJpTCf9eXd7faGrNrd5T7tJ8fnS/ENgGQQft5SNv8vsOuJe/yqcpE4KvkE9
70rCF7iEtdWkALV74XtpHEK6l2WHXh0Ff5ICiqHapeSwkZlP9UW+6Z/P+syaxnWk
vr5mGj2HozmIEoQNLCK3jaYT6sY0DapvCz7lo31FOT6GNE3m0R82E4WTbGXL0th3
Qz8MnevEsNGTFQBjYQu08ELS4MFiHXt06iGl+jzrRuN7rCjKnk2ZBGvn3PbS/gE4
xwh/IdtkHwiIWmMX8UkEytDGPDQJgwoguZtdNAjS7hnbyGXHl44R/rc9TZd62BFo
Xwu5KyX63b+pVnggdW4R8jWcvsdjNYis72PLy6OOvJihLWVwkwULXc40bm76ux2+
QRQkq5wARwhrr1pt/gWKwtUt/sesFUtTNZvQy/FW6M2J9crihoyfGWYjBKXKa/gc
xYv31XiffcZBBLUKcWqQ8npslTl/KctAluqX6ZteSaQqOjGwRleQqip8rG7SWL8+
HyvEQEqYBDpx06gTRDmJSL0n1CV3/Cqj4HYdiyh+9KcrcXnJjsq33Ula434iFpG6
KDu3ujeJZqzgg4PbAHupg7RHo+32sJ4ZqnXm/X+ENwHOJxeAao5IbNeIqRMZkjIO
Q6dqn3Vwdj6NtjNkIT5WMLQe4OBd+6LRVdiB17R6wZC2hElVtHqLzE8JEbT8Hb4t
h30pSZHjcRASN4wnsFbWxNcy7b3s/EmEHgjF8bk8OiXA+h4b6IbEgig1h3bM5APl
srO4bAdUzGUAZpmSTJKimmmXI1Y3mpslrz62PHPj62xhCaLP29txS9RytxXFGNOT
r8Z33Eu9BWQNGQsMKsosbImNy7i/F/bpieZU1nmRBn+VMnoExoyl0tG2kxjj7lAe
B7JJkgXbRikIpc2pBvQIbANOv4CCmLR28tDQN5qDDRffNOCTVHPObM6ShgbsEYLo
sPjw+Ap57wRS20qXeBLSPhxuG02NYhRT8gAWLgGXMM6RuQGWbttwmV1qSskZcwfF
AAmcqQJGkkSsRlbzLIfKQANIKn0oVL1qwlZjVFZHshPT1bn/EFhnbLst+4UjJ3n7
IdceWtpzCZo5Nh0/BdMlzS9fChFnWzWag2GIzBAwfAhOaYqtIee5qOV2PzAU1tMu
0/s8dBsNhyWYltvq4XcgDAoDif5JbktdjJ1tji0oonKXBzv3ManU1FNWYPtFWtDY
Cb8gT6NGnEtwANlojroc8iJ54xMyM6oZpaxKjYxqW0+Rdiij2rECXET+e0fTRO5D
zml0py0bv8vDHpejkCxXbPGo49opE327+FS23kNIl7jnvhaEMMkRUUAtcHokd1Wo
S5tyV5H9BWm4oVa0kQjGKmHBEwU8wT+Flv7SsgWsCMHMcrHV+at9XCpoIfFzxMNs
0TNWjrAt1cGU+d6guFJCMag8MiFgLSUxbCAEFvA9i/q/JDzaOm6o7I8fHpKUAiO4
CNx3pGubzcUHLwWdMdFQZHLzK5kVYQqrrtQJoDDa7NJpizfH0GOBH/efJlbQhlMD
Rfdkr+0OldifAO3GaLrCY/eA7t/twtf5jJZl44qd1vNdLmOlgg1Nv6ZZCFxd1Uvd
GAkeBggTKORBFsnFmHeB5212crUU5Fvl6YuWaOdWWOnTXKUrdE1gxZHjIJYmFJv6
HVsx6zKI36fUh1YzNlqLi+IiupvhxvpziymqaCVA0EunhTkIKXSzq7kwN1tb7oVq
xzvGI90HBCQyJOcgiJYI+PvaPAM/Ks1A9mVBT090OL55XjHyapNV5fxoH97HZzOT
PIM4DJgvs++Wa4vmBkol4nqNl5DOeNK93qFD9+BRrXlOsz6YRrtimYKeDQcz3cHQ
NEwq9qJkCEI3qOXQBzC5eYv9xl0eBlh6ALsCQ77a0zq6PEl0r/cT/IIAp1N99kfK
3ZJ3dsAN9Iqu9U1eGwyxAUkwLYGcuF8uEqpJwDE5fxyjYX7QDdmkF0IHuEeuBy/g
ymhpAPrLiNjyHPcpA1evI5hR7/sEU+Yejpx0GkdwOHE4uXRDC82b9l0w8mh7LVLI
vEq7spln/8+umHuth1z6qhKw2JE/kv5xV6FC1OExG47IlzclxjE3Q9riBrHqWmWf
iWrJhF2qg/rAyGmAgQGDxCU0NKiXW6hMTzwDTUr3Q2LDV43nO0ve/8/yfPhsZnub
w0eUqQGfVFtslvkD3JrBjnMaKngS5+3oZrv0Zyhj1VnPSwtjTNowXqMN7X/HL6I7
bSIddzwXyO8Ef+qgt9Q/dp00lAg0VC0Cu3f9cWaUD7R/FSPElzZicQ9LjGj9hneH
Hut6/861fFDdHWxsCalUjnbLyPHxLy8jTZxvRgBzKykNkXd34y1lm8Deg39SM7lt
bm/hMgiDp2pvL0SeWXx8p0+c229OEyRvEJVJ3KkhxWeeLk+xeDeaycNgZ1M8qZ5K
gJSryJ0OoRua95LiYrnD/EH7NdzJYq+p68W8V9RHmyzeDkVtMUsx4YoJIgEs2Zdn
BDfT1uCcMGiD0J7lvO8N2nb//0pM/zdoyHMtZLYpuXtICarYYY9pPAejb8rVUVKG
SXD+GeRnB6c1VvWonYqQbaUGqXnbvSL78LCuJ2ZenZ8SC/myDfer+dNt1O0FWMBZ
8vBgqeWMd2ZxcmQcaVJYrFYGmP0/hw4EXAFlOPbdaqv96OqpqQAy+vkX4uPyo/I7
GjylY++Q/Uu1VTYtyCvOJPBtShljoeqZaRFJh72i1K0ktGC3/8n+y/Lii+OY5rz1
/5oKq7MYvcHt+mmPiHHfap4ibwoqZNOw/aPgY3RdBH0q10BZOvtZwWJOmoNZA+CS
VL995AL7T4ubu0gx+6Z0xZWxnmgPZz8E8wo3q9b2eI8zH0wzn0jG3nRGL4xmpUe6
t0XeJZriA1W8GOE2UAG0qTPnkFWEFeYfXzEt8leGBH3ofdoDYe3O6XRP3Wr5kphI
A/mUgDk06KUzJ9MbZ/ESObQV28dG4m4UDb0gPJ2wrrJXlwBPJansRjPRmc0anulD
f4jqESqxT0OVMJuJd7KlBqUXvGYu00YmzTHn34rdvzM+jqu4bPeQ5LrpPUc6XRN6
4uhKriSzsFiMS0XqDjUgmcNKeIcQmO9uHju7hOLHq6GphU7fzH9CNtdcsXXwwNBo
Kg2jcJ53IWuiUGFxZjG8gdxvJoZQeWEY8VcyO1QZz2meeOqtEJoLbDdjtAkGBNFt
F1+hhn8kAY07PRHIujAmgzvKQ02LcseT3Pfz+3HluE3R89nT59ugyJUWzRqaQZj3
TfcDKiNZcLB7LNivrRC50maz7dDjvO8i3H/Xwu11g69ELD4L3Uq+OVBXB4Brx8zX
4wftJoargsMf8ihvrXS8mdqnVO4uNBkx3AJdJpgBDdEGuZfQ9WufGTeZ3nWOllhI
KaWTaMgPiFBBLYYe3Z1kdgVNOY9h8PugotFfT4RA8eOiOD0pJ7TunlGpcsCgOfoQ
0sh961336N29+ONk7kVUHiaR9eJaPOnP9tVdmjEltDZG9WSVrndqYbegAQmCp6Wx
I+ActAEgpGNZRx4Dreu2xPdxYrS2CtmI0me5LM9apS9GQvQK5kF6rddSLi0SLtD0
iBPGNhxgcJaWVL0mw4ypXAgbjr38nNbx9rCzPfR/+/+fI5KdHkc8ECeNSbNAeEQ7
8KGikhj/0NIObbGWN0GRjieDENZActGKC7P/j88zTEhMJ/wGBulOqSUR3BnMMMPz
CQfsugLJ+CIaR3+8HsCL3CHuLdF4RU/krbTtfnJ1QaPecOF8ln+DTi5qd/s2UkAE
VAoR5gGweaKkLnHGRpMVqnaRgL7wte6E81cdc9aE6+9zyxa1iMpVrClerAT5w6Ly
4oc0wesuusPv8r3BYY96UPqJ7a0NpWi3K0d0LTOeebQ/hiQzckrcGa7EofYvBk42
hddN5MuNic5o2MOagx2JypfozbMNIEVgbRLVUapMmj6SUuh3p09+d78kvpqexN3q
zwbI8LZCG1CdMKmbVkqd1ufvIWyJZSwn3/VFsuzxoWeCp26okfFkUKCfd9CzZ7Wn
5m/YxoSFhwDD4LbcQfwrBwuw0VHwY+2qtxSBE/fvE6MZ54vVDPmTS9+5HWZWkY8r
AB5f/Fzji+4g5Noi26rhrP+w/EeXiK82AfpuhGbKn++vgSdjLF0GhcCg2vjtlZ8c
eIWYMJ9ZCSl6EmFo6NfnBHAjXd6HPZqFW/usCLSWAmW8CXtfhHyfe1xTcpZkA+La
NGcI7K9B7+8e4PA8Ym3+hjtvNCEWwqZ4MOkDHczATtLfoNWDogxoZJZJxaquZ/VB
M/pk3sI9ddgeDM7FfqBgHpqXLRyPSagwP4E7eVy/DMM2Ax8GIW1DrpfRVeq3/rs7
z21R6UQOB8KHolns/Q7Whrp0yAjWCtnA2FIhGXll1FLgsVe2FrOhHdJY7Cf+VooY
ERxvkqFumMPk/PqP5C3UOlY5PaDTm4LU244N1zr+RD/ieRJkqXMqAjAtalWZ4uIf
Lu/JR3UNGz7rgz49DF2pePJTosmVWDkLMfaMwwJiJayj2wLbUIoXQrNB+eD/orpG
fQ7GtqVl4fj7wbTe38clY+njldBXH/1WKbkz5sgkFWwzqKGqSfJqT1Lv9DrvAGCT
ad9YuN6HRbCCarpoLz0t10yCEjhckoy2nASwsYTYYzEw0Ff5ZFF7O0566jqv+RsE
4/5ySe8yloQU0iISVlMo6Bx7SpFKObI/UNpmOxm5B+A5V+fuybDEwXHszizEDRRa
O7ehVtu8SMQc3ORQ3EDIyIJXf6g6BFuNkpUz6m6NMGtIU31kiggDtt/Zz83LTWLB
Ah2X2Fl9Xkw1LXr6bNAxX+EIa+Rf/MgaY3RJnrI+56pA54MFdB6xf6XVg56DkCud
NkJ5gdQXO70uREJ7vgSaUwIdp+Cfnsz46YjbFgGcrBESvrf/qVdVGGX4OLZslZ5n
Lbgm8zU6CZT/IVgB3GB42MY82Oj8w4wSAS9pM1m/yrFZmHylc+37ZKLrOrOpXp59
g0q8rZo0yt5OweKlta7Tr0JJ3BhnE36YYTVWWqj8A69+3DjsTe6+Y91JpSbyWui8
8LcBYHBaP9vjzwDSg2cPMmqVdWaMm8qjZxP2UUoU4xi6qJqREVfHpZdTN6dVJEGe
dmcWn+xfmXZ46aTc4oJwQQnyUIpEmtWLLlI2j/GNmVN6MzPIupMdRG1yA7j0j5G0
rPuWmjXt6ZWsWzrWuX5whep1gJ/ZnnkFzrmDetZVE5iz+aK/+VjS2ftMp/zQobu4
170MRz6c2gTKdKzLKxoz/Idr5mHjQTlF+JkPNH6e6i4jeX/6xQdjVKb1sE1g4pcU
TPOXW9eRSHKzFpQ8W/1cn+cK/7OWzDy+bq66Y/OscyhaILFEswk2mhSNVXby4FFB
ks11ZfF2KgY3uitA2B75xaYMMGHHOax/pQP0FQKoDTo7oF3QtxxEaY9AyhpYFmjY
n8AdwAhN3dlCoY5HjuRbLpuODebXs2BdGsOqh+NQMvUUCAgW3Y/MmZ7zWkHtUY6e
yZ1Hh56JXBJkZ3Ur9xtdsUJJpi09h/s+C3mKAWcAHdHR3CnZkix51nMIZOZmf7NW
AYJJMAWHXm3w+EFxYUJfRcmZ2s43Pd2WN4ce4brRmVvjNgWLLqmQOveDuAHTFHdE
IRL3XPD9ylcZt7odFRXGIVql8sEP8no8UbSVibfXunH8jPbnZLX0jAetpUp/FrDZ
LhFAekTRM4HiW1bbyVAbiPwXb/pe0rftAsCqW9ck/ij96Q4a5QB8lyh0AWtQSAzF
AIcMPjZ1tQmbwJpznkeYHaFbBe+iYR4iXpzlQ8WN+1psQdm9Q9joZY1NV7WVOY4G
UyTKNrA/zNG4FMfcr3qXbb0Ne21W1Enxip6fcA+qmtqtts9cRUq6fPst0EEMFWQR
H+PpD8Ft0FRq1f4Jsa0gmM+g4TX9TQrUUxvxYpBpC9okKp18mgLvaDB4hrSDDIyM
hzYc7dxhbkgwCvNz26LUT6y17eW5e3QuqQhsR9y/LqtETdeseZwsRRPkBRzcxxTy
4E2zRqSD450f/s/kpxSAGbOGGmzgxZybrHmBg8bDG2t3JTLClH6eHGA23gHx6Qh+
hLqAa7UMiwheZRKmKhWdS9i/Il20viN1kDg0lCbNZ0cqxaDwwwDTfQPAtLKmlD2j
vMqcB0W0MK+vKzpJgmJN1sfUY8ha9ArXEyV2F9KPtUGMIeRhpXOt72ef/I4cVG6e
3loOKuUAOfi2gbeGYnJa09pDywMTMhG/8YnhUiEx+n79tCiL8/jnvBlV/AVNvZ4h
qZhX+38F08WVipiThYSviWMDyCczswgXz9cr7dgGcj8LqNAGlwZALQaenLt+/6EQ
nVWVS4dGgUyEqa5e/8NsLFTWocLDjbBFMQEkdD2g3PQtWDM+0or7UeIe8JCjVTLG
8z+WJeK5X26DQZ1Y79CThT5Gcmm9BzG2QsmMQib2jB8yBbzfD2llkRs7/2r+ZI/0
GFPJyMc4O8PmssHCUv3S7b5RjqIEh0pnnmfYIqkQEoPTz9oIwZ1iUvKA+U/A1P4F
tfhP+0vWqbzyM3VDcSOWp6iC8f74/oklrzhTadjxMvdygqts/VZB12l0F2ch8sCu
thSn+qy4CAzbCMml5k4jo3/BS89++vYVG1neQGpM7chKHVgmCdNQVMmaGAwaUMKL
fbLlOjeIzulI+Y9AAo2NOp710C9kRrVC9y766TbESJJw1VwklQQEByhWix3NZoz9
3bq33VteFVdNtniUi/MNlWNrxJ2sxNI9TZttgrDVx5rdrYKe0vDUgReGSauYQtRb
xq1qPc2DRMHoOiORfwPqjsyp2csER1F4GTwoCpfJGko84TSRgs0CtXg2WxncesmW
cWezEt35L7CqZTq3V5JSlO9NUAhlPDlVQwRV9KbMLd1kUGuvLUteEt1nL3vYSkNg
sW8Z1XkzbbhyKGTtXwiAKrr7pFWryAK2hoWz1fLj5TRzGx9F6MOkcx3TfCO+Ygvh
Yas+Wle7HeTiCz8PO70MB7AKC0LK3PR3cuxx73WM3rHmEiRBsjRvXI5f3s5aHINM
KZ5lgY6Z6yj0uEQN4OHo+UgXDhc8JV7lERy8HYYBGgO3dzym73ubvx2G4jAwWgAh
cRCFVZ4h+Cgg2pRh1I9CrDIUogi6w/ahfpaVaqTLnstUjltCySld9MMG5lYf3QBJ
rnSrqanwULGTC+hGIy7K/pzMi3UfSvPC0SsNhXDN8orfqR5qRryzq2vjOIbmwp2H
IZDg7hhu04RdeM00w9UVjINxInKn0h7zBECK6cwcJfzUyCMCA8ZZhNTNCF+uGgvn
pELjyUrEy1BOK22iUvER9OnWziFS76OQLdYgQuG5wjvG5B2iilBFrBQCbUtZNBCH
phWq99HFC3NK07u0hIjcvYNpESYAVRVhZcCiQEgRgGH+MBNpxjM+kwvQ2f58itra
DI6JmVHT4v2l8bQqfc3b6Rk7eHENS6z1MeLnCoR2EtBnEEtfUoMJ4b6v/V9q1+eb
yvtpjWAwMdD3qi2IAcbrKGL6j2NDGKzQMfD3yGxGy1Q2ci7z0HDM6Ss8uSn+eIB6
nZrf+/B4K01IscHIbSqvhGQV7fyr6GxwTgHuo1w1wOssEvPkHsJFr9n4fICQvr4p
imgdy7uh4TlhFjUjbjJC3kIy5n4DMIZ4u320lVlReWCqRbj0iyTC9+RNYgEThQws
M+arLhZi3yZqfh1orQ+/wzAf0vHiOss7y8EVOPHBF6zfEippFXJIQpaOPS9ofq5x
l4KVjE96mr2NY94+r/E18J4eQv3Dm2JbuwgSuU7xTlcT3h1xbG+LWWyhkFnScRJW
Zwtq1eNMYbLVQ2i/9wBjgYgQsrNlTXJHU6/zQbBf5DwdSeR4dXgwbQQIwg0ttAYP
oP+i146kmXrEjHCjedIZHQg7u2Ijc+y3eWcQ2EZ4wYt0jtP5yOOcjlcncQweKBvf
J82THEtlqwuBhg1ubFZNAsrI44va7EaWLmziqyjzfLmJomI9DkKwFB//jR3Cws1b
wBjazU+cYdfYn9OQKbzsNSPGmwBxR6z30j/Z3RxBfK98lt0H76R2zqQR4ClRkVQV
Yq8YpYIw6w24mw2kCOFnFRk8MZm8FzXKcy2qJ6zjm1v9HUKSmCgZVlJxaxyGSepl
aifb/GeyRiye9ohAVlqHfOT9V03R5aoHN38Q++xOaoK8inlHtUMWvMeBrEM5eNrE
Z6cCop9FpLxeIv7/ofwQNtr/fBSXoolcvV62KJrsqADWcG5mGeGdebgcqOlldNhS
d7stXCUXj4qMxP/YpBuzoBVTBgYPILueIRO0nPSn1MIN+CW++NOIcvi+xGvYldxu
4Lh9aejhwD83UX5gQNe35U2BMIrTaUJGKNhWBPNKrd15e1mMVSAqGm/wq73pDv/8
0nSvltAx+EvimP0MPHD8PZfK0rSbVP1xj7WGHf4KCGEdh4158HHIZ0WrYyHP/FF7
oFwqiFJ1JoniAyuVvk02WPYoq+JAZY+Odj9ifjaPAWfeEOvT/H68XmkLqk23uK2z
ZB6v4nxSTXcO6yfnhifNaqJwWeHR2bNWQPt43x8Jk1VIQSbQFm1uyUVpaog70QYI
NZ1zxUW0VVSqMTdcATNynuClNrnn7XpgmBO7Y0DqnvSDNjSr67zjM3+mtPeroULV
zgvqHRHtFS71cETJpRDJwa5zLgn7bBr/T+btlm1RUuZsDGGpbQYdQZPJrsBcugVE
BHPLcDCpk9MfkiABPrp1il/SWQyn54SYajq2dLS1bxajA+gSIHllxlmdDXdC2GVA
VUYp1fu0kkF+vxK5yybV97nxB8sNGKXQHhQKHbIFE9SEhevgdTa7Dhi+sUYg8BTd
XYXxm0Lqwr8ifKGnv2pGzJjCm8ampd7qdj68aUXv6EWTPmoXaTueImqeqqiA67xb
5gQAUoS1V4b7lGbPf5iY/bw0ACB26OsyiGhnqlsL52ozyvPLju7B8OxA4A32u6Zi
vojAu8wA7FLuPKyQwaNhWHyIG0MNApcBihWR+PNQLuSW5+5KhKyfdJMUSkJYdinb
4758qNUBuncia4YWP7lbLgaIGBJW3UpHxvhiVhCM+bksCfYEGJLcPTDgM8NpceZS
//16I3P27bz5EoXoXhd/xBdKLkkmLcALYyeNmh0unHlu93hU/CbQtLA53Aixc6VW
f9MLtoeA8d1O1dzLRcRx0tw8ZnxluaAwb4pzCFYMeJziZBp89scMryVu0ykoz8t/
diB7kfVgzihRPukD3WN9O5/rNQSeKtwCXL2CzL1Fi/vCL3Tzm2+LBfemWd8cyHew
VXniGVxbFwA8sXMliUZjHBHsg3XPjJqjLXA49DcMrQYEF07Rb/o0gS/Ojeq3T/sP
TdifoyZ/QLQRoXqrBFLnZ1y1RtviPtQ5Cd696ix1yEbX1X35aAkQJbbjutp3IPlS
5U8H4Mg8CODJsVmxJz1bglM0pMumDn+D7vNzYs7bJLM2F/shgxIxR2sONPWBYoQ6
f4iMM4KHZ2TXnggppc99stzig4mRs+jLpcRFg/vbC5MipmqkozvBcvIuFDfpcWHv
10Nhk4RlG1u1ALeFsLPOciGSfkeOPSB2yQQZmu07LR1RvcD1ed8IwO4LPNyozlJM
bEPwxAPIl+n90yvEh7xnu58JgLcssymcksgggNsu0v1C9SJ9Bkmew+Clze3ld/Q3
3chi9CHc/9e+onQkMsvMvdzp/KSGoTMocYP1UtHyygHcmfQt4b7it0Mxo+abyk1b
e/Ys0ONNnqpwo+ScbilFiccQNCKTeEQyfr3zvaxmSWMuAxa+ubK0HtT5ve4kkQAn
2hjhEt30lw6grChlfX4NT1koXwr1jgcAed3X7k6/bBdYhO7xOeOBcJvYEVOz+q8v
+sIHHU0BnzQJDwtd/KyBzLgLuT4e/o3jy6jaFFsI/BVB5fOkgH/4wVCVIJ3L8Qem
UcvaZtkQMD1LYaY4/1BWx5Yz8qxFOhThRNpomNM4tCJ/phxmOA5kBH4yotFvQIJO
VgmUSVYM1a55XgtIcQvXyiNVhMOBO6a7B/WvYlLp6On+1Vpl47G3wLGobOnNOqHJ
jyeFq/FW35jUUXeZQlkE2Qbx9oH7vDpGi41Zk9JuflVpWnh+S6Io8MaUQoS2g3E5
A1jdnyvSkRVtVe96XGf7frqxskz3xUcZqPtKs1i6KqecnJtUfYr/8vJkJH1HaLn9
0M+cD33M1UvQhDZZZUKH4TsuNdNDcymuTXL1zhmpHHheqXoluPMfFSc/sAfoQ8Qb
RiiM3QTVje7Xujn2YAFfv+BILCcwNmhM9PTtlJqMZE5l9uDU8pseT1MGR12bx0IF
4ox8mc3Lxadozk29Txh4B2eKH1S7H/ywIsUfUciMzgtJSAJzi0810Nm1Lw1KwqzA
539j881PHo60PdCS+dNYggGvHY6MhxhdmifNfiA8KrjUk6UeEamjcLV0jvOhiAIm
7ic3yQavGRlhZIn9SMMGCnzRUPF1ro/vk2BspVRcx2dFlgh6Xl/oLaKZgEG+4Nwo
BNw4JiZUQyv6EW+22kBzsZ6BTjC6gFWB8DLLfzX+TWtyYfeOaSiA5CWqVyaqF3fR
Qk8t2arVVTeNeL1KNiViY3v4wxn6jV9qfHUaRX5j7FUy2Qbd0uGUN8dIveQNVRP6
0fz6X9jBluECNsOq8BfDyKDODpXb2e9jUOQVgQpBb3mNT0mN2LF2IHb6iDVl/GCS
FzdBlcS8Q44uuf+iM18oh4bUB9vAhs+INokykOAnfgT7CiUPWxCOAz/IV4slQDnX
UnMq1R4mBzpxAl3hOW3wrHibJAnO7o625zUW4GvyOzlLLADFUlPfRNbQA+3MGurg
6T+ZCgecBMVJdAGa8+7fok060roUU1ydQJ4DhagCocn6wOSUJj5mD4ZAbVg5IsZW
UH3Ksv2i5v37ylxgcM06BqeI16mIxRdD/LEJIwKyTpu/7MEvChsURiJiNE2n+CDa
N1o2vWHQML5GTkQQYZpkUtBUGK9QAgw3PxYFZiROJbZSvip+Oq/EZ3FRfL+kpboh
RLy6tdI1MGLIWQGdJkxAcsM4qKT/sK4grt2Sfc1HTvbCaOClk6dznBO1VXn22U0Y
Wor0Ud4m2cokQRkpBnS0O6pOEi65U2DGaAH5JNOqd32NwPDXS8tJOK5vj6LF9L9c
O2ejEquIIMQ/I6QOijMqJRH8eRbj0NfdlTq044zxsOUkhizokmrzq+Bt26kD714d
GdskryAEixIDVavERWrpQczx+f27RDyTEp+9069tuoI2RDYPFKhIPZWKSLk6XVh5
jyPHZJRQn43YzNk3c15CmPGaJ3yX68Cr9JDffJJv4FzyTtN/Ev3qAEldwqC629fp
6JDI38FFybomN+0piQYStlCyjF2Io5ehush3Dxaf74HRE2d4UKO4ycwZVk6RW2lX
HTf7MeylZr3BTj4aMA45zWeLHpMKUvI/zsWEC1PgorpGzGvYXkc62YKAtNmB2qvi
jVGZ5nRfKb0ZJ4tZOqQoQe1o4Aj2lBYSvrh+plEUINpu7Foz7qkWpa+WsOVEW6O7
jPNCnUD4nYh0WDbQSgQSAenXYY0QfmB73oVP7ynCBrPgRbbnTWUtcBOAXaBL4WLL
uoNknV9hqJgGXksJ7eN7moYC92iuKjCCAl1NjddXB7P3/m1kGwEObsHocN+C/8wl
xemIFdvsXgsWTloY4NA+9saS7RXkgZX2ic6dqpgHS/2B09XwqGWXZnpI5QaWPeWP
8t0E8Bg4QA2GspCWC48DmDIkMdstPyktHrmM5YBtrX1MKChg4U367ACLFcN8SOgq
BKTkK4K04drvUBubzH03N3UI99naIe8Alof2Rxm4SHvMINz8ZPJ6ckik2X1kSy/M
0vy5I8LsQAbrjrXfGPtlsV8xRjb8qUI1onZZzRpyRLF4ZXghIS/9CT+aHU8zqE1H
Wgh/eR0g2YaNT7GwnwkpRbFaxm4bvkLYV/FHw71b49QxZohdaQU+nAodFjy2PVlV
d6/0puhhmgVk9vQ6MvLhdyIVIII6wdnA0M5YcQS8YxaXE8ZSQNGthXTTzpukLqq8
Dj0rZL9uZh9g7t37Zzr+CZkdgzj76N64hMUT6pueat96cTSo8TzVXSt/ScWAraMG
yaWcPClKTDAIig9zb9ZIW+sKgmq3bc6voLNA++Rm9t4Xr6rQEbLoH0urdyiXbDi6
3LS514MwiT3JkT6dKkEAhnlx+pKiKPbHEXUI3GGbwDHceaNNwp3oXDQHhx9yoxBS
q3Q3qlDCSzZJKVh2pqXc3W8WmoyapOOqLBCpuQ+oiKM8qxmTggIFMQ7FnHObMKY7
Q1hyMLfsqPk9sJCxUtlFRvMLPwkFYZz8fr8Ol+UJPrHHXBYujL2xx7cO6U21jbjE
BRR0Nt29whDVAfEjNuf5pwFwFLxlYfWl3/2v101QGLeVE0aoZy7eioaEmhi/jUnJ
0oA91ptWz3EIWFzPHT0+rIX2ADE84ZjkuiUBKXM2KMZBFUYVNfpljd/MYSYxsGXl
5TQzmMehgZG0VmsWMKFGJtuGjQY1swMUrhQNvOijueEjdGmSlA7duP3M1zmgR8JN
WSRgUS7SBBOLtq91L7uNMzxoH/+mskhQGX5AjE4s+vZQkMGfOvuNGIMfmYb2Zslk
ZWB+FODv13wVqyT1NTwZUj7kYq2cNMc+NPOaMhrHT2FyFdm5cTz59J2umqNBxJpk
x5h3umxa3Ov0j4k1s7Uw5y6KsSsrWCFd9Ob3TMjIyGSnY2AhK+TdsLgOSIdjrXME
z5mI3HnF6AkgP9SpjsKCdyAgQbj0m/7mRdh/fRaDalcHg6RwrAilDu+X/emGQ8z7
IQxVGvBXo/5h254bHIzjizjI7nHb8m/fwbtNRJSoB03IFQl2XSMFKlQRPA4rhvIC
iyD4DI6JKRh7GgbiaMqpnRvy9/Hj+RO05veqTkMVvh9V7L+TCc6JIcxjlsaZoiZa
pMyo9zAfjEAcwstUCi4plDkLifjbDmDrjaWHIbDZ55/UdKwmCuUc+Cxl6uZMCkeq
jP0bu3bMsFKDdk3EU8DxEACpwnS7+Alk05ZS01eipAQ+Be/wBOZMQJ+UBz3jxLz0
Sa5ZnqfjI1HSBxFQrhFDTTR7RWUOYOLOhCIX+o075RiUgsmDo//iHc0iivK78wZf
oGaQPhfW8Bn2+N5oWethKVIAQJMYW4w1t90qhUvs7xyw82WiefvIIV1u4aY2urBE
1GlCM3yU5rGEei6kouSeaKXEDzUVlQoe2fhpHqbKY032o48o0lzRiRXOBbdH3oi+
2tJ5yn/gTYenyIg25VlaoRCAZnJWyHdWKU/EoeayE0V0/Aoq8RCfEtcp3rZZGwEh
wXuXOLq+O41nlB/EUIY/2oOBLDc6XLy2SCQ5f3JuqjT0IMv4CyAIj7i/7d7WTrnE
U/f+HTApzOAm9FD+BqvnX8EbTVvYbwZO95LK/XQkzf80B8k8eKwFc1mqPFF1yNT+
YS7xIS5ODtYJfFrg+HHbiXa5JnSBnz0pcaTGJfxjKxkesGL8cC2cLzv4Dwl3FcBy
TPWbLhr+8zyFFwJFxiMASkfLNOBY716W2V8bHeVC8w19NeMhBWwDJGqaJonxcX+i
UR3ir2Ql7fO975ouIhu2Wj5eyGStv60feGE2aigf7nRZeOQiP4V02Te+2lg56Gtp
fbK4oQfL0IxqZkwBEk7HxZfUJD7tjZBp8s9nL/HI/nF9qoDE6AgEmdwTIl7pKC2m
ELzYbRwvj/soE2y+29C1JdutZO7qBSGnl6ZrexYshwkV9wxhm49km2FxH/MVAafx
Nj5OIyuZa87AoZlgz0/7NkOofgbhtRnFrnx9uvs5YvluoSm7TBGvlVp34tASnvRn
GEqIFlagR8COODWRrArJxZpj0975z7fvfz2tZSpcimoVY7dwgns6NgSnrM7ouhW1
yXxvxWAPNoDhY6PzUxANPxV6f5wOQgA8It8gSQyLk8buNd5+X7zspZ0PnS4DvUii
Ld47w3rE2msjuF6xbm/ep0R8y7SyyXTvOw7D0VcUVLW1I7UIMB6eTa28AkIOBM1y
UZL7Rag4DLKMvoOHMO4b/RRuuvemswMqkgQwKZ/XNuDBJ7L0f23IbXxL7CEks7eJ
sqQRVn/ocB9ccry4cRQzLmenLwLWi9ku6+8weJLe4W/jukRgQ8SZyJ14pKMaFqug
3eYf/4tdlZX6kXMOBwt5S1Bli4aVWtFTHdQF6OvJFPoPss1D/c+3rcMA4bnB+YBR
r5ImBvtgzvGCg15vvDtp2FBiJuUpp7/rvWEbEjYQP0QkMdhX1B8186Veh6TB4u14
V1b3Tb88iE+A0gaGdPsP/dw8Ugs90JMspuscFeMl7zX79R0cJ3Lgone9pjuW6mWD
4f/AKUygcNE04HHECntrQvuSHZ6Gce8Cjds5FVzwUliWjW8gyJrc4DguOY1od5on
x5w0S2/E1Lgcz2mt35JEW0Y2Agda+NWRn2QvjTbdo4EWdsjy8QmVb3taDeeajPbi
ipkbwTheMdVigQWQyIt6K26APpn+mAxKBRR1cAGXP+KEG7yHaXVemwpyLhN9B4ZQ
2KljlchElDDWDLHf8N97uq+4yLqCJC7f4CqdE13QoImND4zXOX+bmI7XJRlq8Jjy
Z8QmXqaRbDxQIr1kzbWgMHLaD+RXprlzM2yQzp1RgxKyH2JLu++vooNp+tVymILs
L7oBME079qT4XAYBCWXStBtQW2M1yNTS/gD9Wnpn3AitNBEeBm7MYiyi+7woCA3m
RUoLKlIfY5vT6SGi5Wt+mNP7P7JJuESN0Eg6hThXL+C/0a+ic8LvorIPdYAQtmQi
zghrWbyT5iQxE6JM2zdQKB1TGgX9wjpEWjTlpWXsRSkYmMZt3nf5+syptW6jtdm6
aweh5+vdkyRUj5VayHvKY+fViKx4MQYK9G+uOT88/TOW6ySh0RJhBksrYrON+/cn
vykBgqEMDwlK0ZwcDsC+RG8ydIFLh5VnK/lHvDvPTa4k8oSsO29swsf7idLCzsEo
e7jwZ7J8gBgaWxWZM83Ti0h2Q6X8y5MuQyijdRWNVJO8Ulw8f0QGAEMEe22+CXSS
P4RTysnylRMb140LRK28PEHD83bgHjZuLNViz2jvydw7Typ6/dUi5oKUBu2wTEDn
XyD7HQYHk6ANyjUXX+chZEIo9ky1KvDeHpe9jCpvOdFtqSR3KZOs+g3ReAuM6xuc
U3m938qCw5BrSPb439OH+5SL2khe+qhjEaKq0OEVxQ37E1DPgH3mxjXOeV73DlfU
xy9Pxti4UEMvSQz6hPfL72VYgKKVxbt5GLn+U5dOd6dcKNq4M7c7coN1RdaOusv6
7mAABrOVb1WTMx5SsNOPTNebiA91l4/ZiTyr8DA7U+q+diQ3wSmSJzm3Rw2qdlLn
+7i7dvpjlgOENS4C0lcuaYmzRdMUBM70LM2WrGdDNLNFhmA4Tj0MeUqWO9PT/0G6
C13q9CXZ1r4qL0Zb+/MFzEVLIHa96JBCyUn0E8SBCKyMdYK5I5dhpnMbFesEyWJT
D9yMnTPA+ZcugaSpHyer+5LmAVHfba8wtOrLjoEb93qkurSwzTee0wuyH9ft4Xy6
GyZDTcSQZtdM2MMwsFSF+CY9YVAhAA8sHiHz53griTJa43p0785S2VuKnAEOcJTH
scSwz57T8qL4UzvWhlHbkSLJFCWR+wexNt6ou5BkBw7C+A8dO29p+ajGGdbpSKEQ
c7n977d44Q1FVFWC9YfQPDM8CDQAs3HUA0eSMzwlGbr6W21CbRRlxUZzS3LcibSp
EEQO2n7FkuvQaKzFxhBjBUeLoBSj0QlzCliyhIG2EqgtCsJO9mDu+xLSKqzT55BS
1mSm0bCyBL3A1t+7zwj09i9GpQJySSKfKFYwr6ABXvZqAs8ni1PiEXTi+bUE0Bdy
RcV/oFNKEf5V7+HHEhv1iOQCpI9iE70jb/8NIvHKpV5FQubdRkUMAJjabcaA9ouY
sFUx5nox8z0PqvgWjdiexyQaZj46fxIsj0CfA7HIRAMCJBj6jvB+YRYRVCrU3ALO
C4w9dcYG8Xxy80sdVqemG66Mi1y0uaCJDFj8ISckCOAlVuzxuk1/zy826xe1Flac
io7FtwP7Aqj8q21Pw1YWnqVAep8k9Qu8BHRK9SH8eVEGJvmGhWj/5yCFQLBLnVA8
74tTp7xZ2uZpuVqOAhe3ao+yNxzHB4RV7ukT5PsiSJH+F3OCRujkbl2EaesVMHYJ
rNYUrJdSNumgsu7zf2oufi+BTZIcpquouTHHCMVr8DkURmJSt/WLlWUMnYT71MOu
454KfOWv+P7VUQWFF/C7Hxs8YfBorV1rzV/jBctA0I/TTYifISMUrRp5vAbIM8zX
AW7avZyx2fvugC7TmHVLRSKWNt3BfqwtLHfO5QMNHBSrgX3yLt+gzc7mKy8041FS
YFGaO3S4I86pARKCY/mjwOT/AZv2FPJ0aZrwMHL64zIeJ6O8Sl1xcQUoWUSOhgw7
SXrLcRUvFCuKXy1gyzTA8UFK8FAEydjLLWDzpVJwHYB11C2fHTUAHg5z6LemAf/9
cU3T9ffX1YshNgAjbgrN+/duhGIn0U6xQZihjBV1EI/S+5iRpvhYGZVI1xmJ+L75
98uc/zrZnlZgms8+wStR3GNCS/e6kKAXUJmAWzwCcsFbRaflS5Fdmky/tw4xer5W
jgjj12uUWGKkL3nxmmLULbHweijFWnUylPNXKlyRg9uArgADLRsLk/IBFfUlolJU
5rjICWtfxLSvBf/2cAdCm+5N0X/a1e15zPeBHl8TTT64JJtGESMaQ6war7cAqufS
CQ9JG3APoQ2yt0/Of/iUhv1AmmGFMXrKCfr+b59wmuXGQKC/bIOshzXm6tZj1yAX
Pjcvtd3ayL8JkHMyUrOOl6t0kn5LtfEcVjJPWqPbDFkQLppCrwic7X7QwR0Y5qci
/cnlCaXLS+wHyRZPMUW/Uk6hVTOSh5IGMK8ojY1f3Z1Tk2l4xbbW24SuKe3Lr/ya
qm1wszBUpwSyT3W8zZTaWu6O1D4locHRHFc9RJkzMBcazlCi1W3oWI/p3XVoNkzd
u5SDURPHwyWgPinq9kCorhYxs692VtJ/OWHrUuRJrq0KT/OMLhfi35k74Tb6l7bf
bepPz0NsS+ZkVi9bYvWJ5ZKa3sLJZsbH8Htxgv0JJKo4cS3yVSEj7V6MFsd/3abm
xynVj5ufYIOF9dop4lwE24F02g58Yqk98+TCPLNL4ToUY6/gmCG1BQCQKCly6xXw
VcdBq1vziRLJvfbTWT/bEZW3y7QkrYAFEfwoCFgIhvH1mvhNKX6hLiA4e6xSh6ty
P1x2SCmXOoWqgh3M8q5qkwzm9d5wTgAcRGH24iBjLvAN+SBlUHrDZhx+K+SSp7o/
BxcHJjjqRaz68lZ9V8s57+WbcRpFyF7/OTyNEHzS47gZgX3Gq5WG3JKK3LEQWRLP
w+mw4rL9D7VxY5mh3/C00AXRe8M5dkDhlPxgL750nYdGuTZsrise7JxkLlw4Qw3c
6TZN3MSmtpYNVZEE2JBWUc+JMEZzJ7LjcG117cFdFqRkKqDC+dEh0WFjFieroZ87
NNsSyPHaE1EcWyQFUBpij2w2LnlHCZeCC+1wtapzdlr0YyLIubYS9zDIfmo+Gu1X
zRYRMjTlEDBer2PxgV3rVdteRfgB8D6l0eCSZ3wgdYvAJUYIrGuzQnjyUJaW7uQd
9aoLTtijlhxaSF7qV5WuGEDiO+IJ+3wXxxm5iQN9jEgQ7xMg+wYqDB+aQiKZ+7DR
fngUVG6kZlOuEaFDCLw2CJFAFhOW1xFge3j5UnKkiQhTuraQMhng+y3kzZeSqg5N
3XPzUiDSpUOhvYp6Vapm7zMFAKcGrxdC3niGdQXE/m9oJY0FNi6zQGbbX8WgyqY1
srTxvC0J/XvV1XWRg6DrJXXSchD0ipDvmSoMJhj5w4sLcr0ZHUiNmi7Dwqp8067t
/9sQUmACw45UwGZc6eL5x+b/8Sj37LmSIzRRtCpSDJURuZ59+KCrwyouVQ8zBJte
FfHaMlFA5D7ahi9SO50MQ76cdgB9G9zAYJp8MxCl54RqqhCMPbe6AVmWYShCXabQ
0EGGCas224Z/PUQ5bOFcVW8Qoxd9KvILtJ5ZOJAmJFajVSrLaER/NlNeLj/c8lCo
OgHar9587KUb5KyjFL2ZEy81iAtw0LlOkpw7C4ICi0DxPw7y64ATvR75xnPjGKsO
AwP9pJSX509qlJVF8J2VymIg4v/9ZGqKCSQRTY3rgR7OpemSeOqj2BxAey6rZCi8
XoUjZUczfP7pScZ1CvXxwq9cxgkUKgJbwWlNvHMlsoqWy6e3GvuZ2fvAocfnkR74
juKgMOGA286bB8oXhuKMH2CuoEOhjXLcnMH9BVgDGYl9LVSOy50FElTuBDfQV5wi
aM/xd0u1cSCbyVJDEOn41HBS1ghEIiOVZUSSsIYnp9mmB64NxLLHDXsQ37I8UnZh
Bq6WO3XE5Sjpl5ZGvrH0ng475cesU8yQPns8vTQGttX5xEPX2zx6hE/QmdaDSQac
k+CyBCDe203aK2nVoG2gRO+6fVU3T8GIZVNVNrdKXGEGX5g0oGfPnWx3230OMHuR
X31QQWt+x+fI5CbEq2aE+Auvn4dzvZFlEd9OT2qJQpuMv0DLjBf0gzHamU+kj+Tv
eVDVMVpecNWFQ9CtyhWcES2MHgrkeBAYmvQ0eZMiYP86Lu/Z9xOUcOvmhE5xObg6
oQGUhFIoUnllrNoBf61Gl+Riih+whJ/lr5ncW8E3JeJjnhfUWeJ7YSTsbQxBO7aN
5CERB7LsAtwAd2QVj9g2TmMshlsIg1pGM7f1vaac7Y/nOuO0SWRUilFO5A65VnuX
Ianw2QTlJEVoCV4PjbdRN+fvJry8wUcCElaPQRXXtE++s9A8FzMjx1+6qmVF2WoI
nZRcIPmqZdeWNA39iHIYchBCHmfCP2D+d+6lilyidHoKAOeI8OeSKwjZMwqMZ1wO
l+1SR5cYwS8RLyPgtG9wpJdf88IOXb3Mfo9GGqukzEbCLZSufaeOpWR/JUk/JNxD
ZGwFIp+P1qNXLqY5Zu46B25SbnheGnNsUVRnjj1MCnuVThpSLupsH8fAbeiX3gWU
9P7m/4o0fL5+VJQocWY5ifMmthG6SEOrnXuSU6r2xTTNOfZ99LkyuXkoG1GHrmS6
/XMoM0Hx8tBqJozoLXfZwS0pS4l5Rmrg6u3AJL27FsPxvvQ0hCF5BHr5uFKeDDZs
GNQb0aHxeNODqV/YANfGTQPG1FJq/sLH4mJuVqWrimnucIUYvhUR4QHeQVV6+TZ/
UEpx2JfA9R0jp737962rsflsOG4VNDV5BaVCpniDvvic6UQQzYhAuElqXWpKBrVM
H5UAE75q3NITFSYvY4INYnL0sr6nC3BOByBQ83GuxF5+DfTNBr71VhuQbe+0awpR
9pKw1/PLOyk2rUyEGBl7wLYpm7WKs6VB8FWmIe8djq++VdYyUd9T3ztOsabdckoS
Z9Jq6SWsBBABWseJPUnZRnGonjU4DNTjGCvbBMOxoDs1wC7l8rnm/kvLY3AtiNsX
cIo7UMxDdgoFnpUQm36LiJ4syF1ACeKTlgEaSd3l3kk6Dv706FnLrhCulbB6kCL8
PXVVVp4zwupuxxZplChAJjPVxMdR/4AFFmjz/FSSFNxL0gpgZyq8s9I+od728lOz
VIVwIoqXSwOKbtE6ziPesiZwRoOjofXRjQ+dD8S4eg90zif68DOxMP7ltewPJfyQ
Y7NzpWElMTwNE0VGmA9/Pnqpo5EMeKuURRscIggbdxmftLKkdXFWe04oCTC+57yp
wPHhtNiyAERAYWsaRNAdTK3NpiirGReHx+dZPZdoTD1xfoNvzRwzP+CLxVqLUvdZ
niKq4d2V6Jnw3H+aGe6h12vJAHDTo1KbslRChcf9y95/jUkbQlftSPM7WQM59Kth
Lr2PWLmuov0uLYb9+3xU3b7px2NODvwDALgGTBlu4bkRnLHlzxw2Oa3FVerHJE7G
ZD83pQw0LDV/eaWXil7P21h/tLmambpmJwkf3CUAjgRzZ39ZexKDOVtGlA5d6B7j
/wn3xvbdlcgmwA918wjVy9oDQt0uI2xMz7mugwwj5h49+8k1JqrPt4Xv6OsEJUte
APt5ZBxGVPqGQteAzHm1XpLIDjHB1davKMEl0HQRzBk7LWuZQWqQW++CJToNvWV3
ZA6wTIjlBzEyEtk4R2vH96WM33sQ+Dfb4bWIkJrGikqfTIBQGi4Oxv8TOz6tOKuY
r4VcrTvBLoLEV/w4gy6uhosiIdmZc4Z0Y7BFya3joCzZuaxHA4Qur4o7NXqskwoF
aA6Tt+0+VB1IvQC2ptAD3ehbQmg8ZCR2RwYDvg9itBgM7F6nonn78UJSae/UtjXS
E+/bizbTs9Hli8gmZwuBa/wuerDIx4R5d5FwEA8ujcXW2O0Lc+llIMHKRjr8GAFn
TJJYXT7+CIAA2PJL4P+HUpTSCEGJKGNyUb0qcdvHFP2vLKLimVl1TaZ4R9a/0kfm
lsCaUPCurmRYLiZBoSnUHp+lMNP9ileAi8nG2sZ9MBZrinxnOZ5Gu/I8XvE84I5L
X8UErBdvCsAQKoDGZclrf1SCyNNUz/sKvVXlahe7xfq8l0GIsg4/CsCOudsGN6aV
4aWBuWmFueykfOBV8LVcXbZyCOt9hOuh978GHDzoQfnw5p5xl2HJZIDNOALBpAxr
bOqoyD0YBK9KyLAv6lX0uEsxEVLqmjLLEzivQZQOly4qeC9PZLprjMzgyZT0AJm/
G4n0Hu99MnPkoDQj5RwfzonnQ1bY0K/Vt+IOFMh0HPH9SovKFizQjpdwqRlFvbzs
tw0yzJStQFmLWvqRDTnYfmxDNqktBiLUr9S36JnBqXG7JiNrRgvqexbL5od+KlRr
vmd1FBbjXhZe7Rb9hLCRT1fAIW97fEv0EeKJ54H1/SUF0QVVfJWM+nPAGLO43Rpk
/MwLlHZFG8puKJF/i1wUUp6bSkGmrJkVAXrcGTio/r9miBduIURdj9JPzo45TEwj
iCuLVvbLT5puVa/ooB53raMLeZYfu1XLxHvKvTUWaGB/2gOcv5uOM0CrB9O4iKV6
l7F9z3WH/A11eYTzVSYr+abGlMolnXs1FpNPf4A1052PvzvBKYSuQL2zBtilkOl5
UFMKudHPIEQpGYEUczkkjMT0BYrscSfQvabv4lUyynskm633rpb2yo/LFrmpRvvD
48unHdJ1At3gPAcMLrVKwntgBXNe0uKXB0rmLY+xfJFe9NT3/on+9e76hHeDoCwK
2vxKZwLTm2uA45BOa/qMf2C/oO9hWu8OtfnT/PuTvB+QfMNdWniVSm5cCqBQvuBk
QMo8yioBY1uFeP45PsYfXJTjgQ3Pl7HDJlLmRvvINKSol1MaGN3TPV5EEIEdHbw/
gV5WKuQ3EnjYNXZzlI5/XDlCeS5LfThuXtlvfX9WiCm5GQNT69rQ9cQzVko8j3Ys
Iq2BfEAN6ha4sxBJMc6wZ9q/CFuUslnb8lP7+B+sTPT/agNBXDteRaSycsu4SEMo
VnNl39dGfnQpS4fPkCbBicTkvjBC2PUxH+yXl0BxB08R3Rn+Cxg+GzuJassBl2Px
N+EqdkBr2ufPGH82ipvpXC3OafNtLt0RBJo7dbXwuhY+vfL84VsXM3+3Gr3XgGM2
lFgwUVD4uGiGz35oRqs6Xzw44l5i/b7mWhSfCjsfLYnNQs0UHFmR6i84D9o4+lne
ovJKJQRVpVSwdNfz0/DhjbzMpcuQDCxNXx3QzqI8VfGsoTwoeVHHsyxgyHDbh2lE
rEXQzC4UvGzpUHu5gXXp84XD2oLqBPT0k/jvH3wBH7YcpwwRbecUIftSn8F3qwzL
sDmPVnTLczAxqm+Jsx7XSSnqJ4UgxOMZuS9w2OChrvgY7DBE7Kpo140BrDIpLlTq
o67GfoVBRDLQBYDVcvwHYN8qZX83LisSEYA5OUkkjHCtsa8wvR9sj3GkIb51FtNP
krDDOntCQn86RrSs9IZ5+JRwMsMmHkY4VloG1AfIVZln44PHN+qDEmx9s0rgsXFP
NTlvhmDv9yeFM32pybEJyeqWG7e2lB3B/lqrwIIPVcbt7xYokm3tJpOiLW9Mbp1F
HgrSZe1iPLBctTgW4wvgJFXamfG5IQVbXEys98Ky+Cky0nDaBWwQC1M8NtC0qUzL
RuwcY8vCWyM5dDLdN3FuYX4m7fdcAF2S9WjiIQhMLnskOraYxWU56u4u4J067K3n
/pG9XyPdNpD0oAD85laXThM+IAty+J2iO4l+mZJT1RCRzjtpcIuj1WyIA/CEcwVi
eg9L0ZrRaU8uSre7J6DkqlZA5Fx6R00z3MsblAqhgrzA2lPgs0trZq4756EEQYGt
C7DSdPZNtUh0ItBNK+RNsRlgltt3EasJNNsT9wmq834GdN6nwrCjuQsAPb5lDZT3
38Uk79l42z4sNdoFxtpFB4LnvMVtztg5gDS3YmPhhXxhKvav8ODKxyrlrDzx/5CZ
MLB5pjV/N+158K64mvo0xQ3XKC0S6Vc3rIqdrS1xIq9ImdZ8QCMgG4TjxtFyWkT5
wKEdAB3r8WYQC80MTRGMjYqboeascJjkIX+GDzycXQ0TXS2A8EYJd4GXXxiC7IYg
cIRQesruSgvWWVo/ouOw5J48F6uSmqJrgb9KmNaFHJP+HN0adjREDOk2z7nidiGU
LTzuzIk/7GuF/pt8A8yyb/QXUMMy6rEZ9MTsa3VKbfqDPr7q2qStOc2te5MGb2zK
0wcFQsFSUsG9PVTstFOEscj8Pi5Z2jwwwtmUQr/lDm7WnaTA71D7XxNp4FKk2CoV
efByFGEC3i9E4nKK4OAOxSZ8UuXY6rlU4DycAFrSWK0RLT+Dov1MePtL0bBMOCnY
ElyoEAII5WumlB5mEmcGeAIZe0CkBZVIz9ph5pb3bbOsiTubGPi+O2Dwo60r17Vb
XmbgmeQNrcnmnUYtuYWtoglNlfDh8pV2Wv+bR1AZKzM6QvVGmXTM+Gg7lsRaHR8F
4oAC8+IaBUnefmxhZpx1vY5CfW8PdRLhbIoXCneYuqen7pCc4Eb7unrpBGTfkDSW
crd+lslE72ERlguZy30H/nYc8b2tNANqTK3F8gDGbJPoEwsvYIsAskk2gpwbDQEe
C3K2rjU31mq3AF+yDAgKsKPx+SwXLJFgcweiB7Q4BUaowC90QxgdECMHs4NQe3A/
bWnXnXAeJnkCzkF6SGb6FGD4H9HIAVsklnrkfP7PkOezXXW67pDFwn6mTsU/Hgae
yNKoIpgzzors1i63XfxTSADsbollac9UdPfu67wYGvVudAbCmq7omiE98fGXY2Ax
RmkAfQmpOhQCRzbv94QEAof24kGRHa58uwxPDbVbzRTd9WswA/goSyQtNWgvEbxr
T34g7clAiFuPRUeVE3LildDsw8VOUJQijviBC9WXA5TP5p2bHNnlkQmHWJwBMhSe
jywBfViCaKAuSNtJmfg1nG3ITgaV2zPD/8u/MQLR5TYpKb0Rlndepu/AN0XZh1KA
pyCjJHagJU6dcMN8+AbiCHQllFm0H/JKEactDsYi+I+kBrW7D6BwAyPCWG7Fsg89
4a+Fjc+WB4ejTPiWDrmqy9tEj/amW6/Ke3vdnhtw90SlRhhqP7Herykd1oS9LU7n
7WJkRjYdGA4YQLPuov9a7TjKAFBqC6fm+gTa6iUoBeBK76472lz9vvVedHvPLsBX
ulttmnhj60Y+rBSN8e7lB3UJOtQ80G9prEq2M+dr8Kr0GSLf6yXo36P1blTrRMpF
ZZdzR1D/wcKAvnGeVluWVcG2gxhAQKKrLFVY/mdmH0KQabyltbilmPjSJsCElnh8
KmYc8lowkD29SS8SQziI10Tm6wlXnAs5Vl8sdgSKcbiv+eiuyr5lvpgtWChS4kxn
feYBw2QQVbMBtCUYviweuh6qJmCqVKnIHkS+kraOI5U5dZG3pq3NVJxzeZK40XGh
/r8axIO2ZGme73HdnnQE+Fu7oMTyMCWhONr7NJlAQNChhMQBCU21wguBDsq78033
xEpyXh1FkwDL2s65JKC2XkZxXZmgSs4GS5D5IwnQYxYpyMGlppAkjQGS13vb2/H8
14bIxtxFVOHlEUQCcYzg9hz3K75X11SZju1ic11GY0yKvnRU5hR0EUFrB5u5BBmw
Z4CuKTR+FLrWw+lC1z+VtglWFsb+mODnyPqFGBICUv9TGy0IbD7nHXNDyaKwqz9J
E5nTwsCeE72/XSah6NfRoene7wB5xgIYLq233yBsORNfLeC7yhqC6DBP59qvifcc
LBQtWfageyNNm00xzcVQ8t8kEAlJTSqh523jEVT+1Jr6gnF/A6pBQqvSVwiHeaOm
GBooek1auJZ7gT7LbtWMw2U72tCxZe0uIbhPKLryXn1/bFHLLYFwl2iPtbpeRg8B
aICDcnOC7xn5CsOv8Vj0BOmRJujovH6OyPRqMfwXN9kJA5Bk76IQH20qsPD9RTMv
kkORav32znpi/43aUe9e6QMb4LcGqebu7wHDF4c1KaN3l+z1cYLgNuvSgZqpA63I
pQwfIbeywAPDZhQRWW1hls3ugdgPLiDLa37p97ShpLsNbAB2ui9Ji5E1SYgwF+EG
39yp5wkZeib1C9x3vI0XVoiqOo/6dACY5bgT048C4o5Ib/44jj5cczlblUDk9AhN
OAV10C6oEFtfBJjghac3m6RxPBcTea3FG0r/6nnmHEs+Gj8k1aMQhp7OsKhQk1cB
m0illDLT8BKDUtn1za9QIOVc3lWMxikQFFs8SbinTPDKOLZOc1oJn3V4mBrZc+t7
oywvArdHP0m4BqVS19WlDsA00DjIpUP5JAuTlmHvlk5g9BqDbBCeriYG+qv7j72N
6xqCaF8xkydJk2EnrEgrtJFTlf1LNqGU/g3tW3Um12JnQk1nrmjn9D8uUS8BYnD/
7TmQ0cFlpkGeov0SRWjSNtW360AA3wIc8gqlN/PU97/lHrwXyp+YwWV8BTD7F40A
J2vmc1AbPWgaN7hacdKYoRDnOkEyAoOxxPDepEULLsEJRo50i7w8boLCCDeQH1gA
fsdLtfH0q1zYzalcm/Xol4D5c6DnfBOoj3rfY5C0194NGzEMVFZrH/bli+q72ART
trE6BNnWjShrJIHONxGp8130/YEbmrJPvsCnjHKbo0hKA70ku3m01JwwCW53lKmB
x72aJb5bAPFJYerhyhaeuNllFzL8GTwzTMOBHu/vby2nay7XARU5vc0CZsirnnII
8gRk7wWz8Kw37R/dwqwUCQhxo9mChymqGGQrH2OZOhfW6a8lkQni6mvIaXkS7OZh
wS9idCADKGYew9m644VuRu4AiXrvc1mCMvcf8qUSgLI7eNqlmJ2vvf7KAsgmhK6B
NYzZWA4UPgYU9abx1Drhkj2+V2LKbiemdhKRSkOVZq2gdeuoIiT5gTl51ylWLPLO
HI1vLYaNdW+wV0A29idlMDwSakONw1hYbVYAuUGfkbpyWvt59Esm2WvtfvOqlK50
NCVPASycYsZeVEF7OWhduSuKOsDM+vOpotnuIekgwpCwfcryHOk5LDtDLpVZW7uw
Gl2LuAsc+9WHKiP4KHRRysMyHvhe3zM11TltcsacffalhZFVjIl7CcQ+8ui4Tg/o
dc2jLgRg4K75SxFKp/SU2dSzIK2QMER/9eKR9qYxpzgDMJ9Oqnd8E3zr3EDaK8/L
yiaG0pzPqiVfh38zCk8hc7zDraU4fpLlJVdlK55p5KJyR1lDN6qOdDYvdka1Heta
/dTgNYHz5JdePbR6d/Sm5oIk5TKWic42V0VyhEJroewpX7OAqFRSepW5AVGBKvJF
4F1FNP4eqI6nsK/o8nfSzUkaetGojG1pP6U8Lk5/SMxIWvWgFNaPZmrGYvBGNcND
UYtIGhSRNyNtkqq8UHsn8rV+M/mWPY31g6s9MISr4gid+K/o1jv/EiMENMuRWhaw
xK9HpaJonffnuAjefysv5GMWeV1FEWfazhxYUqXL8rS63oMrAPYlmLOzoZ1nlbVp
Mg6ZwoiCy/qX2nV6+Zhul5mWHtH6hbv77XB4nLeftD7T0gFj2yXizUhpVj+VS7ZG
BeU3jphc6Gyd6tLdq5r7vob8SwIqbi5CGYj9aMig05gC8BUmsj6j4NXGt5E6y8v7
wsFvfsIEhNV45o9o8HxCR3zo3ZVK0FflYTK8S0ojb26vAPz/cEcFcyboMNRAwfEg
+NznoeqF+Hddx9KQLJcvWvq5/kB93b8JQnSyysMUcPwGaUeWf3lAPd/3jqzDzCuB
KFtyx6fFf14c2Urr0VD3rL2NlivQgO3uLt3OnKuzdAUEAEzyF6SsglvPHS0VKmon
yST5z9tzDOkWHaL/nw9I0H0riWGEk320IP/Tb4oeyJOFyI5fP1qhyReFVaAETVR6
CeAIERS4DN/u5K6qoMpKFcl529PzWFh0/GHaysIGh88jstPfV9V1icpsEMQ58sL/
/6qkojNrg3B56/EVsaDwxKeHgLWHcU5jEYw9SczBGte9rUJ322AjzAq2B83OqMtB
yrEUipyspkGCDE2ij7Xd+Tq/g/hKtoxJiJxFv5uxcY6tLZJ/u6T5/DZjanai3FUm
2DL2ipty+Ls/IdS0C93FSRivivys9364fZ/nI3ykdTE8YpdI/lk0QYiyZkfeO4wN
2H8MWcxINvkgjC4tRyCbtSTU1Eqn3rq6rOJDJqS4+6s+Khc1ucSJLPo2Z4Guc21h
J1W4tRtR509ShNMko+2rwyEMV93NGkbxT3m7qVpV78yg6v/0gYgNeWZWNVKZGWsO
uV3+oy5k6tRWfGeFxfbKaL98YAVUqKc4DypChAKxdjjV4gemSmSbvST3P7sct/Go
I5kgjVm0LwvID49XYPWuzx5i5gGjg9kuEhgxRIYf5TCGCY7uJfmKAUMGLj9HeZG3
TLCCoimdzqUfcGxpdyWcEmD3FNYXmDqz1MOjDEmJDEB5JEwsk+clYtswkvRyK31i
fN6UnOywkIQqRfTc33k7JSrDjogmkm0V9+a+SoZWLm9aEXH46BMtOwjEGpZUOSZf
yFakdH6qaiwmjr3BOfUcgB7hChf6llzbMKSGNWJh0PX4yswjIQwQRpgKDI9kfCcq
hBJShclC835IDKRaa7vQrCdqiLFqCWW0gapRi4KUDnO061Trigzu2JRgkVFOBI7/
LORIE1vyo+ualZINwn2MWqOXKKoyWsLwcNOAp14XUgXS+UFcKA7ASFQP3pzXKFHA
57oUXuJjZ6fPfqQHxeLh0S/KtK0NSvoXasn+gHvm/0fjN7qCwEy3yZjC+pHKjVej
+qu5U9WZYQvm0RFhLX6RZVG5Z/N5xsse99+4NVbRTSrH0xJ0d7eBsD9+HdDj6+2R
eAF0bvNFi8d4k4rp+L2++8Nz4FFT7Q/ZtGsGzXfLS9PP4JPxFVBbHSJ21azH/v9q
Dc7jeGFwcPkr18HIpO9/jwWm9rb4N+a5j7OXaM6Jjf1FVEkL+1C3cqaFyROoJrvy
o0HGqBsvCvIHvHk8h6rTOd9v9tRf9VrolKIcqN7+YUtrjHBdxu2CmYLtxH9MrJd9
Spf67xEidE9qZx9L2iSv7zQvy4iQVhKSOPjDQRycEA0EtVYQye7Ewk0pRbwwfoCF
nVR0msFS3zgtAnGQgc+hRqrLAQYmr+TvS2NIreTWsYpq/uO647RsgBT/YYCDJXa9
+6lSzfZ6S9C9EI90hr+h7f/nWGwY9LOEkSiU5YSQn7ixxiEz0qu988nFu6NIDMgT
TlZXFvhxjNoFsUOLd0ZDjpbTTbJmxUFhY76AbLT9oYIP/4dd7JxVVI2yM2xVBc+k
XEw5pPOr+JFJWdI+u+xV6Pkv0QROtzR7pRZz+ONr+Xaa4UlJaTBSB9aP5oT+h2A3
BejbGaOqbyRbJtbCqjiRfRh/jdvgWwIpTLIyxBgNtDvxkk3xmrAeqjFZCzDhCz7r
aSmTb5NbZG54hmC77XWfVe5Z19P10rqnL3Tyx4+F7q5LyuSYxmPbvnlbRjbgwRXb
pqSMo86uLYcAti0mqv4Zfy1xpJPHb7mAs10G3jy9Ot/z7g3/swn0iFsj71KgzyiK
yPXjy+LC4CQ2yBIbHK0dHNqVIXT2sdvT9310g8yAUWgT5Mg8QWLgKXVCij6VeCwH
8gyHlqED5zGc+TB3XntTgbdb3P5eaMYvSc4Q80+JEtldKtfbSPvqafNw/9h2a66I
tXsnhCvUH0PXvSrtPB8Xz2X+Wom+RDECkTzf0g+z0AzZ5Dav8P3nCcwWqoFxJWlW
Ja31f/RxkNEDlIZTLQ3zjuWoRK3ZF0W4avBCfQXZ+RC3s2lxaS6chclIqR9raeE2
GDEp/eLPwevhGoL8SxRGw1kZ365RlNloZ+tp5if/2/O+Zr2VKYcdaj88f7Xu3jEX
/WA8J+S47SDt0mjDmd7RY3QLv9xuMPG7xOd1gC/ja7d4S4QaCA5ZcIUrdTIH+sv3
Mt47qMu5ZEL3vJ6P0Nj54kRwXx8cK1q2XcxY9DTkWlgZzOm3XeRsFNvVfkbg/Ood
AHcEOv/4nwyQE3RcR3t0Od7ElpBmjIMIBS/rW2HH78CFmKPB3Ifpyg6qsnb150xt
d17v0mZHWWUtRP0YO1D7f65uJmKSjktzz1n6DYbb2TT3eTTxbHrWL61a4pgQOXDy
Ko/RlA/c1PMZnpxLt+tcBeLewH/BiXvZYNHWg57/W88JD0JPHVn9h8y8ZlJFrK9o
rFfgJLhRh39N/HABIkNWqce5b65suDiyqsi6RYRA2gYlFI1y6tp3K04cyQOTs1YY
eLX6igLKhTE+uBZghO8Wbv0dZ/SAqW1p8ChRocbj/pHqxtyKfRXRkTcXiD3AsSOn
2i0PTD88KHPtRqQ1oe96CuoS/0MI9tZm28bb/cjvm5w40cFVxUMgTRN/qYbncZ4G
pqHI0LSc92h07R2owpDqA1KnpZV7N/+M4dAVOllObfd1X2KBX3a3T2cE6O6l4jyM
G7xhOr9/3qjdwcSAXktjP5HbcukE3OIUKuC8ScJTlmPqSyCyAjejHpYBP5N6JqkI
iNLO4DSGaAR6R/7u6NByhxmzBGEPSNZffdCy8B8ABgBZEDeFhnnWaJJ235S19VxX
BAqRrGfKBkSIvx7Cbfqrron1WhNTEvbEHUmkfp3z1EPFht82fTCzM/5SYgiR2guT
hLYl5DsKs+OqsHQyD07EFRBae5UiXNbMIgNvrxMvhqd5x3qVqf/iuVKUFOliw9K8
ZRb5OlWRxa7aOml7CHGIMemwWrWAevq1LQRdMCmxEEkTiRSdDYNz1BDrLI9MYs4E
oe9ietb0UjjnsLWeA9yFluKc+ux2LA3roVae5vT7lh9YaJQWW2RJP82rNWdeAeR7
6CpaZCJbyssB2PvtqleO+NsxMId0W16hgK1dK9wzhGrYIA093A9TtgmWRvu9OwLG
mzWFcpSE9uaNLFZhq3r2tTv3OhJa8kW6fWG8wE918iDEegNJfv99ltcpendy/jr8
a1pjKdcDiJa/8bOHxFm/pyr/4BckwMKSe7IE8+7g13ao5PA5vddqWx/dYBZSyox2
9VyEH2isfZsUVrXL1Y3wlGUYbvjkyUIXEoI/9phXUrncu+oLohwQr62tujfzmafs
OcApOcK0AACoNp/xe0Dt3kbb9VdkscSN/Y/4SDioVlxdWIPHHgI180/QgynxGVs7
XPSEMc4ybHmyOfz0cxxw+41DE+uoCeQEybXIFpFqBUepJOygrdu5a+6BAawc6f9T
b/Gfbgu1NV95IWCP9c7Jk/BXeqt6zoOL+ubndnpIWceLPy0oR8zw4y15XB41Yz9X
jURbzYNAJfFgMPx9FbIe1vEYgZetW2pBCGMVEWLNjb32H3Tw4JOt3b+6C+uWcN4c
APNmgAsgcpVahQ/Wg+YgwD4nl8vXhONAW8/vXnFd8jk8kqpCxC+ipMAEtrqQgH07
iyeJhT0I6l80qZlhZSrSQ/XMwLehbcTECcdgz7LdaAQbeEPAdIqVCs4z3I9gKc+q
gb2uoMLAKifWac8yGquRSpHfJiPZgMy38zfNbt94+iHkQ3JoJnqXThIe3tbbXMDM
qgX6k9uGIKW1c0bKyY2vbaKFb0igWlOVb1FrbqLGuZJYSfbdGBOm7yjuaEOkcAGt
n3+OMNwavSw9M/e5JfMyxsox3AzOCwCUxdXLDgo5aKkvIc+X5/J+SlEYJ2A/T73K
MsJXH+8aU7/ZtgJjoktn/gUqrHMb4TNTSwAZMJVH7Qri62hme0f1HQYREQvK8TEO
2L3OjUXBm7mpzOJLKL1fpNHLnginmejR4ANWQVkBpAc9kT/0LJy1XF9qkhkOfpyk
KwmR3x0AEtu4H7YZ1C43XVjnviGx1axXJ9OUCe1WOaRNfapx4VB05CZoIW49+asF
aWlqVbtxDJqboAhFiwOgwjfAXnX7T3FQxj52uOoI0m1qY67aDw10qvma3XoYkIsT
MgJgz9zN2PdFT1wVU63fT0RcRIkh+1zuLzIdtbhqawco5gM7pA2sKGfAgcJfOIcb
wH9v+Fh3zl6Qln4tylEULz2GBYaMrQ1h/UV+yhKUOl6WO61JDU7knwcZoyEZDNN5
pudnAchIcbJ/ecK3VlUR+131b67gThmaYe1NQ+MeMUIPzbLOWK1ukZf+u7R+4Elv
duu1NZeDHDNZcaqYDdAVmEXlExVpsBDxoh3irCA25byz4tTnxcZ1JiTUG0gt91dd
xlYcKmlJUJu0K5J3EJLHKCgbMb/QHfyt4btz9EQ5bLJC6ibLNyokSEAPJWZlulYs
c2mOw9MF/Dk/6rDBldOnholG0QVnu6pZ3UGL3DZfbzDxKlvYc7sDtSFdBi+W6bO1
IBbIMMLGZVztsXigtWlDET9YNAI8yjuPxspUiV32Q1mP0dZqJGMNs+3mZ/lprlQS
aYSEEV3oNzWZQJwqAaV6ueElzzprrjDAXW7D3MWwWQSIesX/a3UDli4VQmieFOqh
j9veyCn6lAS9yVYNSvVH4n0KCwpzYAQ7ewP+tHZ4L3EznMxCEZjdupt8wQiFpv6x
1D2oSqvM/UyV+Qup4Vu6Tv48IyrkBOzYzajqzzqNeJrUPFoZMWSGv5kvqBRgdJET
bCd3ZCxSnkiSNYcZUhDZ2LBqDPRizWJh/MQshuTIMHHKk22WRwN4borx8SWr9k3R
AFb1zZ+OIp+UOTCpMp5HKPccwAHFTSJhUp4vdqi6nAaWSHXkTZirhlloz4/dKndK
UJB5GmbOuzqxMn6Xam2J6QXyZeZdJZKhFlkkWzNAvtRXtn47ONW2uTntwAw1Nl+A
uQ6Eck6cG8BTwKtocsYkWFGKDDZR8awUbCO10EaQPk9b2CQB7qE0pCjiSIitFhOK
QLXqqiyqV5i0IbuGCPdswCsFtMZob85VWRrPnash32wtcWDj1auvHF6qk6Ij0jrm
hs0SjcXnkbXZgv8+dYRTd9vD5bku03BRCu1pCKU7xwLnU7jD9QeXN55RGRpy3iuh
HjQ2DaJlAdkE4bJp+AqdSfxKkDYsa4IdCm6Z+lfvR2Rkn0hoLXzQnlSoqPSHx3/9
XdV0Iy2l/zTm6728Dg1CylUJEleYW7DkJHWPx1Ymf7cPVDVa0p0xTAbJ/5dguA5w
g0OCtvM5zTcgt5QfIZiaE/wYmcU6BCRcGn1wZknBc+/fASsFKynSyAXhK9z3GKGn
u6Mr6W7RfpYC0W7EU3DO5w52KkOarhzbCDhJIiQN50rKTawTuzm0cByQkGYHFvXv
FvJAyDKbv/Cml/eJKfsYLmQqy7vM06kp1s6soDDg7dAa4C/E8g5Wj0+A4BUOg/WM
Z9dcTgGDgvUr2URwaOZNGoZgZYFuSK46Kn/7khUBiyzjBdY5kDVbOXLjkeb2rJM8
ssnovUXkUtx4ASi9wzMmKIPYZYoK+0kCH5baYwkmkC3K7DkweWyXY2Paylh53z/M
kyyqXLg5Te3xTW9pXoYK4HtKliD7Dv6+R/aqxJsG58r30CW3TewiqcQqLWLVsdE3
98eg3Vddy+smQC0wMKz3+sWm8jsXTebANyAQHtkV72ortVxQrFflz4xE+fg9qnGR
I2Hud/m2BzZpwsggrlyOhq/HjqAhUWChHXOEAOOc69dtg90mQGlDlkOx+RXXE5rt
n00GD9JEuMOs03egyFVonGDl4BdQG8mxLYkyInYmYtbRBiWVfL4SM+vWoBBRLOIe
M35X1H2aoB8fXGWlWu+4QrdnlKSgyngdLs4dp1y6QfmLcnLWYaZSgBs84QVTZGCa
Il9vdnOFHSHhiN29IFneoIAiTerPrXm7DjU2r+b2y90nh9kOrESpVPZaTEApmXsS
Nh/SvI+8fBS39zabpzaE6FTxBLmkFLEHWvTNuNrfueNUdtU7B8PJ/2BwyOlv5E5Z
dL4uztJlT81Def6cYe70Ire7ProvNJz+9HvCn8L4C7GVlO+gxvomij8jwJ4B+/el
KACsD75I3Kuu7n1/jFvegDLsLAkEIXEhd1vFzfMl5K0gx2rZ7Ehq+c1ZmMfvOsW7
INQrb/UdKcLsKq3ailwyVNjS9HuOnJkrEpFQoyDLQUqYsFS8V6mVh8UzEnTmReLR
4nTmZW2ghDICXj2khAVArv36KLxKxwzSjgS75gEsRgtC0mfjh52MlUnE740wR2/W
zQkifVYWL7JbdRssbkX9hePEyNv+bhPOa60gy76obDSWG5N+ulKxqbf+DMcYoy6c
d+0qvYLotxlybhud2D7sdJhZj63rVcS7Giqi9RsncJ/dJZwu5oHhyEdm2AnUelkw
SlrLKok9HTjQKH61Mjv3VVP/blTeG2d+xL54KaVj5aSgsnWUKWVr1kDdBBG8nlwe
v7sjuD3uDQ26GzwAo9IssvksUtjyGeECUuB2wxCYF0AKNBPl1mhLb3nqBOJe+Y2i
/p8cBGp+59wfBO2oaocSOqXmeO3/n2I9T0Y1vmIjEQFlujj5tPMcPtbDvlSfFs0F
7Esa68XkpRBYuyJMJOjUy9w+t2+6dnGm9F2cD+aoR5F/w2ltiX2a4xDCnCEAvpm2
CfwXWV2n2IxevTMmX5hHxi7ulRU7Hfo6Xl+Ucl2tzRqKVjG/DQmIAH3SKHX2BoHI
phrxDPW70cvCBVIKvKHN8Taz07uIptiNN15OSKK1PT5NJ8JwqG66g8ulVH2fCPNp
XrD9L8G9W6KuBK7hOY7ImSC7KUsHWa6mOVbyyu0lHLt5hPbvWCjlzgs6SRQxjVwC
HpM3d5x4lX9b4CxdsK0rIZtTYBIo9t/ubB98mmCYJtv3JJ+CVRlucmNw+A7tODbT
uXmKuXRTGzi56uHKiB0ZNhbP/pe8EezWOqaAw9ePjYsl2C5jqBt30PgWd7EQBfzC
9+9KPxSBOC0VyZfAHn4HWHlx6hiX881W1wQRbE4GQBxvuMv83/Ixmwe11Btj8a5w
fRG+xdhElnsf88DD018/4rjFoGo9Jy/2AlnbpW/H3KVF7e28TtlvkQD+XdpMBUqP
OZVYgUgQ6n6DlGJvpiu1zJYRi1yLmX5Wu7fKuQvAFQNUaQj3/7TAr15kuhwgkMle
98J8XAf5AfDhCsssY25Ify2onHYipOHOif3HKw8BJAQK4f0b/ha1fx+DDW6xDgOO
HI7odaqlMQ1B2Mp7kgNGWRfDeVrVYP14O7tDDt6xzUBEsRM6gWkrXstDXKrVZfLM
1XiMch/hu4qe1bgl3Cns0S/NhbfBrHSqb+s/1dwzu++APBvsbfcjYk3h8dzlBcCE
/ixj67CO9vS7a2AHudUcKpthmjyp1V+JyZM/c1MiEkltwXHBTnI4d4JUCS7m8Za3
sF080NPTmHfTOK2Fk4WZMJD+J1snzQXuAgyrHgK30Hx+PbC6YMOkXYFepPLVnmhl
L5vJmsQwqQN+qa0y+SMyQh1TVqk1g016ja0PTF32ymRzYF3ExiO0Pzx0KN8CaWxp
ei3eWprdp/Fn4KPGOMol50HtAfeBTuxmRPWxpo6XGxyOBzRvOtLNaNm4p/qWCWCq
Uw5qINA1rPHb+jtyfwAG3vRWiudccOAIbUMsPEX4QcWABRbVeymWEO/hdjfKw0Jj
makfNzPT46dW7z1qNys24ML7kiw8P8jnKP28/YfhmkRQHej2FPRvWHk4lzW5EXs8
Q4yYtnOSjHryAA8lZi+c1KrDsNKeREu8vRbOPNMh2Z0iZF3u1bh7n/Da6mOR2mi8
LTBLfjX6c1be+gsbSOpL+HPWxYPry4BH/OToGic9297XTNRp+zA4HyfKZrByy8B2
Njm7aRmFREODNqhuehuTHxAoQybaJ24SzKe/Sj91W181X1ODhPOFjrYdA0C7iASS
zoVxBh6G/jVI1lol09oaK3acv1IHH7ONTunmVHoWZaNmibbpqWTy514Crm3RduHQ
CAvaVVZEYMxZQfLwBeADN6S+bMWC5J7mVgcHH7ryt0jRdaTUy+ORRiYZ+FQIoAF5
pjGdLSEiceJs3JkIvcBKXFcbiDF3RYZOraLlfJykwVQy3cvc2vvbQ4011IFGtJ3Y
Mmh5YBOZgSTt0XDlbD0CN5gxw/8vzA+aGiwnexmqSBHBqR2yikjzEbyVyg68to56
kt/KFtdtiYw6H9WC2xhzhzo3/riJElkUEA93BYYNRUihurN5brAH/6k4WfM3UzoI
oWyfGJPJe+at2pIv0T/Kb8IxhVc+4HubY89dOX2qTvfUBIjEbAUc/UhDIPFiPcNC
RVeJBNJEaZNZTHiD9V/6ql+rvMt8Ig5RT6qU7/xpFwe02y41L0nUVNgiKRP2OCyM
Mw+PJQwb628kZ3NLK393a+AC6wIlFLaREjQgakV/kdhidffn+oFBf1SX8p10fXOc
Ptwi3b3cut2EzApTqK09WKYZOfo6BQgxHI3UDxTF/9uA9hb0RneZjZOEdSq/H5ng
oxPxOJPyBhab/kXJw43IawESHU98WBIdICohIA3utawA7vYF/wr+0bKdysoOxEd3
j8RVsDirA/aSYL1uT9R5bpsSb/Mueq40MFKACz8Sx0WCCz4qhBkPW4t/s8zDetzB
qneU7ImEXub1PDJiw0+7txT02jjBdUkqEMVUveZ+88Ii0SDo2xvbFVVYW0vJXZAQ
I7dowU70RYB/CtVGOfCZM0YHeVw/rvmrv4o1QDZu+P6t23LJ5cCEsCmVyS5L/jxn
n6VK2suQlD4znmyUqLVFZGsd13tX8bm9MoWujS0H3BMsxX1JOa2w1xV/+D7U81Bd
JroDXjaEvs1hiqGL2UirxV0oNo9Fl8egMaSrq026+lqxUr5drF0PPPv/xICdunAV
L1zBhR0wxJS1AI8Eso+wGiBsKTdq15ktFXN3luvxCumwWqfmKlarJlp9yUM0Sduc
mUwQ7+DS6gUSUWvKVTZMUA2+HhwbIxWxVSGuDF71pG1vkllKrxCbsEQSEP8g8BTU
O/dBNMY8kJDQEtG+o/FRx4gxbBNUBwjtHvW1JT+itThYr6QXGm0qp88tiRybVaP7
3yrlMKwmd+oOQ+O8XRKH++kHI8ARxbA32KDxtg8FW1R50Y/9BsUqrkjjPQ5ydEt0
/one+YPQDQjsqGL+AxboEnaWg1y6uAjeQW3F/iDybqUJzn0PBqySjz4US2LoHTSw
ntJ2GnFxqS4MKF7pl/32VjHPovlebz/XAnIROsukxna6DAjVEH653oEM5KvaVRPX
hh2W52MxCfAWEF2fsDdkDwQS7kXKo4Lw8RpmZO3be/Mm5FPgdAsK8qFI7MUxq3wU
inf5ts+eluAAkAI7qgT8ID9UafV472FidaAttdRV8yMRHFvRHd/VbEQ3+MSc0Rp+
7fdVHmWRMAyHcfSqt9mIcLeN0ywSMpos7JxJieoCVCqQowwT1YKYnX3/+3xhfZRG
Vir54kP2RkgNgMnq3tihnm/hFqLULtyGH1PEYtrN+CN2Tk+l3VxCchis+vjmlacj
mDR9XAQ+Feb5Cd5RGhZQ7XsQXCLnGteYOMWWYmzNrPOWpFfR10OKEqYcUM3XhvpH
qepJgvgEcKy+zV9SX9AJFi4ujrce7at3gVu/MmqI/8a0sf2k+Gjd+py0N+VG/0JT
36DvemQvu7N7O1MijoqPWUmKS92w7XgW770y9DBjCbNMHMbRictI7tqvG+HRJYZE
Sbhwvre6nO3D//QcHHNbjtqzJzE8wgeHCyBf2FJkfMwnjPW1eaFAo4jVm3fc+qxR
f0OAkR75yyaGiCn78ix/evyA2mT84cH2BkT7u+Asu3jjkpW1UkWJdGg6icn8ypDd
a1ts/L83EeiD33v6xcvs/iQmHDW8bZjOpwgjLb//C5O9qUn2DEINLpp40jYs9LOp
pcHur+PE7fLePu4fCoKZIo5fPlRWisATm1p5rVm92BtZh7ozXVV6XlDHngVtkJqO
XEOB7CtpLUx71LgavsKbgZnZSfe06FqBdtgi37LfMdvj48TzgSS1bZBH3U9WKUYD
NAwL/bclUB69O17GE/in4kJLzz/u6y/m6Ag4P/JrSzKACwGWLZtAiLUAj/bq9UHS
Uu+hAj82jpEEgtAau5A6vt1CiLt0cdTkNPG1CMAgMMmH9tif+8vqASfgWdEgbnLq
DdzDkOy09qyDkYHeQ55uxXftUOu7I/8iCkRuiyDFyIhcvKWcPTf0qs8Tjk5IV9Xj
B/pmFD4zL5ZhTTU9Gs84kCrp2SVRYmLnTPwIb9L1HI/RlsfsIbrbGRtP7aOazUOV
Ir3PhhGvKonmayO4HiHzx7aCRKyeE+dQL4OyAo7cP+PTPQtprcfyxCSfMRNAU79u
O3+Y6kvcj+tdQ2nrj+4UBNI9bXLieT4yU55NqBQWChc9xHxVU+ozRb9GIfDM1OsM
R54hRm1e/OZtL7Vielw3dpHyagbxawmyVBitsQ54TzItL2cLhUvMyRgHtWVEo77m
rhHvlZGV3s3DFP6MQghKSpQAutqM1H0kO2jKmk2BpsXP/kmDBpYPNsSe+4g0QQCs
DzPtc6A0HSGM1TrIbYMaqBCNkYLgL8NUssnoFPveIuW6gRMNy6lJ1wTuRY1wLASK
g4wvvRq4Z3ZLEAU2HPNuXe2gKbqXoboWpIQbujKs9DgRKQXMhbk2edyLQBrTTMD6
HjAzB9NknRG+0Qti5zL7jWD2aX/pFlHxhPYpUjt+PMd+wSFz+cV5By78EP8/iJdB
MRQO13umzWYCfsr5s5muhK9PAGle+sYRBt7oaAv7/ldFGUyAUe+Iuj9mD1BvdEtu
awShVmu/tTXNalGVHI9LFn92taNAhMxgrsRFw+D8DrDRozy/u1+LQFkm+80QI1oF
ihwQDbqzPDUZ1GemoawNgvTzrClnAHLFxgoaLjP519vmwczwGvIPE/kYhbkcY6Hv
5s4EIzPxXwpFvvwQVbl8IJroQdvbNyAsx5Lid+VoOiIQ834vNrBx65Pj7ZCBdxSg
z1n+jwRaySApWUuFn2kwpFdGAMxLFu4+1QIaJTWrzTv2GMvAiusezPXTs233D7m2
1zsSPhfMF8PWO0pb0ouALKrY3/Fyjh3h7C+86Jlx/K56WLyN1hzzhGNGz+fZ9ojZ
3Agv4jAOht4fT5M6F4E1n/e9iBsGEmFHJl2793VgRdl0xNOIBC+xHeP0J62vZRJ+
jWX4PkUA0MmF02pJE4HIcA1a/aJZuiRFKwVRywn5qiqRCetyqGXZoi+vknMW4jJg
rdzZ5/PXQADT+rcYbWyZpc7inPn9tbutSgIfRXCIehHepsgFM11zQRncWdosDume
o13xAnFtHV6NRIqu/LL/ZrmSKZ7YGqs1uIK3/Jw6T48r2o+GFZtGDShhgG0CopyC
ddsDh8mHjzZpetBuSPWKt7kD9sfKRNu74HgAkglE5pAcXQF+qXMwJjS80RxLK+1Q
75Eayfc/HQoMUudqJ3vIp1e8VUwnelC+cBVNEJbPHV/YaSU/jidpMy1XOZF2s0ED
+PQ2+nly92lMKq/mWhF6UZ+9cITef/2JeFICTLbcNcXUwPm0dl9zVn21BRKZJ9rT
1sS1HtJlLkUMvp2FQhVp+DLJ2BiLcMoc9jJvm1rqqVIPKd0XqGa+j/xL1QC20NGn
N+6uxlv4bJGwVgo63fAufCez+VM0xnTgMmohbzWlSgVA60NmZMJeXTXtlbU6RP3a
H6Fx87nFVw2pv+V98RasVrh5bjxfHYaF1lwJUwzKJ8Bmp5T5wkIJon457AhEmYMH
QSPY9+xixmWV+R6E0IeqoQFaEjeHbJVmsqn+hclOTWePt4HRapzuRCbz9TYyRx1/
L1rLD9qwgJ85iL6LRadLi/uF/Wd/nL5GVi9WULr1MCj7PiMw48AQtmXyL2F15OoC
J143D4ZV2x0lbVLZCJ1ezLFFiqm9DKDigt1sHI+4S2/+Bko5bUbFuj38yNEt7H+2
in7qaz5SeqTaYsafhC62ZqMZ/TNbVNZLj8GN/pWw/p/FevlFuYDsDj5HYi4RS9ud
JPiIzsGLzIbGsTRk+ZGqdy/4sADQo2VqrvRAeASfCKKJUd3MoL6syHG0V8yJ1/g7
YzrwzDtBRxvz5OUOtYQeDVLlN4KO1d5G4TkX4q8DcOfJqTTSwRZILs+SNPZpFH6L
bSLNZlH9D/zPJoIeZxm30aglHa5l1QJtlVCSWLKzfofh0gSO5OUh9XKzU9SlLp6U
1csdOGGjNGF3JddKRQxT5P0DZQadXdrCHzsrkPeZ5TQOF6IPqmp9WJi0Bjm4Ryby
TBpTku8MYWlq3t0aA+GV2DiCUXllC82Dg8nLlzKq/NVZdHYBMRha3JuVCYskimWa
awhlQGiPCbXpMDkFuDvfec6w3aLpqk/rmR6FPiTehHNxnxv9PyEvt5W8N9/AngWr
5ncen4EfG4PmIKiH1D6mGRZMUGSwUKIU1S8AefUF9Gxmo3w2Mq8iAQDkuLxFoWbP
wh0JqlOs/snbAlxJXV6xamybj6gNtaj4mZxdq1sEKiKHx1gFZBh2XN4EPfurWObn
1Xg/D6mOjQ78HiAag4H7G8DjSPsRCGdDh2PiaxpvGjgSvb5T0vgcO+XcFp7aydXX
IM7BcZGE2puu6qWekdlNChKYZuKMceQEmmMFQBdf5YHolOyAhEPWWm4qd1FD0s2L
9BQP8FHf//709shc8NNMAQ/MNlYYNlqA508bSysTRMUCzvwoj4pmKYiiJBuB7N9m
9xXHCQPb+NDd2b71kNipRs7zUjo8QfLR+SaxXkmjM0Azml7ZOMZBXrnD/Rwe/mXe
9z3uW30RWboEHD/WDg/+N+6BbJaJreXgmMWaAQ2dCGNJFrNrz8wpVTLjTslIQJd+
iVoey2vDPFpv09/cAP/98GIP3Rq+anG4DabL34lmJ7fEjA3onFJ96wD+JIl+ohJD
ekpy8XN62PFki/6BpBSbR3N5exIvjK4zZ59pS9SEvnq8cfLkdwdkWxyfMv9ywhR3
IHJJxWuVKm2dRJwwuNAGshlP5CEwAt/aEGQnWwiU3aluRIhTvLijZFXfZe6Qe+RZ
FBCoK4+liOC7oiyZ9ACg2h+lly6GjgWRUqpIG+oN6qto1nnqwNm7NdXgtMUbAxos
rZGbaFei1P8y3iGjyMBs71R1NwrvlP3nVjloCqXT/EYdvxWMcj3NSKk3g1uyprig
FeTby9fr4FWpSHluuY/lP2xhG6ca4qfjMgw/yYCi4g7qVndmzX7iNxpcjfsZ02Du
T4MjLEUvl7KdAr3cHYqhIagEo8J5te/LkNPMoRbI73QJMRkQc50XBlY2QoRrGs89
SWAyd6TrfiI4xB/TyWEkbZ4QUEVV4q531ccySgHD5jsxmXX2XZu/TjK41t0Lrx/z
1Oln/8luMm9qujq3gnPbT5tYTR2xwIcsMo1dFOxg1bZ9L6pugmEbsGeR8rN5tTs5
MDKpNNHIbqXrsfZimD1KW0zShW61r27DjuaviBQRbIkzaEayUIIAhRpvOuP+Lr3a
hYXA/cTtm3ERhqSuvppLOzx0PatUXalatN653pZF9ovkniozczGxYKP1TYdVajpq
Dzbh4xWULE6zEmCzZyhnUGKXt2HL/j/WPup+ZdXoxWHFTdT+RPht97uwas0W+0hs
VJJBaWr6KMJhDTOQQoPcuA+svb0Pk4E/Aq6rgTrHZcohsG8aZdGZFDUxyhH0cS1i
4rjv1bfNTiV9tJlddHyiVuWwWT4kZc9M7nxyQ8YLMZF8iQ+ryKMbTv6X8asvjaip
gbLlG7lynPZmdCxAGPYyqxHBre6f/9OhdPVE4DOLkJ2j92ztLqLhGWFk0QfW067b
mZ3vJyJ60EnjKOC9XSrAzT8I9sCtgzFH3Nel/1htAJ10APPhA7ym19y4deM+1ssr
HIRWroAkg4TFJq+4x/b7zcVTCwWa4zurQO4o/tJqoydO+XOGGtXCqH9TWhBKZNUd
W1jgBqPXY2wJKG1kNEs7p270K6xWzNSF9++IXbgVQdDuWiQuQxIawnGzewIDqnC7
36YRsInxs4bNAqRViVEIReHGOTVDZSmzQ3LeXSPJ82XhOOozVNrUg2UKyo5dB7+B
+uLXpYvArct+32IlitizEnDGdQXWovQWp1Fg6pKHfe66MVLEvE9Zh/jAI3kX3mlM
kQmlesWeAeZOu17grfpv99qzRFAxUnJ/+/hHMomn8ho+KUu6WtsMs/iUjjluEen7
K54vrOVfsyUSB3SeJ1bssuFo0+MNG7t7cI1LwmHFyH65LBiF7NM/4seRLdMJ+E6F
XVoqMcD3PO5RJmy0vrZKlwVATNk8Y2VkLqEEU5iCTz29HaCJMSg1zYjiJ8wTIc7i
bgN6Y2z8RB2/jAwafhzZmmPlGWcchoQmvcr11Q3aXR8BNPaM0BbcTSzNiOoX1NYo
gs2Fu98FR4aCzUmXtEKX9zIEmkj7QN6fj0iOEdV9ZYdNDCrJJSbI5g4ZwzRgBF4F
DrJE5Ad16OeDklkmgDyb9izId8XSRXCY+cXJLlKREPCVWXxsnNj0yGS5HclBOjiK
JQ2rvTX9p5/kNXrLx1XnnrmzD+pbOBLv4boTIO54hxTgqdyGOYIE8/fZGI2QfMVa
R+IDgmYy0+oue8khT+UNwVop8Qk0pb3RmfTaPAuSwnaOYr4hyi9U5Aeys3jy+Y4W
Ztz7DR/Y2R6/OWMSPr5VuWPYNWdcpOONIqbfxt2Ro8aH7D5bj9csmp/YniHyhoty
Fd4lNASWGVAShMDF2eZaD53dRfUImx1EkRs57ttYeSyHOkEzJ5ll3jcfPvXMEVL7
8RzK8bbqWf/uxGy92TlJBN5TzjiT7Ix5QLDrE0liZkpt+of69OLYV8oBc5ZTfXhy
ymJ9FZgjZWm63yVWa/h0SAezjX23gNIqgadGnq1kC7YtVYXxFTqbAZFyuZ7d5Z0v
yoZ4w4UIV9HKKIuie/Yae7D0aG5ZaS8yGmRk4ADpZ33u6IWOkivRp444vZ6y40/t
Oo2uT127CeoYEYzCgOSGMhgjCMEinxQBgp0Cpy2yaGD6lR39bt+4dJ/YA5vrc9wr
0s3G0DVF8QoZeHBTe6D9kJPx48sZdlqBgyGsI4whUNVVwH0ln0bBZZR2SlAFJnil
9lvDNeD3alesbUErQzyxasiyzhRvy97hGUoHNZKYLMN992me81cdUwaIe+3W1yIO
IDJ3bz9r05Bux5cNhjYTpxpd9qpmufHuZtw8/YrNRtksathw/fERm7BaiGKHDtaX
HJ1lDBGYpJYlbh3nirXtBoa++eqdq7RG8C2uvioz+b96cjW3PpzwXKMbBYeW8HJj
QWzzoXtsU7X9FyvugQ1BBjiCvMK/dJYQ+2KKlAth5sBBGbKFLBZ1v+aNfW0BtDpJ
FMDFHbkDqa4yLC3dN49IUTdQd/K3MOVFPZcDHXmehsFvDD+fRGammfKg2nU4q1ld
vUvyBCOKFmLHAtOdMWMHA4JuNI67skIJYr/bVuUv71fUyLg4oGMHC+VCSvOV8BnR
9w2rfC/2/2ZuL3Vakh/K2jBUJqqsTKT1leQTmmWnD6GaiDEjc1eJuJKpcRCn8T/6
4sZZ+IR2BCSs8lE7qiLw8gbK9IuJCbSgWU+qq2P+c2utLwxuFfMphLUxjQMvASq7
iTiIxszBTeWGRH/8ZQXiZ++4YvUmMtB0uCBsnju5Om8AUE3NF0CgfxDieUs3WDLq
73nVg+FDW6xvoI2Jl9HiViMAzPWzY0suLdq2lVdjQLZNkLMK52pdGuq8oUW4p2nC
PBMkU3EmJXbMJm1ElAag4mHUp8XRYdYk27wSacCdQ0Wjo8nzVNZ2vOHo4Ls22Pdc
ciX9uMbetcskb7nEsCZLJvmqRtfS4Lr5hIP1RgHOtMRl2eytMRGlx6XCo1l+fCvc
Ub/vv1HhjSxIVhONhfBUkAx46RAq5rQA1TA+Y/hg0ORcRdxoEqCxvsuJ3GOabXil
oeACJFZ1X9Lpf6Zu/fm38a2eWMQXYt0CiHqacYPpvQDKXDS+MVcUr1P/97C0r0PO
acEsNuNeS9LvHUfxvgYm2spPZHwuoeqfojsAEuu2x7YszfcMnbSnL7vSUC+SN7Ax
oMDFxAgl4BryMizE9YFZ6bg6Thfunz73m9yWzgmBWRcaDuQnv47Od25Fxlx31KPN
gP6qQ5MahQYxA29YA9bWtEbcL+8zGPrAjvqAzHhdkp2hHmor9Qhz0KLt9btftE3n
ANhoYdIPgNJmbdrXKrb2xL73ZN0qXzkT5wnhssJRqfj4zbsviwVrAgzqvOryzWhI
pYINulG+2yk2U/jVsLkGcpZ1n33LhL3zXDki5dmiBORp+iii869+o4nZKVO4F6+M
84bK2PnJ0u0e6Qq73pIB38VKlYeAjn2LdO7J2md/2wBOmxIcMKVqWhG1MiP4lB/L
rKvh8zZuHA0CpynFmdHLPez7ksO5s1bbxijQFpNPdxX6G+kivP1JU/eP8RgyoZpW
P4ir2xc9/lhRARMnoYb5ACOTHL+Sbet6el1WlUG5dt6s6A5YmFRv5t7Fo3bsX8tp
UdyWL536ENEJYX4hYcyGdQoauBOY5rcKon1YcDppU3rPENBw1sFV8BzO35EOh5Se
CCY4sfBpZigTzmFCIWpGR0yz68ui3ZomihD0nRQc6cbpAwksXLbhjVIrF1cYLL62
Gj7wVmyE5nZ7tPvteX4HCUvBNzyblnv17TfkZP3vnewAN94wiMX/vZGqHzTyD2C2
edSH6guRflS2d7ZvjJNLhP2+FbbKyXnXYQ82DD7szopBnqE5jCxUwHScejxh07cj
4CIrQ2/tJCES0H8Ugl08t161v3jocvi1J6vA4skQnn2Y0EwuoDe3aTIdgalRJJhU
omAH+uULD5lI3QxRqrSxTnIuejLwV+CD01I22QT3WbiKKreGJj6Aj3ZJsp1yNMXg
0aWYitEbsJ8fl5Wc8RiX2j0YDMb8A9Xi09hZyd4ZFsOJyBlDzvChI04PJZYdhbp8
xokKz/5L8kMhgG/q8dXz3qEYg7VwF5L3n5RBxOlHU1J6+e9CI4xeUnB9CRUlDxSW
rbUuDKVOUo9CQEIappohK/004SSfokGLTnWDRyM+9ZxUgNWBZtQkBKhT+umI1Mh2
RqOs6uLgjnIIRYHKw/rEgt84s4t1nN0S20jP8VcZHZ10Sv68eWIu3oKa75yFQDjc
O9bDcgDh/6dhCVF9fT9ZQtoOObaTeVzgSL1wdjSLdZe/mLMV3IE7BLyOAPErv8jA
Kr5bHRO29GTp5fqljGdO1zhcMySHu1QuaLtimUHNVPxv1HkgEb8lLHhhXATzRkp0
kQf0ZpefojnL+PXShgLaCfAFlQJNO/yV2u3X2wnCA4ZSX5Msxnxp6XGGbx83jYNA
0pMHYdvUjpPY7U4VJt5fjz5+tgtFcCXyak7XxrjbNpudefXRVWxkQNElaD/N66hW
/BOSkZuBeoQjlpsYDgjFeqdrQGAfugccZAPbqc/YU6asSJr8r23OaEurwVM9EcC3
kUlIqQcjw1ct1yKVt/CHOKRgTg6Dd/PEkZFS1+CGgszPpVV0/gPkY6yd/u4swx9o
weE0+fPAiT4hNvnZYQMrmaLOEaf6HzuHmKfNzTa9tHkDC6Np//XHUDo7UTeLvv28
rzR+xHb2r7t2lTRmFn1G3L/TPXvyDOHXLALet5ces9MnIKjPrBS9bP2oG1XgQ8UO
75YbEvNJrlW5bqBBcK2C6ASbL5J5NPeLknJY6cBkmQUEqT9C2NoukckeIBsEcygI
JoMRAhGfV8xJyRBXZ50/yZF/1Vm+sjQwYBRGBmmo4sv8uyT9Uad6U0xGsHSxWuxI
ZYUXnWkH5IzDo3e3wTXGd81GsynjTh1lMwDtGMrcqwN2OaZTNvhzkc4ijBrkUinu
ZXFTw8QlO9+0z7a+rP3G8GnrbLEFgMHfX3ywR46YG7ccORMe29DeLxZUAIMfEFfb
TUgRolprVSPAUYEGOvfyO4lU3NNc7eb2mdXhHo/lcx6z4twmAql57mk33qFhBBbh
lEOV8Sa63tAVI5v8NgHxGK/99caUhbLcYy7nl7PWQ4MU7yQ2wdV1xRdX6eKQVsXG
yjRJ6KreI4S+psUcoz969GHL44RdnDdJmCaRR6xNxbOyNGgrcoLaqtZ/aHx49TOU
AW36tnIm8bZlewttcbWKUsUHNBsmxKcOnUSJqDPF9PC5ZWASiGj86QD732sUzeRd
B1ujqXJoQvDSA7apf/AGFnG2Dwiewe0p97gv+fZ9bzqgqTFEeQnMJ+7fZJcDFBMh
nEQ1IGvfahoEp71piAG6QqTSZ9x93q4gAGkD8GXGp26iYKVl6NiyFWhxnWT2PumA
kTX77HnpypqpKCUaylnt8MttpKvdwTaPZl6hw4YKRyJ/YoKhyhq7CNN7bZoD0eod
I20xUNfKXvn8dptTFGJDhs7O+9zIdvHuqyDEGXk8WNfhF6gxjtM5tzZBYvKbZ4ov
8phuWbBGR56NZ15s7zroQBSLhVXr6V8o519YItInKoGa0Gu+dAFUzOgfrn8NlwbN
wfOZ1at74XJsqcCtYI61+Abnv4zWvdhgpjY6VRshCKuFrDCX7UIaKe9rMXazekH3
dpeRoipHowdrgWOB5Tp2bjDoY/TO/X7Pkxh4m4KGSLc0t8013/cHBmKPyGSNYP+Y
AFOOlQDpUA+jsN8251bqx5YAWY96B0dQVPE99MX1dGQd0bmwaPCplkc8JfcgCdb3
Nlt1lQR8ZvPjP6XGgw1Ge1xj56zdhv5PBHARC8rlf005tcGUOd8/FBkZ2j7L6ies
RGbExZwBrlJLtEyeR/cKaxRhNeSx9acpZeO1DBBXgvooqXgD3B+rgOz8hjiP7D0R
ssWHiPOlvRIPuT7um4D8nTDI8SLm3aMLd25ThZlxixCHJwCDCNcoL7QiRYQgmnTZ
vog3F2+gJ/RvUnG+FE+l9QZCDfiIjo1jXhvmESAzvKuehQyzZIu3yk0x0ejDvl1c
xymJNnn56ut0DpD6rm6Ohejl21+/6hWTpwshgOrSltsAmvNYHf1sEBqAn5UA/lkK
FXDyn7/mMhSCNvzHgNRoYccZBk3qEpGEohphqofAmjfs01CSBSfWYLJjpmThXr/N
s1wClkE+D4X4nwEszYcuCQoQcmW6HkML0euhduD4dd5cKIRFLBdo9SqjxDg22GO4
R7m/8RB4RemnHcIUSxmgSZ7LW75oFjw4IMMByrxGfJHINbVz/b5OovrvuIIadYXB
Mo6QLnX+IZS3nFogdiPjmSy6pL0NKFKBERsLuxrymT1NVo6yPGE8gXW7QsMyghP9
WBTC6umjcupdKoGyw1l16S4Vqxfphuityu5qLrUutVkG5Co/AES/OoPc8bz8JqEg
mNjFT0ep4xdClJdse3cgKnc7BPoR/BPFdqiVlFLCmj1lGJFamm7n3bDo8UM/daDF
Icna5yw1wYOZTum9j+oNYnjusrI9ZHJ9dpIrv9eTjo9TpYESOVbe7gWaHrY9QMFI
pFgllC/Z7vsjYjkyxOCk/MWcdIhnGDAVDTQ/y/zxa7/Xh4Vh3Lvoc796mOaGiEZV
RKbvrg6PO24eF1/XWnUIlIIlWzWZW6F9tjs0t1m2Lww2mG1oq4FTrfSWRS9QSYmn
HjB6lEroIMyGliQas4/oX7ksvyrcqTqGjD750G97FnbKpYfMKoRd8tzhSEJ0r1+r
eYcq7YKQfGx33APaPYXsj50fxW/prfYBucQNBT5AjhiQRZfA/gnFmm1NIr9fTVFu
RyBonv2Zuj4z1nWSOob7wR/QHsP2lmqfORUM9SDxikHsyPqRI6ogejjCUOpeCjXk
ikLP5XVaMfyZ2b/grWXCpW3Jvds3M3IMSyMlJmgZ4lZ1V3lOVUKAWubjx9+VEvzI
L2Y9PXDGpdp999OReOo2qI6Wiqh/yy90nhVhDB+449k4MD5snmx21OW3rqz2uCM0
LCYxdB3HAUCQYWEGpjBgGVHtlLjGShftuPJG/l0IMNzz75gO1h1WNm2bAvcf61q0
ke/2ix36CfndkwX3symsrETkI469x5sHXzKv+AVuuZlD1q5wPv/ObXEAWfmNlnzq
UQyzqfdEWRLfZWArImCZYh0+POnYhWXwd9ccWq8zZ6WW9p4tQTe97AnKp/SCF5Y/
Q9M7J3Qn42aOVPDd7QgrTRA6lSXxGa4vm6z+N3biwTDVROwiNZYUVYKkRYnOExGm
oComFLyyw/jVN01Z/GU0/kYQgX5syHfxeEdJnS5K2hiWXyeMDTM1+TGeAfAZ8Jjh
O3p0gkwus1jPBCOBAea43Us2ywKqnPla51sQLgqsskGP8liWk3k9gl+hQW4D0Ibn
6MkP7wQwqs2MbbNM1glkktYQo/Svzp2qDV9nZOfYCPFbNvcICeQBM3VW8L5Weq6i
WgNxrhnHv2wyhNio2TJo6vj7nIxB9mrpvdX7fC3rClT+7dlEmWs50WzuJLKI3T38
u6d39B8c8oPDUO/iJbSIvx2cmlAXt/+B4ca6EQyzBK4dCIXpXEB3KQ/x7z1Vq8X4
GlZyeoxs3OcKyIMFrv3SMEyeTicT5HfK8tOp5As2ojm0nZ0Uadn7EoCxrSeJ7gRY
VdhMFQU79n9na8QoK8LT4i0cuqg3KIVgSnzW1GV0Gd9VF3yNLSBbN9WrLYHUn0YB
tmqEtAuoZgrWetjT38knpUEUFgeRbSd+uT9v46K8nZYuYDE6uugG6KI1i4UGLPtg
Z6O7ON7eYc13WWDpZMpMQil/X3h1b5USgeNTlKA4gwd7L8VdXTkvb1yBHGTgERyu
NSll91KOIjqwf1QlbqdRUJVc3XtYt0LMCGTtzYNubbiLc8YR/zqhZF0SWnLMq2k5
KWRC80uiGPaqT8GIVysOJAno3Ot5FBQbEyNWdT/hZduDZNmtflVi6L581TbDJKpH
9vur5LdkJppQGJ1jDKndXcqth3MG5xaj1z4AA0Uv+0iUjhuP5zidDsLUAEUWk6do
wwMQ/hm+4Fq/GMXFqfCLORgUXzTu31HNRDYU4HAnLWtrsBfLEMPZnw1wq1wykaB8
SNTWqpAddAKI7YicefPJNM5A3MLcmQ6qe+5XR/mLHU5/6wbZ7/zklnQ3WmhnhfAA
yVKHwynICBxv5HiyAwFZZwobDC+bGFjBoWaRjFk+CSNbgG/OQQbu1jBprqvac1ee
c0SbEZseidMaIXEhSk0mnPWbWrtj4225OT1zeWVWNSoqFU7Y7+IuUCG573KRaBjY
BUIdhdRqY+1ju8xdZnfz8WL7KVm+eexDx4ZhwL7xdbICWr89wc+JkEdgMLZvdJkd
DBvc6WF7bFjTkHTbZuKy4DSgEi7aaiLe+oNppYMy7ij48mnL/DmFae2QY1kJP5Qq
oB+FX9EQaATqX47YUoJUpJ9TUtKZjrJBC4i5oeB6UPaw6rAaxld86cM2lA+dTMpZ
e/xkuKagjQEBEA6GUq4E3nBACgWUMxGsWE8ihjaDWQFh7OePIhm+RuZNoU9vsht3
/aAmLs7ygDYDEoYjKM0IU/AoNc73XzQyRBuge2atkBYwKgp688Q0kjRTnoSEp3ti
2dI8CGPHYqiioZ/ZQJZbffJIW+z6p0ERdSPOwwxn9QNRDIFcrb0WO5/IuxYl09eS
HzXwnQTnS8YvOkz+3ntZ7M2hGLv+7wVTJNnRmcWSBjdKmlCfDIuSvkTNMH8lpnt1
OOrimPwO943JL8eabu/6iNfeBujNT8iOVHlQCUNdLJQaif+QqR7g4Zz5e07352pQ
FPzf9YSoFhwAPmTq4YVvDjF3qxztVQbBvKit4mtBbj942uqYUcECzlS2/oRejDPI
BpXVfDrth04G7xwuFrvDttbgbZpvXadrfkSHnmgmY9JRgVwcxk/HMh8ls68wIL+8
+Ixfyr7VKLPM9rvEuft82mn5nXt0KO3yV/h/EbOmQbjPAqiF/1YCkOhvI1OR8d1w
inh4tJCuHqdgPFXlL2GSfwGrQP0m2kyDKT0KydausgN09tylwdunBJIW/f8EQ7Kl
MkBnjIE3GcE8eA7Wf+0qr3koPYrNJteDd1u61ACYm8CZkkZv6S3GSVMRI86weVNT
jBx1ZUh8FRIepBVpAmsUOIT2ANN55IvHFfHrpOqccuPlCdfbKDJgZ/4FEGECMafD
0cwhd06lebJlvX2rvsIXkX27cdyvyviNhpKJR4RmybEZw2HXZOYBZVKiPXimaBwI
YZ2bf/hG2U7OKHFFxTKWfKUxdBAY9b6LrR6JLAzE62ZFLl5iEhT+kAfSsHLzwLWA
50kIziBMDwN6V0IR3PSQP63VQYJux1vKnaC8GsRSiFPC8Ue5YerAfQVqlzL8SMj0
l19cD7akMjSJWG5lmQh/YsFK3eUXrzHCEb60NxRXnxG+RaKzx4QbkeU4wlE2Up02
umLzHWkzhmleiq6tKWSjSdB8jdYPK0L8H7gq5CSD5yON1vuCTLKx8n2xRZ7I2Ocl
3m2slQW/a8UNSe+DgR41WmmJKJLmiWqrR8dvsFidolenWx8lKtgKx9lb/0SLsdR5
qpUk5Fv1SQfGx8vRmnYE9DI99Bc8DorGGTkvc7zDK8Op9Lm98rcPheiJL01BaHvN
oGNiozaA4goEEKZuOecCilGQNV8tQ8mYlUQnzL1j0rt/V0Q01LTBO+ksRySh1NkC
yxuRvTdrogAdjXh+8jkpZDl6tJs+xYceE4pSoLnjuUs1REPB5cFa0WZ9xbOq2R8o
uTZ5SVEFB42rVGvFEoMOmIOLUG5gJkiqyzt0vRl/jndNSfGNpMrdHBKhEJC4binE
OADJEQl/GJ0oA5qinhX6ITF4z6VN6h/v51K1gmtyPRK9Q0+exgf5qGVqwzjk5dDD
RZdlWrP27dxvgO5c2Txoy+WrwFjHkfd2+hA4WfmMZwsVT3/MhFFC6gU+RaiCoIaw
iSnk8kBAYaznwi+DSipxHLyxoZ4jsWJt1QHALHsH4hHhDxqYVxIhwjXusfq4ayem
tbky7jdfUWbbwA29+jaIZzGXZJ2pzLRoU2616MgX2tYJbX4UG1yWT0uh+XG3AM00
SBPDrL5sfMWym4SdNphQkadlSxNmP8zTh7GOTeqHBA6N3GZWqmY+vCtZ1Nnjybys
V/2X0fzswsPsKD6KGO6mUjPv8ZO1Psm4inRLxOzPFzs13BNxSF/xEWhfM9hwRs3x
YfOYaBrqNlvS46yReK7mZLNa8BNhiEOf1kE0LV2CeDB56J6eOEpX2CtRIm/igsBl
zZKYrU2zbqONxLddEeT6t4aDHfuvyr6ueFrEVH7UzE8sno4US+8l0H2rH0/Jvw9Y
OCCdNnz8gaiBBDF/mRvFdltFo3xdiwIMBe24sL4kVatuDwHR+tQ+/u7w9dgOky5n
la5AIk1w0UT/x6kyFm9R7bzTUyMMt9E+dbPW7eeuaCJS/AwbOW/dcSQcLNLDMygw
pRO4gwny/ZFHlQ836IJJ82e4DfkBPa7YdiH+Kt/E6c/hiLpUj8N2T+zR/kpF1/rN
sbm5tAQAzqLa+uUDll3E3iKX+bjISRxwL4LlfMrHFIgMmuszbJi3C5PYfZ3jnUmS
/9qX7vzmLJuTUgu/QO8bdkE2kVdCLmLMefIb6zQCgJB7dA1JzkmX9sDQ1fFgPyfr
un7C1Yi+5KPYK82PwIUgaespw7CGgDJaSnpo8cBJctBSol0p6CVuLK5wEHqoOw2b
aGVRrNweJ1p+31rGZot3BDKeTUskODNdhFmmUFXm95KPOdWAs6KmDJBdCkXnsSiO
8QqPPae7AGOjKbwfhKt2l39wHsAYu69paVVUxd9AodNMkJ4+fqejx4pDpLKbgE4G
q3X5Mk8I1zf8W69GH+BLmCRlU5R5xlILefWkiieJlwFgrykHkueGYZ/BEzG6fkvu
hoged090prcg7VIBQeOGPnecyhU23VK3+YLeFHB9/rxcCmGudcLPsXl473Y5VVtq
02/uYXNJbg6DRNL2vB/cGSvJVMpcE7QuyNuC9V/kDOFAqyEvLEuF2Vs5qk3vVlyS
BjbL9tcbKuOapGZc2vyXxoHf/30C0naVQxvb8MyCRZLzxVQmig587mIigfTpZoP7
0XW/65kWS6GzsZXsl6POKRMkBckMZfIju8Qkx0bt3J2RJ1gbtq009Z6VkW+eY9gY
Ghf+HdU50rl/nUmblQK/RD4bFtJ/P6kVptngwVxAf7Hokr2MkOxZ4WZ68fQecKxI
JPnDda0eZ27VkxEjooRhhGNTaPGMquyZ2tex1I9FyIQuV6E0jl8Bf+Zz1HOMjqVa
an189DyNEX00T0uX7BKc5KR2a3mbcVmyFmQwHX/ekZMsiW5jsoK8nshL1fK2ISCn
D4SvDkRgJyIRxg8GAJ2qegClskP2LIDUpNuuu4n8gT7DzwWaiMmo0vczXWeKw1g+
9UiF6rNKn74m3euTbAsNEX0o2RLFZ9MDR0eWmnW4WT6VNYTH6c6DyG9fbOBtq6GD
6/e5+x76js+yAZeDYWEFoKKOuq1xX6D3s9T2KlmisRebnWEDeS/4s+2BEB8oIyCr
q7ORg7f3ZAbDsk0eaN4EOMGExnjNwN2oG9I7f6y6T4AmEu8Q/0WhtlBqT2TG8ZFa
fIaSKGJDshVEqCPrfJTh7Gwxv+v4/kois1Gsics/ouDACyXiYH+slISOUCxLYEYi
gzBFyqYt3CHZtkF3WeL69PmmNVojwKX37DVFD9Cy9rUVhH7UzIKFtT/QiICOIr+v
rMhKUPcJ/M3kVA4+RhcRf5yG3rYueAWmXsYxjO7G+0dLVI0QFLPv8JR5qWzgXX9V
ywYubDtbzjf6qmmhT4KEMSebaH1UiZRnif+jhJYheusXmYvwOeaZnX2u/R0peEgn
uGDwwLcI/gRMj9HbMBzKkpFjEbprOXG8fG/jmRKweNDxZpQ1tMfn99biAD1hndWt
szy3d6jEjKwlHlQS2TLbBvdhNLyQ91WlOl7r2ObfKPFvG+BqZL4l66003lHd9gbE
xbv8zhVxf09Os0+T17HmyJr4DN9jW042ufmEsD/9OOk+Hnf2gvky0EHNzz3l+hvD
3GriQu6obbS4wBrnSozhq1PCsC0LUGavBh1FVEXCLRNyJITWnWsLcoVYFifrwySB
GeuHtNESm5i11zn4Hsikkb6+k68O8Qn66XLkbMjuJ5I0k//MwgPyI/MiAOGahjpv
qPYGJLig2xBWUwch4NI9QTTTFNZDW9iXjJqBW+/1p/UXt6h/7J8AckaERT1NDDPa
ljLYgRyuFy8DTeNQVDH9INB9uIahVcDyeNDrqzyzd8mNGQm4tCcfJfhgmREL570i
RwjcndKO2ANhYbgjL+ZyhUOdAicvdNQxpIOG3EQgVaXAwk3UmRFotkejC/q7JV3P
Ip0AiDkj9EyXeomKaPaBNC1FohtfFux28UPGvc5t1S1UmQ5avk85FfJUWvfaY7fQ
CsXYD8Rksg1JYW/pj9v8S4Ep5XaOINd7kXLtQn82R/VIsI9FTzCPlUNnshc2Tvar
0NZ4d9IS/MHFW7WpuaSSIy3hHNzGDv0DXO6WcDA4ek09KhDPWSyPmU0FkvWd37kC
kgfzSfS4ihPbKUEvK1ZLRtnkQi9txlM47sj13h01KyiH6j+aJQ8KybWbc4nKZ+jR
UaPFBh/p3RbL/B7Jp+k300cXIqaOz5xQ6dik0w2cw8WduBs3NdwEUMmXa9JCajtl
IFc3WEzyC8BaPnSKFmOOWoy83Zf5I9eaMTt712+1gWR15MscozYYYKQ55sHDZhiG
8nrfl7ms64cVMwRYatDndhcgYiY0wTtllE7cjly49UqB/hhOWH6G5UZbG1CsxmgL
tTTzYkrXLrn+sBgIJzJ6jO3gu2kfDsCVzCs5I+/ODrgmx1ZlEYm5C0/B0hEiG7zU
QazpBnoo7Ylsi4h04xngToh87eaIX0QVl/c97K0XI/YhkpFI9whV/jv8nzIFfbiP
Sxy65z7JmtRuHGzm6AIUH/ap49hFlVtMY8EzEHzwWBt9VoyzYyKGfhwq7c2Lbx9g
o8YRZwtGPMnY0B6I9viMvgwRNJSYeRO1/UxwVYQRjb3ABvJTy73KlSs7Iz0IpHDl
Nihd9zpv3iiMyXf+fHsce+T0I9yfUCQ+9XsWl+CUM4xJnTE6J2+apzNV/XA7uEGJ
TbnYVTJonNkXYLpy1zUdexXeOxVCYzaf2S8MJxQFhs5X0mB1Qv7+huqbe9J7xvSD
Bw9zGN1O/1cA1tLM0nfjJBc7aeYLBsaT2+ZUmAUaNPPpRNI9ga9dy1JpYbvJt4n3
w47IJYRheK2g8TEQNgr1UsbpKQhUKKObHyWiUxVCdZEld61yQ+A652ATA+mZaP8K
YiFCs62/kA6mCTl6hzPkkTmzYRwjAzEroeslVs8vRWQvt1LiWNviqbyLs76ZCOdr
4ZS12zVZ768qc2LgQaqFoEoOujWMQjHxrTC56SGYrbRWOLriLSGmf2ZwI6EbRpMf
iM+v1AmcvuH3VHFj7IGTvUe5rlwQDjsYkmA4ug5KBwpOJ1baYX1+1XRfseDsnt3m
V76oL8HQppbsXNgkxsOR7r+9XmIiUwgWPvUufxy6z1MD5ZY0rCCG93e1QdTrkqSp
9nanyWZfrfouV7R07VjVPvIhLoLWv2q7q0x0l8TnpuiFMBlP2SkAGwUL/VD0YgW7
BZo/+DyvaCcYQR1I0MpBQTT/S+hMF48Em/HOT8quHga4fL9iNZ6BL+0flnHFltwO
ynD4mI6j5uk69lASqAmsOsJU8Pcs+twjID39JF2gjZlVimDCnSAj7KUp5IMjy1WV
frcEQlPj1fDVx57bk/copH3qCGEGT9EXKlg/Ocg3lBGyEvOsTd7SdubxBcu0xnds
/TYJI7lmFvVoVljvyYpcF8bsmjlXqx+TDB88iVB97cbVqhh78+xTxV63tR5d2zjM
GskwWgOXd4KYbX9FG3wNZ/3uAMKVEhWOuhLNVjsslLjqv2Ytz80moJKZKcriWdhh
/eFiYBRh27u50COnafghKbQaXz9ZQJpphDAHgi1mNbyuEln2wSI315tuHGFp+q5/
ogApdw+/YDymjNvk1k3GNzo3vFyOfvESwjSROzzJYL8p520yXKFVUa1ptuMEieUM
CJJ7A9Sb+fF+u3T8zBor9YbuaF5yO8PI34s+kUscvhJP3e6T360g/NDtu+OvuRkF
vaC9Hg3Q9yUf6aVxAgKC86yEJrt1PTmRImI1m5ku1wIRmW63dhdMOvZJiex3MOgF
JeYX4Wdu3hUI7cSmR3b45QCvfgBWGtV07OMjD8TB3ChXYy/bjd4T6t+e+eIJ8SB4
0MMZDXFYchE95M/zCCspXtdEJ7GA91G+m5AeZ2GxiaKYRgVORDKbXygIAdHmkS4b
WiSYiUaheXSHeIzE8bZfcna0DB4S49MSkcxpLq9kdMG3i/Fr5JvSQph/e/1mkTCF
MJzhPzLCLOIBa2tfzreF10b99A3h4tqYUksN7y59+Bq0AsZQSE40Of3sksjwtneN
+KLRBWSQq/H2bMOCcL4Nib5Aap1nHwQyOR/ssVhhMf/BUwUcOb55BPljIWotmsU0
mfJKLO9HLHzMqKHZF1UKH25Zk/g1C1zS+x4SeRRsgyKY5C1OcJssQeo5ppBxohFi
MRAd/SYH9dxe/cDUX0IQOJvucWxYUJ94pG3cds+J6P1B1l2WuMA7C/RRMJm6cA9I
x+bpoIbcYHa39NaIUvzsJugpnfo5P7ipkj5EInDn+p7jIagswAQJOpHJZtoDCEH9
y4VSlDGHUAYqmO4bFt2CvYWuPMzsY5SyPldKflgRLFY8CPHt1ukIkN35lqhMxNeo
PqyDiVO83T662bRLdDO96zQVwSVdh/mpJqTfrH94JkSHBzE9GYhcJuU/+4+AFMlT
+fTTDKebiIvWXK6GIBnZzPeGfV8z2gxtCA424kwjau10YQq74TLiqs1IQ2C3NNtk
VFLqgtoTrOSeYyxir8Phz4OQVUI4qspZpCOeeIrMorkDQNzic4DcviKiXBtYcCzd
2muA4aTXURIhLoe5Qn2Y8ythpl6BxIaggeEkrMb3aRTUSxOb+Vy5StKvSSwTQSvv
gnSGpadYgebh/PYAvkT4OjGpBcSgmrSj4j+GykVg7zkX9RHARkOriZ8Mi4SmuxWW
XTDKTE6MH/4kymMLSx45AxKe5MT41KXl1SW8pFZmWUBcbTs3xV1TiHCGnF8O/cM8
fSgSr8NgUBBfYeYZo001XwpdHBHjU/bGYz7i+oH8dW4UidpbnctuG3AkonfBqeWr
GrhNxQvXuFp9HD1VcqIrGy2jVLk12vnJ30g6auxcgkfifmszMeoSLB6tw12gFCvP
teKDLMSCHHwmuLU/OOXY8zFyQwqFKy7M8YSMfXfT6/zuuLTXgMX2UsMMtb/b3T2j
ShkdishQn/JVEBKkvWuLD43KhqMQjFYfQF2WgwlOV+X61rkDVtlPgpRnhya8mXT1
qcidQxdp6qyvRq0WAd8DR7tH0LT34VxNamIMf/k8R4elNDL8Cia67ktS1I0Qw5Pj
ZygTnySJACzbBRLRE9T6ZjsClzLX6P1AEOz3LkMDn8ycTZAyTV+9wFwcKrHtnld1
VVg0MGn6F1yd3KJtmzIFZ5Ma0XenGFgVYpOy8eltPEzTgoNMPVhX1YN8QjadnG52
vRkfREe84mqUp4bmfRQLj1RyAvwlqKRvWt5rAXTMNhFUx9i7/jt180jQq3lYts1x
6zpRi19X4DJ+5oY100EQsJLAmP8BBl/fTuPYrR4PXlivziSleitFWFHwnDBpiVsu
pHKsv8BYyqyKsoCf9xOPH5YtI+ssfQcKQgM5HYQSv+T49f6kQ2qA7o+swBL7pfWo
vIOKtus8pNg2sh5Rf1PuVZhm6yCFNuukuYcP6wzh6HSx5QWo33YO3dfDqMpg2WYn
crSGC55/yVjpMK55cEC9iUAb38z5iZDSpCI9fhJFA9PaYIjs8IfMsUkEkxrXLjXK
KZA5lE0+yN0DfyPV+7YA9npLGEdmlHoBwWJ8FoB/Gp7Frz0l9uS+LPUvnjvKSoLk
eNqMI+mZSOJ7Yjrkgos8hSa3G0pqk+sA1XdW0h3rf/+o+lA0WN9lhDaUXascBG+t
RTUNsz0MnuFR7Qnu8k3jkxgknPd4DgXQSaI8RSFbzSXylbRDj/3sMWZf2qWptzvl
HPhDMn7tuhqohtLp9l+3GzgheW9DxSX/+s7xRfQ9wf5VIfM50LuRj6uZCCOD9jSQ
d0nYp0PvLQABUU8dt+V8TQilJn67hV4Kp8spyybwh1K/EXrDEjAtzRqr3OHpP6hD
82T1pjG8tK14NOp/YoKH6jF5PWZZxrt9YfyWYLkSApoCFEGn76efVR/GeKcLwtHx
jFuD4QAvToc818FcMjWkvyhiHkyr/YYrq4HSOtRtC2Mu2uFsNOTywQ+25aw+kfbm
4LkEbpUHySiPItAkrJq3SFGIAkDsr82cVAkGa+cmaQf+LjzlyKJ5+FhjyMJ4wcFs
zj6gLpN49rd7G7gpaxTR34GGIDlaWI+CbcWJXT1y3zZZN2db/8QOhjwDRMYwZkJv
6ihskC7ctquINvxrJKMvvQO7SsMcns0B0Sfv0VPhegV6zEd5whsYzTY5wHSyPUT1
KGLMjONDrdkaYGuu6uOKxxoB3e4nf3xor6+oLhrXJ6TwxQIW3dik0PIqkwyYBpk9
Ae0e2XRaoWmDOHhuT32mG9mxjwEfVOpG3Nzor7yU/RK7xxHZ4TbsUvnTpnORWh8N
UdmmJAU8lvW2+m7h9EiWwTbl8lQuiww5SkXxQCrC4o0Wh1Z7Qy+XmKoL+FjhsyUD
WN97d5dW+z4u6JhT2dIbLHi0+d8VR+UbpH43ZZLcR2tKbKNTzq7aCrbkapO29jQZ
WltcHNO/nxgN2As56cPDT0LZEqhEVkbW1y0Mt2T4imsPN+4rW4tE8ngbZ9jglPyZ
X4iAjyad08dLVyMkumgmxS85tEX1K2XztJZ4a/qnHpaCbTJpye9auNJGttHhxRQf
DKEcm5IwXEndHXi6fSE+LaU4f+CGc9ZuIt0nnfqYF+lzSEFoGXtNbFamSlw4Itvu
XTAzfDSxBb0pihWVUAbYGlj5Ecu6CEGyK4IAjO27KcIfbvCW8fG+9QJRWfTZjIrC
oTPvDn7W8M023aZzspoG/CD05Ho4Q4/ZmfhMSPJ/+IQuey33iN4ZmCpcMPEqtfao
K0AGllR17dU5QtIekT7sGyQtQaD/nGHzCOAvZqV6/RWXpMvdxlbNMTaXCRVMxxIy
3KQfzKGjravOfJxNYf8uWdkTO6zF+yj5CYnVcUDBeQo0YmiNQHNRGx8rBidiaUWO
caZnsuzuiYdno9gaCyDbbRLGWhHIjMzjC+qmGBXqvqHSo7H3x0doz7CRroU2fi5Y
LdxWfJIJYr9d3i+j8BOrjsYULMEsCacPAoEpeWTQv3iSnqZHwVguEsfSrGWr09eP
M8sCPntqhQYuGophsr5QqGMahz4R+QufpGUjHo4E7CAhE3BTiT7hEvesItxy+WcZ
9hLeQvNdzZoMj0LWgUENMHh57RehnAM6IbSWMDegBP/EEbhpWGqEIydFob4Hxsz/
ihv0PRkGUtzpc6DokMhn43rn9B7+PXEIuu2DiXrFX6PfxMJ3DV47oQj4AuQIBoJl
Ak6zIOvygGrX71bP7rgFD6gdlKH2my//NfiPZuS6Bxa9JO3MPKorrN9YsKrAfjzC
ryx4o+YuFemnf3ZUDubBrXs8AGsW2PACiSLFaGP4BvulQaNur+T3fR5H+PV9FlUm
86mTksxIbhRSR7u56kXtyjodY5spjExkg0stav7v9qdsBCmzQ6wdYXkquZ1ExRis
xsdvENzIrC0LbEaO2kq1x9irDvg8nJy6Vz7Ew57zn5mjoZyNjIVV11uZtcGtugXj
q8vYtEZcxbeHwlzdQZhNyJub1pNw2VwkW2ZwrxQ7XVuyRzS375cehJ8FZ662eg6k
zyfDCrrRsvUfl16fjGOiAY0xS1VNuljbzUxaq+TRcZPBhk4RpankmeMPpliunZ46
EmQm5k9A28x0kCeFrvQU5CSyft9mMCAnaW5ENRWigH8mTPDSm/8xsmZSdsRkxQIV
YC7PUI2dTgu/yhDXAV8dHV00/aNcNaPT461NIYfm0S0WWnOqTP5wZayd8kUJ5SzA
F0Ujpzrr/RzjDEBJCfIdwjENjOsrV8/XDNKEmCC8xm7MVyLaGt2oQnSIzqOphwU9
cDGwqZkodacqEIF0JxPKmLNZ4ofuNcxzy7jwRPEMpI9++0UdFeiVFHTHENHYvI6B
ale3dAI25blGcgy2/2FBclX2ukE8RtiBTmwFb/8QBj3T9xHukFcZbBJw1orHjVIx
UBMQES8K+FwNAMJZmubFJn87Uc5gEDPCdKWT0dSpF+Oe42VEDGLls3BL+PxTGysC
XGB0n7nm0ybt5ehfGm48R2h83rFqOgd+oJXBEcrPRDnkNU0QTuHffTl4LxrCaMlV
TLfTplPKaEWYS59CiHz4xsFBgEdPW44yWcmq/yjYkYaCE+72hcGrxi8v8PDGuXqp
KnSxO0nIhk0rfq5lfECQVtHbvpZehffVErgzlNoag5HPVJIC3zMx9vBYCvvFg19Q
rDlBnTFpv5dvCOn/YNHwqRC2Nf6KnkRKil1YEqLL11Y8gSPuWxTJ6ihOiJobs/o1
yRuOWR8AYdxwH3uPqQWB/MEBS+Y8gNsdWoTxy7f/vo3svJ0bKFqB4rCkuw7MesC4
Aw5Va02GocyHJ+9Y0YfrGZVmhC6gQo9hKfxUOozdaiZeeBQqo6pMoJcsnli7D9g4
toPIwvrRJ9ANefSx0lWJEcPDeDIbQQUv8i5Z73SDLpFrfJ7HBBRZZ8K7WnYtYCy5
KsrvDn5czLSv1hMzshcPPNIbjOf0UrBEzDHJep5+WrlPpor4WiRxN+ap5Iro/yO9
8I5tuBsknBj60bCLOdidgZyT5JD5OMlr2u06WJmEshAvHoEAVJ8ObUiXguM0KWmZ
2X7a8KfRsHIklMNqYs6CK4332mUITi90YNrsMC9scBhixfPetCDXBpqjxWSHXQNo
r9guxpykrb9UwuTW66dotUBnruUyvjeT+kiFxLT2Y+YOLoMnaQlBKqVWtASPuBN7
FJBEm8g/jCb/is/GKeb3ACQvZtPqi+zHP0EA2RVNCxBlfPor4nFt6a01Ut9ERxfr
5dMB2wTI42/oKPItaEb4sBpuRq2YNauy6XWPZxLd1u2PBQinTeIxiafP4ef7Y8n1
5CFS5jOVyBBf7CaIc2HEh2EZk4iUnRoz65B8VmdXXUv/cAXSM7UzKnAvedPfokLS
9LhNy09mbI5+pEXNF+XezMlx/I+dblJoaUd9wL/z9zeXp44cedAHyN0jq/XkWdtD
CqTDR2h4g2ZbaMIsSbL1uY0X5d0nudd+qjTCe9C2bp+v2EkmeqmQgSLGu9YdF2ub
SApAm1ht8535CtzIOoXcqT5q4U2UbE6ZcB/+YL/AqUAA50MdZDwvS6lKtCfkAZJ3
KPZmRu78n5P0lgDtq04RZevXWbPWAxGElv3EHszKzlpsJmHOdncsBuh4Xu9z8k2H
tC6Aid8GvLKxUJ5TygEbOXbHBI1JDoPzARYVqMZbATDJSIAADU1qKuRZM4Kn6mwF
Lf+bFNEs/WpAbPhKAhKtuYyG1Mp61HXnIlme97+fGX1x9IMhImtzaT89888BGlv4
0MT6Owr0Ov70rUAOwFM0ycyw/+BuHA5LTsKyOHxjstoRczfMms/SB84Ii/cNyL3/
YJwh98geuIj1wbUAt6HU4OLe92oJI5d5CguVsb6460mvx/ajyEmMrSxpgtKUZ2N2
InIncwcKoXlbAhyluoYgHBvnmldX6YCz0caFKZubc5dPPc6Oshf3JPX34f1z9+L4
ufv4/nC+bYqpm+09emUItTOnYRed1W3QDxTGFk9xdN43BJri5vMMG75lBom4dM3a
3RBDwimGaUF6aFOpRFawRVXg+QKNeq1cEMpPRlfWfgC88z5iNy9dLbq4TouqQp1r
51sIRp6xoVSaK8i8LWcnTCU5M6BQb3GG5ZQzeYclNbTdhMw8C+u+0jvl5SZIalO3
3RMCRQQycfWUw/Q7Yb4eUKxbe5C3iddLhNHqFaM81LgIPFPB8iRygqP+gPTP9huH
OQXwkNKMmqvjkXcVxCU0bSW/xH3N30hzrYMnsR/F2LLb8h1ctYrwddQIS7B9tHzH
oVbYPSTR6wczcNOW6cljV2JvBMb/eZTMV8wlfz1iTsPmE124EIOnhd5O077ucHLz
CNa6m6hX5HBJ8COnm8tJ/Q5SjLBkXCmTgavHRXsTJHnrNqyA71UXdzPKJZHxkqn2
9TsV0jMlbClV3dwtN6UYd9R2zjDS44DhPVSdcrBQMPsyWp+Z9U3prN+SBrEnrVh8
Ct0SbBIA0ad2yBTwzgA7RpQP4Fk+AEOK68YSB5uTYLoqdGqhPlxbHThDkrGdWg7n
Rq3MkB4+y0wRXqMlwD66JYN8y/Z3YijSW8bpEYwlsX05/ji0u6LnzV2QVfdmfr3W
QcfPKSYbdG8SapS1SEEn9RmuY2n2Y61CRkLHf7mp/b66ex4pP7AyzUQ5PgPvO3Xm
Qh1agqiowmbaeiwTfFk4vCBOmgXfKN38U2hdd8E0tr1ffBIlGT1ZfemkT7es0YHv
IUTfzN6ByaSvJV761gKY38YfUs3kwdEy+mtofwwm0coLZz/N9buoyvdA9YIoOg3B
WT9wk+6wnD56I5upjmXN15MJnQ2C0dycs1dQQUyMd80KYznCl2hqrra7HwxAhPfI
UL/U6lGDogumAX7Y7d8wXi/3F/amGsdIRyzrKlD/NY+DHBcA4JfNblr9enyF/QYA
hluE9d1o1LZibito2KJHodX1plIEw+eXZ/FxF1oiXLYvp0nhCd8CRGZ+rkzt2+rX
7s1Cwm9CzyyASF6g5EemiVoF022ShSuYUFWgP+QvjD7Apfx2yC3ijRtyvBAYDNgv
TbmYeNNiyiqDJ0abnjZcm5GN564rmdtMY15GOTobsAxsirE7i9l8gbHWSJwsz5ud
5bJiRFFphyzZEpC0mZHa47AMDOvYY6969+PodzBsOiGdQhcXzR3cm3hcGQV687hJ
N2FmpEMUfnihOmlZGeGjEc+9t0nslo7vQ2y8YVCvB2d2tFDnc+oMzZWXY9iQp6Ek
xURr5ZvSiO6H6W0khWtJWXDyk8ZD+lmzPB+TYaqdLFTzxFRHV2QW/FpJQu9mKlGI
75YbdOsxZlvyyR6UPuJN81tzE3eFVk4lYbCULwUVVzedxh4ViMThszbOxSECOS1V
ipgNhKNP8BoDQtNKFYzkIC3xd8niOZKM1zsTlcova6QSMnE6OjVt11/1G7CoyzRO
qJ7uxGGcj5O1ajimQ0LSm1W7Ab9ghqaI+8nKGybmmQ1buYw7Bzay14V0VF+VWuP4
ZOqZ6tbgMgfMD4oTM/q7KPBMRyduNDsW+aeJ38SnwSzr1PnpXekngJf/6OHNq3pg
4eQO+u4WszdmLqRTSpSyXXpCZCcj7nAh1lzAb4iuM42+MMnwsCqxCAd2wAE4HMqt
MbeKGgYKUNcGROL1xleeiSJxwtA44boaFIo3s6amolxhtjrnfQJOMft3tuKePIaz
HAI1IV23Eo88Uwm0bZQcQ2z6bYs1wAR6HWFWfs5P5XvlaWCrsukc/HkgnLmx+2tA
UUUh5yvPmoJ4pjPLHA0SKXyMcyrxUeW/HVF9ANdRX9lqKbnIxo++MnWumwB8LvAv
pjpWdxBJ5XoVmwSc5A1dK3JblIUzjtt/4qU5h/r0I+9uRK8/TNH1T+MUe41KXEEr
H6ymbqiWV42krUI6Abhru2lU6//2HJ47ZM4uudA8x3ZSRyQgfPX4ryXpJYP0kEdY
WJivRrMxFT5w6d5mKR+qA6a8h06wUUw9GcQmiZnp2zsoM2aGjwf+7/ycPvVQV5qz
spDHR3y+r++hd0d5Z0Wa+a9CM1Pot8bZnfB9Qw79wKKkATYgF9iHn0/0sr0lWETX
6zRJqZrHQ8cprjQh8SH9QhLWPZuZ/LzdVB3DBujWfnRSSna0z/qMkNM/jfkYHy01
8cDfCVjKJcIKsKMpnoPVitLXotkn/A7veXioXxesgvNBpSwv1MHNBLg1ipQL6xaF
WP8jICbvbYAmolzDCwLxeTKCzyT72B1dTRmLJwQ49IfuGgFYyNGRiDUhmwMo5Vdk
96Cpz24M1ccCw3dDCNWhbRn/GbYA5FT+jWILHtEfVk/gGMZ5ImJvY7zBQ26bdOBD
vUSHfgX9BmyHYpYRghpjsm/HTWZlECPs6Oy4aN/xhp16Du6XfAUtQv4Pp1JT1461
VfUa5iyxNwlwIM0PGSk3qstivcUr7Al5DEHbBIWfAf89fjsHFFJ8rZW8pDJulb49
AF42+zXSMx4SRY9OqfQs6pl32Wnk269niG+rJJPseGl8WI+OlGzVI09a9C0bV0JZ
qt6up7OGbiAZjSpnlYuZyN8lqvrm+fiIJvN7JC7UK131Ax6QjqHjsj9zn8m6N84z
V8YIas+8AYsbQZtcxEV+ajQgCxN08tESf9CjWIy9sRJPA3l8Cm1v0EASR21nCffE
Gr76OViLI3G64rMPUJu4A4KHo87S/9zTcVq9nf7LrTIljGUOxtZsdXuHXM/Wc2wF
e7Qe3i0zEB0KCDJE7Te3uxDMNWcwPOmOVuubrwRpcXNyJYculwxcZIBPgw1jGPwd
ZmzS7i1dCKq+JCH638hIYwtHhqd/dzkLnZRnRCF8lkdiQ3r5PThaWNLqVMlkYFQn
Skyhu+6XOPFFFNQ4pgELwIqlyHeX+BZmgPLRvOl4aEUY7YLq0FxnXCKthpmJ0bjg
y1hMN/ts8Wk5EbDZg2aew/g7MyGXtHjItCXy3hSCpSqC8Vptg8nlXgKDVQaK+u2r
joyvNvKFx50UE4kVQpVDveUulQ4N5pOGOAuAG4/naihitcc4uR79MKnwOrGJ8IqH
j+fL5rFF0HfU6wsrDhv3WKiKJGEXoI0urol9v+OR79/M+/Um9It6FihZJQPjljtS
MJ0W09du8451ZG4ohLaWcOdVGQELMLJFClkw6E0PBnZf5Zb0K7SVN2hstEvXvIty
/VAtd4O1DHgYUucCUFDXTOlzAcF3ZIGM+StO7JLeoBIwsDjVFbjn0sN7s+QeB3GT
5R039vmXavYbfLvu0Zg/7NPxmXdYsI/3NZmCsbiDddQ1bYoyF1Xk1r+Sjkyt94Hs
loEWFge9P1vYyZgWJtkIl76i/n7DjWkWZz1dmlV3CrUYBzIa0jHFt4GC6vw+Ecx3
axPjZ1Fsc0gojqyWJefTRkDEaWrKxP8aiYEMnZblCdnQ/12iJOpP9KdLRwzpOeod
3yk8sY1N41sukzUygnLBozICtVcZ9b2+ZdALyXalKqKz0SVDQs17iOddXqvlgfTY
4sA85wpW9fjRiowGvkt+EQMocn0pD2zWDf1aCuqBF/8/YubULJswwwVgYYQirZsT
+zDAQYU5qUnlWfK3k/UcFmFFSeXK1C8awTwKu71gRT6zxW9uDWNTSRZX9ksH99s5
ziZJ7UXGwA9A4ysrffkw0ylKmfPtlviF+YTLCBFUw5FEmsnq99M8zaFia9GHOTRl
Rl9XYyQ55i9OmLoh6QO+/2QwBRJ8Hq3mKV+IX0xzWgR/8VC9KFPfuz7G2XAOw1DV
/0kTGE6HJiJqFS75HpREP+WZ+VB+IYJ3/foi4oZ8yinlp/WGqb1RdXumC3mEs1iH
ggzWa4tU2wPSCNtGzjfJXZrbIh65aZvziF96NvczIAOJw5Avln/wEwmnkVZsPVlc
oGAReSdOtlt5NL7zLvacqRGrrmGY+UYTUXYKJeTHy2VgHSid6c0QxdOSNfGmH3xK
Ced9Jr+BOuuzMX5OcMat6LYg+L77UUZYE/9HH09ldgjOn8zxVAKR7OyUCkZkWwVt
04qITXc7nOp0iv2WGPfobOuxjQUX0MI2aO7f+sVqJimxXoeW3H5DZBe/QclOGgz/
/IR3jeu4MJb6xaBEoih6Zou9zhs0OeHMR93HIhl2R6Aozhev7T/EjGubHaZEObjM
aBTN1IduXvMFftHJEL+byqCJx1c6GNoUcrrHlpZi23Qa/I22F0RIFBOCIBwnoc/Y
HEEz4AnPmO2Qa60RTd0FjZyHzGnSNam16mUpAe+MA/F/lcL2To85ZPK3tfMV2lpg
wT94yb+xzpcPD0TYbHDtWW8LYrapgiuGCYP7sNLbW+etWsOSUUH2RlGGTb0jw/13
Y7MCYJSxozTLktw/i0PzCtLVxbhoAE7huFKnnho1MhLqv5wStC+AD6Lhb9C8AFGO
j3bBc7kwtwMk1qywT2wnxC0SRuBS2P0du2DaRgz7gQbNY6vzR7sXN+pF1cWNINiw
LxSEPcvZo9VusTa3cLdr+z0d675xHy+hWEZ835xiHAFNoXlDla1jGBbNqmo7ZHWE
6GgNHC1oRZLZ+0d4+3ksOENWFNlNlLkZz5zKmm97jxtxJ3RPXZXSh+wkmAlVSR5D
nRfGsozjk8Y+3KCBPPaZ1vP53Ci/Nzp6RDt5u5lpiIXGdRyHN2WqRnDR3L/roe6r
kVgk0mTXpT+oaK25XAG7bhwOyjYzJuryHSAxPZwXhKfbGjexm1r7GOGj2G7kFMh+
eacSAF4HwV7s/26VwIueaNskY62xkTbRkLjTMiNK5wEZzGjvzdW+leTaq22DtSbf
WEWXlF/V4ndUYBcVVRSKLjktcnwzQ8TEUR+iZoJR+Gmte4F6WT/pwFrtPXunj7il
COckyDciCrud70cZLDIsULIXihD1rzAAIgf3R3cl00Zev/iMNpQGu3Y6Bm7PJmwt
eDoxoI97W6uRFX93APjm19/RAhfzN2rmXT6bfqcwwNS81hNp1AdkmoGLTpwFO5CC
LZzrLjDV80fo0Rz1AqfiRiHmVe9Rkb2MBSCx4mhSDVRUk7Xh9ZbgLJTO4bOIF6pE
MHG2tTNAtzMVcG24RBfquwTqaYCX27fvbt04mcuHMWFTyxXb/HLIZyQsgMyhuaJs
8cIlWzKRoZsU0dvtJIDIT+mVdLqJfisfYbqGXptgIAWZH08k+scyyMJ/aTstf5rD
rWxIr0cccP4fpKzqDveyeox84Quwp/Ut0I4ktqZmIZSuGiiLCWI8sSSM61kvWxnv
sIe1E4cy4A6ISX2qssjt9EJWtHC8HdiZAXX1XisQUlemKmtIi64wb6ZkgpbRhDsk
Z2s1h76ZODtOWDa/R/PhqZ4OePTC3LCTxsS168/+rPDOeRh/i220rAd1b7iSal1W
OBNIJEqmDXxJzkW9X5BS0+Ex27x8/qBbv4hqIxd35FkenL2huB5liasneZPyySnD
+gviNog9xxhxz6fTFtdHCJ9IQoi1Z20LKPJVT/LapRnAeePlGkrk6IsLUvax45cS
UmxCBZxtxzFEuGLKwj27jXgH26FWkY5Hb1X+SQ0bG1BFsLS2D3cVXohKBryUEB6+
VgDMirHXplZfwL7g5IPLvFDCtL2IgIdRNEOUaG/Qps03obpy8efUYBsGjE9SdShJ
1V5o6C+pcQoLFXjgLhBzeaIy3ziKiuEs65Vv4NAKk9TDPURPvY6azjsC0Q0BRMgb
fYNtNMKLiJhZvXRDUnNFUR8thWKxZH6LEigBaJgAuSKQC+LQVLNLOs2MBovaAYZx
QdRe5+/G3VF7YANyxLTv8FRErPvS7eVS3gRri+BkIfMROPHeXpcao/cGoK2aMXm1
WVcRykwaRKo2fl6IKaQxRr1XHf4Z7JPmVYw0ZcOJ13/5oQp0zQhhG0uTdaVUOvfr
Uezh3RLLFLdCvNjBHpG30uquVBReaRxiL11fwBw5J5Ogtwexrf2NoiZByDQvS6Iw
lcTYlRu31hOqB+O+ZX3Wf7mLYR0yeEhm3ycdvNgo2kaIz8SqUjohl/p+iaTwvA6t
Lts6DYoQc4KkPYNYBd7C2D0UZm3krLCq4q/V8DUyYf//2yCUiCmICo16poy3E8JI
nzp6aSiJu5z2g5T6XpwkWoOErzqk6ZOpZz0FEuNnOk6zAqm3ArGCzL4VfaGxjmBo
5mYDxsbB2VUAnpxIHnp92CLQmVdTmVo538gDg34TJcy9ja/2zAAuKhBtKUpmNht5
adMgXgH4JQ0+8X3upxNZyu4tl7z1jd6OC4+Xqd2NTHq0vvbLKyJ24791pKqNXFsY
zwxuCHoK2s6L5B23utIY4liuJc9eX78GOFvhfSOdUifyyrap09cwNVrXxhukStBO
+l0R5edf70w9Vx+mr+lTST9KnMCtqY4Q4/MUNSqcGkfDBAbqpReXcsYVZQOUu8+e
ZN9G9xeNohrnBk7RGXd82En8Jt4iKgXvYP5oG6ZtaKgzN8PoDoQIuvPoBzbACYjj
IFetBVEerdvhUOZ0x2ZwLTiOTRTso0NRoz7ZrEak6G9aNfSSyOZvzqqGPypCBIe/
To19m3OS8D+8Qdsi1grNCo4bpdk8FllgVTrIDFKqrB31EyliqvcLxizRipJLcvZ8
SucMQR995OSbYvkgTTCsnhb63/OBnIYWI4Nk9vXUmhyJzA04KQ0inuufueloH0sp
sb0ht7d7qd6eCwyt0XwbUI/9bBpcbllCbKRWssU04U9JAWNZsYz4FeOuCMid3ZTC
L/4VFVTVcv7PWGsxlqjIlb6u0bzTzv+jvGj4Z+f36eUGwuu+eXlEtAdisSxuLES/
ReS/oPlQkVv8Rh+bB2J7X3nyWK3wYh/K7G0I3lRz3tbdvyq+TbiTICYUxXDAzHSC
kowiCi7eDuX+U/AGZ0vV/OLFtXzXj7vRnvwFb7NgLUfgOhVTUI4ucJ8mWBbUXhzT
P79gZN2UsZjBdu2tmOnXMMo2dPttOy+I0j5EAUtx7drZqAm5Y4GL65kYdjg6Lhs1
0eoH8iuRtdJKdnvFVyFXvU6x5sWgw6Dlyd/gEXlRuT89lhnVYt/a9/p9eabVT/As
sK9Yd778b7rQTqZbA6ktlIEKvoCHVtnm/ojf0xwuoQNCogM0/s+UPmY7432gzWE/
yZPuubaBlMAaKKbpD8m6pzOW1WwasBX9T+HxXSbzK0Zx+SxZxYE2Vb5QDhPJri5i
3CmjylMPOnMSr8FekaebYcMY7xfbSnrzGlKPZc+CazsEkpirWZ9otbVrvH6uKJvd
E69Go+cNAtGxBoPyPGGJKqG60tH5nwcgnRsPXcWhHIW09FNCJL0xOR4jF06ri0AX
oopWB7/HjrDbQwkFVBa5X6uDtlXJIvJ06En2WjDXpUayTo8YCu1jBrK7hqMaVJEK
kLpu7mdW9aX4AzYvf9AsUyGe+I+02fXoF8i3+Xo+t/67YFIEjiclmK5NysJDln18
6excGSsX8u4bZspKPkNruNoQ+u1pus4HunnBkuX+runcphTsoYR7RpkmHyp1tv11
AJTm5xui7h4Ad3untameGDHlUh+9u/MO3QYRu1GsuEc/zqUZjg9Um7q9ekGFUS//
OPBgAEYeMXdBnm+LD7WPUQxRn40Zo3HxBjbR1t98C2bPHQPs0oR/b2nhc9KA3xnB
p+Ti0vPiE8hya94hD5R10nAqqaVkEVi5m6FqMZ2pKfvR5A8U9bWyaLfTJYQBiyn+
9BRXGxQ9H6TcLa4wZsA/phEZwudKGZfA113EdI+YpxC7/KFfXP1oRSl1fRtf/xuF
YolOviA79eEXFp9LsW70oD0y5RNYQ62HKQ50aDKQxbCpM5PdsTMKKdWQBocSziMo
opGH65G5hkeY5OKPAOavjChxUCrIycLrsnbb5RjygVIZ/1ArsZ3uWFjknCoE4GSH
jznI2AzAQ92fTJP/tiLashsMMq3mZv79XKhPNeLwEhXEmK9Cn+kyYeHFxhUR/QUb
tEXKHGjBKI//ONTHU3X/BEzFmw64wJIf4N5PXRz/qykVZ6yKpAcDFE5oc45GHpM9
IvM3LMeFChUvO3mu1L6rgENmXHTDeDNzpe/8iBDWLUlfMkpTKkEGUgqC/YDh+WXP
jDUPIXfnLSwqAikQ2PtXdQKBcBTNjcXSXdZ1pt343HR2zhBW9Tt9a11/kH5LvWW2
Co6sSsGdR3CHrKaI+Q9mv4ogVx6O9RreMHkVmaNrPr0WklY4B6vJrw3H2sNN0Yxz
gDkyxFpVJRhT4XD26RxcUv4UKnBVaYWywlrnGOeQrmnj+rloIqdr+V1t+XuuGODu
M9O0nBxa0pyl/QG8//QJO02N4noNmk1q8RfhfsP0H8xPxkH12tpRES6mSIGh0rsM
l8lTSR6R0EvD37PB3E5bytQtV+YVC6Q8zfBNHFPERubbQDJMqNy+a888YE3v5RdZ
5gApW2PnZQant25BOSIbzpxqCm6//mecU/MKHz+bAw5clyCEYlWx5hJYttxj4CIo
SA4j80+Ds+Jg7OESo5NzUFEDPq5iGW6VW73hKPCD57KWA67r6h27yqUOS2EFiD1v
48wV9YBPEc5xdpfMTfJPGDp3JIQjklkZc20a1eFrom8M0pxMG/QrZt7x5C5Brire
Oq0sr0gOJ8S9wFy3V6a+K/TSvekJcbLFnevKwo0YsR87NpneftUcNnzLsi6AKany
NkG0YaEYfeeqh5mTrt07Mpc5qwSncGJxLdsnM5jRD/kB8pvuo0lGEr2S7KYT+yzS
Xq1oseDASj3aqpwdcgw3w9xXnblHpvmlxZlNew16n/9Y17Zl3RK1ZbqMxM1mmmBr
YvLCs/ILZYQv/QIVfIv09WT8/b5k3dMBIf5qUwngIrJDq872lN0u1akkv3lk9m/a
Gik4YWQuobumu+KwgfzXUZ12KcKgaRqgg54QJl/X5TkP5TgGdLIH1bTG37F6BFI7
0pILicWeZRv52ZPeCYgU1uQxiL+NxHTIbh88p50StOV/2/cuXiI45QY3kh+vuXaw
iTCYJ0dcROTuxIYLvZxnbJrVqCE+LRczkT5r76H5TBqcweDOkLXtsdGWmcKRoq76
nKfoeX+Kr/8zIoB3HMBJOb4jnWDWqYT6prEkcD4DQqkko0T/+zorm96UZ89OSS+s
FdunKCBHvKk99E80Rw/pAP7Bz0H5gXeveEu2Yfll21hLr4O3qNunROultg4E2fgV
R/YidS3edkIzl7L1Vkvk4sS0CMTBGXdiTW30H0L54N51ax60uw8TWQsbBYxg2xcV
3JLuiD/ZnNXYLyPsWmNzPFjvn0aMUdiFSd8n6PPveFPQ0YbKvg20GvMqlUnJFmOL
YyH1Nrf0LgJfVeu+hwbmzZUdA+rnrWNe7n8o/OuHwSD/OG8/kzeNenqCM/zBlAaD
jmMJeaiqQkw8a02ImIri5nvpRl7iMFfgwPI1ZQuwxtaEP46hef2vducilZhXXGVz
5rqL9E74OQDABcTCmYUlM4LSh7CcFMJHGlIeVQdzxq+Oz3qGVSpBROLah1jjGtO9
Oq5JZBgj2XsiFnUYsoATfJf45vQjBbcnD9ktzxnEW1yLDm3r06AUAosiWu/bAK4R
2KorU7x6DHKwgZFzS/Zd7FnRhZSdNn7z+7aEYFdkrgsynFRL6uytFn38hyV2xRwV
fzqrE+YT0LMz5DoRWQzDk6jln/JUnGQOv92+/s6BEvWVh/JEO6GhH6+nxY+Aa1ZT
UmSV0i94QLFITkMf6SqQG9JT3vBXaYOHn+qFJpmsHe30A2rcsLAAFn/5ZWZaW52w
Kz7cXKXWJnauYqf1Q2Ax/GjU7rBxkdx3oINWSF9gaWGVaK+IpZvhS0M1psQ2SbuN
83FkcnPPNnNB6UjzHZb1Dv4v6lsl7ZBCQN2Te5juAKhLTD5tU1pmv/hc30gA71AN
94FncEWgcVcbCHc4mrtgSmimr0RSOwPFkTlH12wIkaocY5F/XuukK8FElsKI6Q3t
vFSzwLqyBl/Q4mVfbEQGhZwY5umV9YbcO1D3/8EVHviZco3Pjh5tOlvRfBtpvIul
Cd71DaSrngBaoLUfGFuVWrfdeIPzrjkAZ1Y550EQBSjZ3ekzJHcEGkS2X4wyU6MW
O3j8yjdUVDjnu9TA2dMJ+z9L2z3Wvlnq/mGODCv5TAX7ou6FLwwJppTGaEZeWR93
1/iiTd+FWWkLjOsF62xQVfamYQXOXYyCr+InTSSEe3ezjLQ9QJJK6FNq/mZ+IAcX
9LNbmRA/biyEv1NlXQXlpTO355WCSyYwE43dTgjY14WhihUkrsPDgpMwAtTEiwv/
OnAftYrTETdLa4RIVwobGGAHXgZ7QZwVmIAXnxr/JlB/L2QCw0Lig31pYNqe4MxI
IT2SnjWVyw/bjUSpMQV3MytcQUvJTg9yEwHoN+Hh4XEaZC4fboVsuWht4j6HLAzq
bent1nqAmBe8ZhCbHpLGvDkSmd8AW28gP7pmDoL7wLo4v1miolMlfrfg5cohLxrq
PcGWFgJlmsRsju6MZi6uLqZTHa8zA197NxUowj2+SqxzV0HSoeJlcAp0tCfOQW4H
Zs1is5mFXjqgaNJhkYFCV6QyV/CNjfk4uxu1RU6DxLXgX8zi6T9y2SCpsYPVG8eS
i3qrcZX6M03VjdKXpfhqxv6PGCV81GdzsRsRICQifQVNwavDnwp7TVQT8DRWV24g
/0HYJnI/eVw9tnPUdHQPT11BxekyxlKHblb8AOTNHfQgH690xEV3FCYijIh86YK4
6XddFoMhwCGxBUu66FTaZEhq4gohOhsmtAiw6iVeV6Ih+PddnQG6thcHHDL+sFZm
HEeFs0zxFH5iumEHu5QmDuNdcTra/Wz3We0XS7fMnfCqLJk019uHruZRaTdOc2AH
H4qNubjwAGAljMmZq5YFattD4D1lhRix9PmO77h0m6I+KFpkwpFEwXFowy4TofeP
eFy8wHseQFBfcaL3opVMCn1e/BBXQM5hIHS0qRUdMIZd3q/KEn5ZWc/Z3afZsCWG
g5gQUtU9ZkjKl2dWL2oY5NeCIf+hTf2r0PTkPNYS7Xp5e8UhOUBAgPkJpbYHNskp
br1nQvip3eUBt3IHkdsS/f4AuTixjwXa5ci9koQSvrt1zlB2v13dxor8x6n1KCYG
F22jgSW75v5GAcF6YYWFbWYqMNvY8R370m101AAri3OBkvCNNjfIPgLlLcKcnM+E
958wuN/knaTyAm6mao8XZ1dbEnIMJJOpEQR6b91aF1EoRdKdVD59NiJiIn0SAWDb
ED3k/d8sAoKN3omr6Wau3rDkbLzqvA3wkzh0hXr4R5G3EEAT1AsGb2kYXupYkdLG
96mHFHN62IE62ESrSoXVFzhdqwnRRxZmxElSelR/338zqnAzFyOPUsxAi3dz0mIh
dD9X/cwGM5OPKTubBzykoyh8qkMVilj+WNa8x3GPrqkkm0RTTGM/Nyg00mhMwoSi
TCagFUb66qw0RNTf1gn523+OU1gGNckQHItxZqmWRxhJaYr813kNO6Deb5fn4Yd/
eh/0lneGkHdEH5xYyCBfr1cVSK72UEkXMhQw5mLkBZkX3O1ZsgoqfkckE8prXuEg
64VISE4NpUSseLok5WzHpOgTD7K63/0gipCB/hWzMweyGdQhhNqoKPSBIluW5Km1
4rBuRPb5Nw1TGECchZtmmP/0Bx8pk3YrH4l1AwsUM6vQ/3AHDdQcdInzlj9bbtTQ
k0tdQpuNDYqM3VV1Q9jxRQ9ZdEp+OEq1ZKCWQz2GALJ5q6N99GsVkAX13D0c35bU
7E8Kl2bjpKx8BpdyE+ZFThiINYERmbv6a8Y2EMt1GXjxKl6OH6f7V60SOxjzA8fP
Ju4aeA6sf6PHc2kZQWeDU26iIGn/YzOBBRnrzsUwEBwElSh55qSq3031zL48/BqF
/XWK8I/aEC0sXSfdBfJau7LULObWPtqVhgszG9Y6za8aZoy+e8IvaxSunZwAjIiL
VonxcQgWFfyfx61n8zfzy4Lo3RBOIy0AuUy571V4HXqHUolInsh37w3Lyr44US3Y
AMHiujnCosShwW3eHk1xozDea86CVtFvtir/5lZXG5wOAmPIBAXb1pbsO/XO6cIk
f6SY+q3ryyFu36J/g/eHkZcYq5k6mf3BWtNO5RSlQ3x2LUmcGO/MIDM2DK6ZE9mB
e2TMDHd+zulqMzDP/VRRYNe2Zr8isZar13tmXg8Tgb/cmApSK+DTjQZp31oV8O86
lkDpaCHFKI/5+pksED6P9TfjRq6VMOs1oJ80+I05JpIu4FCayFfzCo9Sa0MlMGuZ
fXjrqf4WnKBnVfuuqgzi0AOjog0B2TfwyO85dHQLJ19gXoKF5PXEbRMBdwoiFt4k
VzNYNM9otnpZlv6MU1Abr0duT+By/Xy2CCnhRnmBsbpRf5fo6hiK0Acq5i6YsAQz
VOvR7U/dkCKBsXTsWa92JgOB+S//zk7mXWrg+AWPNidNeK9qQiIfhBJ+xc8aRV7l
yjpdpX0oltV9jNfn5uYBmfRGVrvqxrdFTr8Li6DihVRvzcuqF1ikKqIPACEqENcR
oDpo6QOCiK0JoGkOAcKI8dFkDyCff93vy0tgWO4GRcJV/iUP6SeFypeQv54N6IVV
UPE9ceKdTCgz0frdVaK/rsgcWhD8qWWb0z2mLRt+yxhIBg/SQ2XEIJyVL/ZK6J8l
MUpTG8i0GXa1/VacrWrXXbTOsf6bHTNPcQM4xcQ4m5b+Jk+4arBt5jytAvkQJVu2
qh4HcSAQgit03t631XHUjOVARTEMTxtAAn9rWvuuwjCRaJrCq52YDrd9WV/9bONC
SOOOwgfxgrtGnfdod7Rv5+wTcSDurfzfyEm0GK20yyWZ3FWAnEO4mW0vqkLYg5Zl
Ghwd5p/wyIqCSpKrRxwg7iCKnQJHyURctLjIdpnayWlJNG767XMTUpocxWTZdnfg
knBwjuZNek2Vw6kODgN59ulh7MeYdoMN+QloFiYx74/K0B2f55EyHFsjkdc2ICay
GKHyNvNVqyLMa/J/yKiMc9mmA4hVvliVWrytQLeiA+dgjz/szQmDgTKzWT67Hmkf
2NGiCvGZWAVT9QATS6shgsTJ0Vk2Nbaik6LwKw8FQEtCmKGyM0/XUEjp2Dq3Q1Sy
prqfZXlYq+Q1ZoMStBeAjYPRh9XkVPFvZNk+O4ALh7ZOQQtKhlOtlGTCuCWkwdU1
yS82bigeohw8mpSDqXmLQo2suba2MR1XKrHqk7+6/XoXlKucPhdBxpKIfpiy2u53
qsK1y0VshKusaiXb9xqTh8xWczFFqg6n3nG6KLZcyYzlZ+Z0pLgdRB+cf4H64pZA
jeySR4oIrc6paiGT2YWxSsEI7I2vjBBYK3mgrE725xuL1RSrF8gN99ZKAYcZN5B0
DPJTwvJUtOyaXmC20pKcJ47gJry5aBmPG12+DWHoPhvvtYqEpJUSfilP8Brvd2hX
awHZVRezDm0Z2lSYdOBqBw7puhHhjgf263sdLReUsdvTNKOisXXrEpO9RjNepetg
LkYJokMBCYCLBlDpoNN7YYFkLpZgAYwdiK5K4QVcYYAJpMHuLK9a0XQApldZfeGy
rUKSi4BNl8QmNoz2UZWYiXGzQ0iZzw10xsr74svy8235n3EUc+bcWw48LtH7pWXU
mGEGCcbDZxpJCCyHHqyMm9D4LcariH4SDB9aAebQHxfSdOnJxlPBoWbN90alt5B9
8qwF5YJrq3uDwrFxD5Dl2cSxdOX5fXTq6VJWqa/rwvqcvvr/gEEmHRYLRFpjGS2f
/AjnWeAfETmZxLCtNlyhtExrw6r4OyqkaCq2uMlO3tqPhnQHtCzcLjv8IwH3vu7V
tBU5TBhnxG5ZcassCjCdQB19CcZYcPUlCMZjOdTEQarZlHGqmd9QlYv+JPROSyhf
qxiKi2V5KY/nK5S5Jv9dZiuC0CSJmrIYpEoWTPClYjD4mtm9kb23eL1nGfrUsEMp
XqXK6Y1AiDYVofhs7KqKrR0oMVDKhbwBYcjs1i7vByTtEKy5lV2qQfVdRL92Gprh
emxWweh6YGnpEauJp7JUzNwMmTtMISUa0c/uaqCvN+qTNvPQSz8YONwHG/XtYD0L
OgGXSDMDS+Gj3Q7EVvNUbgzlXyYLLrCINRkkFMCJrRc/1Ud0zmVUuFlrvxyC8BnE
fn4oMJIw0+BnMC3H9AddN7+VNDAsDn0CdbQmeIp9WVnZeyXoLkvFomSiaw+W1lGA
Tidygzc9mpPehbgaSNn5SByNbhmE9ozjwWBq/EcXIh1+18IyLqEsJOSbR5ZgjA+L
bRlnibSGD885pvKXzuQUI+1J1kM8l0RotLtAOGgjAL23iUACPBXTkHZVe4YJyXLJ
W33fUk1ctkYKwMkTR5gy2jW9O1ghKMAejN10FeBV4LOQTrpKUWh7zxVDCjRKNbL0
ixySV/izVmgfj/CcHe6eZQOvjeA4q1zmbADL5Ucdxc622+kr3U2Gnc4ag8NY36N3
9EkJ3hhZdjRr51TzruM5BdFIQF0LLzM56/a5Zgo05RiLy6wJ7XyNmMVdQ4x1txI7
TWYgZvINS099z2MqSQ9FPLLHsCUv8vVqMvFnU16UbB4To4fgTW/VWvFL0by7yzIX
YCYWmUjPO93SOvrpKzUMPdNVDsXTKGfPXKmQLTutGlI6RhhiDI5LJvxg3NfYlPhP
Si2PXoEkLLjnTWOu2Cq3Pq1DdQNSrlUwvyYn0L0b6cEFH5SK2nrJBWvSNgFL9tu6
yBYhMZ0iSqzf9AipTuoBcJ8mysGyzJatq/1LRj6dnmKP8arqwCFGhjJ+0nflE6+L
iTJRttQagqPU7IoMOVFrWRU90Kephu8teyam0mpvD9lPPGNyKorwsmbAGHNpuLxt
kRM6RZOR8RV05zo9iImHtfEojMeZkF5iF3XK7GBljgUdbLEme5wQYMR+emT9lJyi
yIIstR+ljE3vC82ZFfvd1Q8KFw53qgiXGomXLr2hVbqtl7HnzREI6g4W1391rDBj
0MfqmQ3RhGQAaE/p7Cfp8kEMVNyobtgtFaUiD5jPM6FP1AmzC6n9dlTNFDU5jEll
Hpa8BEd7YKgk7azF01TojkZCFa4Azgr32N1sADLE/KNlVmP9kuyw0JMVJzormNgz
3+53cWwW2HY2P+efJLwPpXdVuLJh3imaKQWOHdMMnD7qc0pSNzeLygL5XJcbvceB
BgP3Tt1GBkRCeMs8Jeci0gC26S6oQipx7rt68bTckQQDqfqi1Kt/htgcZQIm05FM
5Reues0dhfRpsXDRO7RqYrVyoTzW23s4tnz5+HWQE4GTCRrC4BcOY02iGMlKD4A7
9IOgeahXycOs0kZCn4pcygVN1ujWWZNOYpN7YTkanzx6qdhX/uceJcxRwwr8AflA
wVM/cbwSrYY1i7lHKoIOfg1mRGmzih0okg8s+WuChKQNExrq9ABoLuxLMUYfsUCL
Yv/QwXR9prKQQWRdDcxb/6IEGlz0KDhko2W8jBVYZhl3PfWUddBpSF5VAMkByPzd
Qzfe32FFoEmz/uv3S3QER3ezQnSDLlUjSPDbPuh8Qk/9wiT9VyJkf4aAm/Z6fOOi
WdvIVoOhE8nelYVI2SdYG4NLTab7b6m4fv3jL+tLnAa8UktofeGcjq2UAlaTl6yn
/ZiyxglGcL96lUL3+lGnrcASA8+Hj/usp6OLjPVIrDJ6swfe+I16l+UCLePOsjtY
sVKgGAOzOHmr+kfe3TFtY2kfSMxoWh00NQ3f2RQbVNuKzCH5JPFtCF/Zx1+PW1zs
o1xYM7F4G8VZyzsbumcy35be8kNiYMCvdx4CYamZheVbRIaK59ePN6CEHXRrZMQq
aelBpEzT7RR6JgSKpvubqZs8OEZHcv8N3jleDkn3YaEj0L+R0quUGDT9c4O+0+cN
0tI6Z4TUHlEVH+YVSMhwOZhPaPdOCyir8dBXFohqpHB6c2+dWZFjfyJvJv9XVOEz
NfuJdk18yfg0puTIHtwUGSMeDOK7VxIGApnfv1/z/zHV8yEos8lmp6PyB7G1VwbV
NF597ex4uiqc4aKvbgFBP5qbzLAB6NvQxHYk3f6GBgUSsVIiYQhedLZV+D7dl+8I
oVZfMTLNqTsB2NxiLz0GE46HacCkn2rV26AN8WnHJJ+gafm/9dQqCx/CzVGZpjHb
cucUhwACLNoO23OrY1m+FNFoqtaS08HqGlGWI+PMfDWpmAxo1KNVSuJpEp77PdIV
kfvpWLwBBoOJbzxdjIldeNdpK0gTpivECMbtUVzzNGvu/7jEkEti04kKvVhuMvHF
lbQ29HgcBafSRWvz9pP4OdH8DHVterFlem5xcFtY/mhK1RGkZHz56qgPJCvwyEvB
D1mUGgSHAz843a5+PNUhg/Nb78JpgzJLOUG7ltJaazuh1/PFooN8bKkJ6glaR+q2
7v2aEVN4DF++/MOIH2fKojaY3CJ6woE51Fi1seZdMGg2W96TK52B4Srf3W+Wo8ow
ba+W7U7NHnaFGmJMZARu0MLo3lvstT+IHp/OP4ob9UIKYeMC7X2Pu9urHBid8ZGH
A8vumgHw3XvjJFNJA9NFDFCQlwF4F4xdVxisbDl4CyfJZzNSo5V/AbNQT3CUKMox
3HtLwriVreB9YBF1CkXIAW8RZA0QTKVrLoZFvrglGfKwtgRTMmtQ8ChaZJ2YxyIG
56GPvtLq3S3PMLPRoFg4H1dtGbaLZZUF8DCh2f38Ga/RQuC67AVEh/F+nUYHzqwY
kgWSgW4AjZsJVG+VzHzCPfnLl1XiqLHKXZRTDVYegGtx7y2TJ73BDWhivljjdyJK
YNLuXmdd6B+FC28yJZxf4LOuKTptCEqvwoEmEY/HaNuYAcUYAGYWXP04T1YJqNKD
2xlRpcpvOVg9yK8Y+qfll4dpd6aY0GQZLgwWnGtGBQWPFFVnC3YljRxojyAmigsV
xvexYVfrLNo7sOoSK9/XkhpYXGS4VO3IbAlxVwtecP7Hfg//nfPrei33BtNx0xap
VI69ycOE63NWoN3d2tcK5p0RAtnB+vvMTfF04NHcCMmPFRXaqo9iEs1gAcxMj/DT
GmWqY1SPNW3M0B/SbwcBDrIXpIHSNoei2oJrIkK3dwDWwREWOuI8kE1UBO+CGR0G
gsU/Qy3yUXdgNJhhKo6ByCVcNasWruw4bysNs7+1i+ot17I6mguBFOAAJZ4PC+kJ
mw3Rtl2HaEH6TPQAGELzPjiEUO/WQRbU8eqlOLSeavnxBNDErd7M6rpLvs2XNkIQ
4t6woyw8DlaFtMzBCPQjT3tqGjJi0U65uKT7UlhUaHpeCet67UJhpqNiySdRSIhB
TnnJKK9No/Bbn8CK/mz/itMZVKGq/tjOXgotCNm684mAbIzf0q/SO+zxM/AL0uFe
MMBPIPafDejmF4DKqaMDVNgPAYyhjDohs0x1kbQNjAj6YUwfLy575JuEOiuRe0pQ
sExkN/T9zO/HxQgXb3yFG8ctRLWbK24ompS3A+gnTYN1JmUwbdWO2MVxtXd/edN5
HScoVYJTDRW1hJTe7HJ/hErVjAYHdUDvKCqNl+2Hn/Ux1HsE0Zhiqh0bKrs/7uyS
l/4atEInoiFcTyDDwC6gHNfD2PX9W2zX+HHqAmqAEr0CPdkSohJuApPULKwFhPNk
0wvN/p9qJ/mERLFkLVz5eetX0oayNFmSaqLkJfDl1Wu3WAte80sN0GNaEteK4czj
sQrNwm0RdvmsIO58LHr3funQdgW8zC2bMVMA0sWDUillFUC5R4Rkpsk8e3qBEx/f
QWkYCDFEdWxR1J4nIJyd6EUU9JgWzdF+EzPShTvN3QkOL6XtW7z9DNSho41p3J0W
Q5uHRb3Dvtr2hHI8OAvKzOG6hxqkXJWZB6HygZOD0/jzYUGXeQFBnCWCHqxPZk74
w9LubT+JUhKYfHaTZh2rCg4R6BNzt2zkaySTuyxLiqyrDrX2F3AO6FEUYpl/R3Lp
X051InEpGJy/r5Ou+OF/Zs1M8sw0lDXygWLrXNC9dnIa7QZx27yg8DiY27OE6fas
mWBRoX53AS5lNE1NHTxBVzxQpuC8lmuUytCZNntZ/7lxkfU+oD64pVKYo4Pr4kIE
9XXCLofPgncl7tJXIpnFmlG+q8OTj694VRkaO67ZZovuvnTlyUzATM84GRBeZQzA
TOJqtVizkPtE9E4uSfYqT5wYXmgfhxJkVuBm6KN1AIYIBU3qLb9jGqEDRoDe41Ei
2CWWC1gplrrt5WO/bk1tqhd9KArUw3ykL0TO4CZZdkk/KTnL8EdzWQ98Tfi/gM9e
pWli5CafTF2OIHIRTLTrSMXCWF4gmoe3xahHxs35WmqYzqXybYvtEwpGPSa7Aqsv
GMcvRvM2JiJe+3kMXZIMDc/h+4627P07Ej3oABC7dIsodLc7029SLChlNamg9G74
uKSzeoxMQGQimcAsZGgZb+RQNO1HhMxx+MBbiGWgK+i90h5R5Y1AfcYMwjn5xYQp
ShEX3v2PMaTWLsIaIkGTWmqHBAp0klQGBR06L/uQrHiBZoTfOabB/ABXXf4Wo8N8
OqnTwfboco1QraEP9OVXL/rEEXdvnpkRLTZljs9F/5Q6+Xkbe0aVT9KvWM55tuLy
9UBoCilGhtTeMz1qc/Kn3tIBVKm1imOHxVKYo6eOJSFjkXPFIFQQfeGLDmPGuSuD
j0uWtqhyAEC4KCq2HVlrCELGvvz2UzhAkCEEi+gsf8I/pdkRb4pZ6zb3gl25xROv
V1EepXDQeNESwHHmUwk04or28cn/AW4PnuVSjF3FGfo+iE1guwsXdpq0LPWS2yCg
mgUfWAajATPcqFumoSzVnMgOOhtPwKxudfk6UYRZgj15Nhg36tsvWJYOF7xq2Ejp
rlLZIK5zEzU9meU8HYGQsoyJEsWrrUE9D8KLDPEcDLZHqhvBvThcraQpelsyDek0
6dT918tI+WA2JV5T3VeWW+Wfs4Q8SwgcrQgFb7xvOrGrcilKoF83iXKcrWdQmbS6
VCSTfqi9nKAMG/6IXalVYgPtKuke4RvkMes8XJl5WCCoOHIT6JOlokxJLK2oYi7K
Gpb0EfnTumyjQ8SJC9gYh43WEmr3ZfRu3uNQuKx2MvQhYQ/ii9sC5QWbp4ya5AB+
IH+gnbHariTV6c4htlGhACLamTGQmW8j92/1xq2kP+Qwz3gXq4jZ02v7s/yRLExz
k0BzAkb6CvPxdBPSMysm54my3sZpmI6zvjj2XfzsIeVtBfK2aXDzWF9C4Vbd6t/T
QzU+fpMjVGFIu61es+UDi9fm9l93NxXQkDSz6kK7FOdmmp9ZVtwFoDsGLZwvwcqv
PX3cxEcTziDHHvACiY4rPNAFo6tzB1/EOnIsOOZgFndbvpavdR9l4SFQIpZ2XL83
66G++w3lTakvpPdoa7t+1agAhVhMASAEE90HA7CgruKHCHBk1Jne0znRJPjYs3xt
WPGncRrxXalFSTB37Zx4IQrR0kANcPUwkIkUrQp5T/aF5YlDfq6Tdq6+gf3P7VHe
6KieIAYryTWNEK0UZw3HawHC3ZxGN5/j56McSk+eALyjVtKjTrnpsGh8idomZSjb
XeFJnKz1CpOb2r1m7SEsFDbKLaJ7XNwqCD/F/3dPZRCyvnAfZNFILblctVNmWE22
yR2Q0857yoMko9O8Qaw1iAwL5aAsLDaQaFTdOyz0PCvpma9GTQyNb1s0m1FRu7Ab
8VhucPUaPXdZVElO4DN6C3M/eKgQJdFNhWDzCK8HSKCtVzS4U5j2kKanVN8Vn+I5
G3uhCXXmILOKDBtwnNW78dqk1FM8hMow5LFOUs0KXGztd5RRASncwrg7Wy0HatOi
4cZK/rrBIEESKDu46o4Z9mMZBV4WnROr8Z9YaXz5+tUtH6Q8lNGOIJ1dVTsSwqAr
C2XriBEZF8K5FbShUWbSCBMmCJ6vzkMJ6aguT5Uxs4UuZJ24G2YsiZZCOGZmnKpK
YGL9So9hmFYa3N9aUB9Sw2o/rzwlTSNerL6jf5mtRU4FQbCqNilRKdzGVAkPy2v/
rLGGE6q+Gp10lzC365BLVhsCe+LtAJI+4xza7+7DE3A1SlegdvH8WrFgLHvHhUJw
HQb51SmBvoHqODH58Wm3W0PKL/9GFc1++d6Ii3Zgy0fvbjPTXjQ5+323VeCqVJSK
Vk9X0sBQc/NoAg6E7C3ByB/YxCOQq0lsJqJTG5nVNEChmNghAvWBcj7cd/YEBGhd
SaCEBD6Uj35WtdPzncLb0Kg1QNKfAc/6Q0Wrk7qLAJWPSqs7GFzGNPkIOjRLJEqV
N+wv0NO5frUK4CdhP4xztxSPV9Jkquhb3T1Qfwsy7bu9UdyOMR05vpdy3W/p9nLb
TgsCl0y4md12aApWclE3vOHFzR5zatYYWBb+TRXybOVwR455AXINGqcBRR+Fi32I
W3vaVMzHihe7AvqSmAMKM5lP2SIp4R+G2eVPo+9N8rnSE6yG/VggZHb8VJjlz5v0
YO5sgdvHgUI1hoSDT7AGtuJHFBTaO+X9LpiAcL863UTr1/0AkXXTQKsU3DlL6Z6k
dnMS33MugM6LggD04KO8wvU5W52kgHDU2CKT4guT+WWHyh1HEAU2awA6tsiWnrsQ
QAW6tDVNs/wIzotqXedoAZEDsXjtfASgbLSf3lVx62LxqZiI1xg2Ya8Y3lnXPKNy
akQAt7y27ZLMY+M3vjaA6jqBFFCkmVwpYMJX/aREF3TXwXXXeUc8BE7F0UBzeiGu
jP7Quge5rYU7P2DcgZeWJ7pfEykRmxJVW4f/SsxqPpH/PLK9u0PlMI5iT6zTjqfV
cfzovGOIaQRC0IlEm9hWw0/L7Hva/Is4U3swCuoYpJWjv3uHsAnMRRGeN3m65wid
MjoVK0K2hUJbbORCE6855UWCx8RYl82NVSWaKZbXFDZ7UBbat8QRk+zVt1IQbtBU
Cbu9Sp4+oC1MLE0dl/GmNppB5su/boBXi0+HXyieIXFy8QKWYaEPu1p8jF5QZYSg
SAGEkNlx+SGRO3d6t77+NeaPCixvcn9my6Z3rZKHRCDoG33orGwI3UYc1bRQq2uY
XhlzEG5EOvn+O7n5Qoi3w5unCyH+RyptmR0CBl3PA72NOMTYMfuMNRqgUovistB+
Oz50fwEyO42jOgc08b+Gh/CyA1cJbFyuPkjd8IUjUu3dFrtPwaFq+OVOJwIzMYHA
pgnfiZAKE8eSfDOoDFN1vIcc2c+lZEinZx7QVIk2vlx5WD/P01+2+zb1H9M0Cyei
41MuMrIt79xKtE4HUn5T/1ELcZuvUBITrxL1aw2fH+6i9il6TZZboaibgHwYDKKT
fa8F5aw5oCNrpBP6fRFSgyYuLFPCZpuDI9j+f/yUajnNROAAQ2Kl0396nhcWYzSS
YMkZBaWOR5tHufO2kj5mlqG0aARVZ0PPqL2mu0mAOwHmWrBs2vyNvOrMG4fYmKHh
iUSyTqfgndTtBvnwtFD7c0YWS9JItTc/dxBvVxq0RPd1LcwPxdkNAKy41Jq0VI93
3Rpj3scAyBf52YaN0vBZsw94kulLLXsF+dvADFgxsnt/hHqMOV5cA3h5Aosft4Ug
Zf7tc/JiKKoLpFtXQw4brz5b/um7NXIqVykgKG+UIsAS11GeeYBva4A4q5Roq/TY
AXbJAbi2KIoO5gtf780JKYbw/EPE5SFCxA34/q+Ir4vU/dX2ltdLKcdg/qS7zDRZ
f86JxmNiJKMZUTW3gZGli1uKgZ0iC/XZ1/OJxWEM24VFIWM+6V0bUPfBLnzwAA6a
AZqVSU2tAAgyysN6ZUjteQ72wKIuJIWigVt5V2R15/JvKMoF3jNCtV2H0F6ivULz
dspWOKbQYmP30tsXNSW6pgZZHYG1zLq5LPrTSDhYADla2OSPqGYnMiTDFzB4ImEC
ZRDRSnr7YykC+a/Ggpz0Wzvj2aM+X6kV/iSYoPEyrbBWGdgzarEHBzBwpCCQFiKe
YABYdVFXvH4ItDoDSvqDTthMxv9w/Ovk3oyfpvQSbzftrxvMBY5z3VJxpYdRiMMa
CzDniCgz5mJ/X4Tu0IJQOqpY9TLeUIZgv4fD21IwdGnXlszaDek9SI9+nyR0V3Fr
Y/pRM8G9SV+g6LP4DjJnzucBjj2qn4ZomyicVvPQys00vcgqEsmHfgRp71PSl7hU
Us78W6JuJBcATyQQQU1Mz3OBM5qQeuDnckmYg772PGe6u/aJLSAIOkh9z0tITSsI
JCFR58v5GJumterX4ec38/wEf5N1o+zjhilBun8pOJtJUViCPwbWPmD1k418vWhJ
t4Amh+pjpQczK47sMKezJXMCDPOz5zx2i/8jnOFLLrUEF6wLZQ/eDDBE+FOeZ7Lx
2O44/xpDyKZtBHNQvJa3DiS1Pr6YcGD/iq+pncy5mhXKeIrVqM7jI7MGHKWZaO0C
62E7oclTxXmDiuG52cEy003QYRozxjCmUgkfqh4qzH7FkxDTvF70Y0PtO5tcdlGC
aLIiy6unXos8aTMTRca3Xkjq1xZvfmjXBrc4AN5mDBDkSbQknRNKG2xCh7JS1Nyf
f81tswQfqDz/hJn3zpKxj/q5QnGejF/0BxqADHqW1adFpA+fgJww+Atp7Oer4aCm
24vUNgy51QJu6A7U2ngO+deZwmqt2xmnf1j4negygdGx/C6ItPFbfIiLGOfuXGG5
Hp0Lf6hewyL21awPU/Wzk/8tLs3dY0bENxQNbQHjYxMZ2Jr6EUwOgbzMluTP3x2f
tXkJIEJB+VHrDLOavefgXRY2F/xcbkKDlN5bN2LaV0iCelM5KonikPPck9mqH/O0
m5NHJO9AVEDGw2AKJROxQoLnWv5wDSxNY9Y8AHBr8VGr6ENYtOGdiMmGMA4rIybf
4a7u3ZBDgAj6QGlv9L5A9b1NmAE+q+oe32s/cDuOgkzLIE+ve+jRk+44WszvPuk6
LJD0GB1S5Xjfoyig3t0+U7VE80jpz2n3duXpExebYjtDYOPGrJN7eeqT31qrs5yu
+Ij5/Gh781j8fgQiHKaeZ91JlxN6BEZq6xtHJZ/ZzYtnh1/Qtz9qMwGR1LziZUyh
1WVz3qK4Yz7Gk4Y7v1Sau4XSWhk+HbeWFWK1qTh2TnP13yLbzvsypulmV5IyRqnT
OU07fBnAJiDoXcMw1u/K5glbaAqRW6u5kJbJDLCvuTMIU3bKYzU7EQOttZFDGNl7
sqfjKYIqKJMyHBZcxhhvBd5jeFAHKNiQPeCTzhAEGx908RKYUha10Rvr/WoeXSYs
TUhqGqMcOZDRkazsowdkj1V8LwO6qtL/kspbAQf9COFOj/iU7ll7E6La/yVItfkS
xeyNDn4mw05vHyyCBLkITUPr5Ctkrltuv1jzQ7f+oa61Gi8k/Egv06Os4385NEfT
efku8eJ0kn9NO4uzzlYFB84iSMuXWsUTs2yoC7JW3mS9IhxlCWPvxyrFcKhfD2Sk
dmjoZB0324KT5g1Dsh8NMj69+2uJtRE8caLVGz7ur75XEl09i0JN6pvrboMhbwtL
iZzwHWjFfxkSjGou3SaQyU3A3uGAzjZ6PYoSm6J9I2ADSTz4NVo5f3a+dXgFis1J
YW6U8cqWowgPyynoIhmh9XlHUitpf9ONiwJAo1pu40zSD5TMhk58l6LfUoE7Rr+3
t92azY4/Lkc7AWuto/m8V0KOHdgW2d7AmYCf1IU5xmuPMGkchSSCEgQEkDOb7Dag
YMvTfykQnrOq+iZu23oY2ihBAz76vuDcdFgEx7twQpIvBIlAWcFsweJ6pgL0702f
0+2gz9O5VbwUJ5wOyjFNJEWPwjJtJBvZuX5o8vhMgeXRUATyx5qtSDLbELHyitZ1
9GTzndSnSDCtq4WFkxGeL79R6K0vEzGMdV8djgLsSSbxEw0Dd1kb2z/mrDvA+NGe
L45M+Jf/tD3LJsAaqQvi9YtHbpEluV0XOt4aVbq1GhCcVRt/1h9t0qZvLRHMsXe+
jQaIYlYesvvQuTlJrN4MF/1ngTK9QIPyhrfrkZGl8FQDl/bEsPPOL/BccGaTu7lj
CMVKwa4CjdTnxARa6YGbM1x7MAIrfAh22N/Y52qsH4IiiwWpc+5y7ueDy8ImDbsS
BSUA79RmLq+aMETShAyp1HJUU78aE2aNfmkiasGndHG4OvdXSzdYtT3d8ytxOQXy
tZHIsKIDEq5gjPpDK1sE/UmbIuG6jqNE6ySjODYRZOADHkMz/UmuszrY5Wt9nOQn
RmdXy2pe2EECMGDAQXPHmqeGr2qIOftGeEyffLYp9f+RbXnvIBg/nzlyputeO1Iz
eAYaZtEYOE8HpSWmVwTPtjocD/KqUz3kx/QSGu0wC9jDuNFs1sC32n5aIyarbqTb
RocNff2ocUVFe+0uF8Nqja6lYDxqF1TOSliSeeEFkG+JoumfdHgBnby7GOKfphKm
cAKRNcsJUC0PSGn80fi0oBfI2KGWltw2y1r2IgLfcOfcj02keTEgXIxL8HkjM044
7Cn03le12A3/hFb7kTf3aShpmwoFR7ZXjJonmEBE04FD08McfIxTkO/UagN23GxF
obv3NOoUzlKeMWJog+a/2CeEtN5+edjxF8lbOpbdqM1B+jC3H8DIeIZ3Q0V2IFFW
Qf/CRL5RoJ8ZvUxV6MgjLyzYGgls3lIuGD20gexfkdQfP/XMf06rZuStvDwIcbM0
N/VtlrI8/1TUfb7XafLJCC08NHxiwC6wTo0j+nvvNRBpI6xRYW8tB4mkgVwvN8or
f80xtZ06I7SHjFQuYElpXUWAxtLWM4TX1l/B2TM/rPuZLwXqWjfMkcvUEJk6ofdI
7QVyC2UQMwDVju6e1OJm35bKdsWJU+EvhOcqG+9JqHkSyYXYhwoGuMZkTmjCCT2e
ZMRTPVnfHHFERHe7KBTMqhwGlqhFRcq5d9uoqutB/kw7GPNguD+9jzHSXYkteNvo
3vViFQ/u6EHdC1G2pM++BQgBDSjgmwS8+WjLHasuhiRH9b0+qY+/fuVAT8r+Kjmw
B02QgnKPUQzY3O4KQSXIVCcxsCwwGsxOzmtqosJXKeNxdFEXpDkkLdkFNCBTxN0e
a7FchWZOPoB7wPKZNQGzF1Br8REnaeHs5HRbvOXkRyDnGWnGqQsnvumlBZgH5DnG
Kn5LBAzKSISyBeOoKXld/TA3QnU3/7FSKR2dI/Ick1T3zk0fCUvwmLPMUwxeB4Sk
/rKGE2M9Aw2wRccw095WCjSCVxySdLqsJQBzbZ+GzX1C+j3zDlbXbGeVP5ceF9Hd
7N9SoSbqg/T4gR2I59i6uWLCBkPduFVptqrZ5YbD4LUZEsNty3+SWN2so2RwwUyH
l/05peKtDLapOKBSd1vzNi1NctGQnCBJbhQ48ndwwCPiqSiWVnLPQNIRbxkfUkAh
vQQtk0mVIV50YtEMGwAl+xOP4Y83tqGPpfrodtEh9Yme0hi+9bEmo6MI3fWYWH4O
0MtZdMafBF3nAotdrNK/C39lSEyhsAU7t2Z7+pmttPoVgsvHqppHKgbG//woomHT
Wjk18vRO5/IK6+6YZB4X1EHWVo3INzIFTntQXDL8zm29OraezHsZHBvPcAsezwz9
91Su5ZCLt/A8FwlwvMuSi+tEcNDi2bCl4VqK4nMBYPGcNSt/VgCijOq2RLBfSjTZ
zrV/43l82TbnZ+llb/pBbHosrQkdchYNeW4bb90a5Nn1J3yGtvZiLCVf5EF2n6A3
OTd/M3xBPVUnDk4xA2dIzsLJF4C5Sg9GPUmIzEeoSeInz7ZCjNSDt5o7ZlGDRmoT
GY5CuXci0bmn8TYKxUeQ3OkGjOg7xWbnKNTNzUg6gcXvbJvDpkSH3jH1HELNVDBW
H13UjQPPHyElwczZraVSiix4asvM07HFiEQovpfYCLtxm7uck8Ajb6Sca03QhUhH
+RN2r/WCexgm0AOKh4zdh7Fog6XEdwsigKr4R9ksc/s51gwA1mHK9fERO4MmWbVR
vGTvXvvj9w98C30jAVmstIThXDTPZHvafV2AMTbYYzIg0K7UjGz/p8YPWkzOS5BC
HQJpJ2qn5xOPd2AFruh5YqFe6xL2OG0oTB3nmgzaEXmmR+uIRuOuDZUY7AFsMWCS
ttkAYMryzCtTcC1EpdK130MYxTyKtPX0jVTYK6Xp/BEescjnWLNh+rge6YChvrN/
f9Wa3EjL49wzjYKhxrDL8Q4pFBr4UviXvtF7WVZKKKpUCgvGuewdAKLyVpAdpifr
w3OZf6qqcxqO9dDF606I8NPcxcVHvYVDnvHlN/ktINOr19crdjehyunkNgFEpuuL
/G2tTKIIX5HgQuDlVBnZu0Za5KQ/EKy3bhtrzhV6iU0zT64S91zWK2FmfvePOD+n
7trL11aTsx+E0+xMRd7FKCc/RqLTaZ62ZjSJYlbVuq2ahxq3qDoiSf46pjQTkzAn
e2FgrENw/ddeEKofpORrkWRd1KxWUnqBqgwb0KsVp0dEeGlfNUaJmrAxughWU2BN
3+Mxfo2ST12L81hzXzfrpFJViR3Y6dEyWt4NUVAGlvpCdFWnpXz5uI/ILjKNHx5y
n9o9dFExu4Zj4Ig8Q0yX819fsNDkXF65i/L222OPk4X3Rcm7+nuYRrxlbfLC8O5u
OVwuQZCjBppkOMict6XAMNUubB17GN3/CRIMZb8b49wRc/D7OTwi+MWJTza3SGt3
W/4Lbx0enoqekz1IhMtLElz3YPWbMGg7MnvPDk/a2E534Iinyd4SzbA/GcDC1aLP
OqQcJI/P8UIzrMxTLDjNu4Od2xpNb5v2ZGP5LWkxS9au6EAKCYBDjjUjRIu3SnRD
Tkx7xE/7G1N7nT624m5yWfb7Tkk7Wl3CU/72cTq9AcHgcwoeLHPsB3Dsl74uO0n1
dKwP0qZUpqN9JB2mdk9mGTfTdEByu3zqgAVXozmhzIPTOH/XlM2SNRE5LhI0NXbQ
z99u5wMvw2JUHamqiEg/sO1m2NdCr84PS3emjeRIsFj4eSaww7LJwY3s074vNGWT
iy3YRS/oCaTamFY6rTKOBw+s8TcB1jQClE9zMFkVcKa0TPrqOmeeAEuLhIqYEzIp
Eeua0ANr2Ya5tEJWF2ayXarinINrcFQmHzg/3f+QZFYTOXKqfaN64OSaCn1EOiSC
aRGptOm5ZViEiD4jVByDnysdRsNFpW6Eq3kw2vGzH7mvZjQku0pWX4AcOZxvVKVE
K5FoiQhs3Ib7x6/Nhv8XjwGda2sUrs4tmuQzjTn+lERJSxV+e/jj2rhZ2dG8OduV
pScAeDJiyPrKLL5dP4YvS+IbtdB3HnYLjYf1WxJzRcKq4rbogLTXGgHjgWrdcfgd
aVa1EdobeJMZOgRUBH705ZjoaVyxc2gwhb5DBdNlzfk35i8Qyjwj2KwIpkMcwRDJ
64KK8j0iMj12oAza0F9nXouLGexxIpQQjyx3JPPEHCY6Wk/51or/1J4/Ajiyxi6d
3hezNPEb/J/bwRU/z/QNKnDkIk+8vl5GtBAn1YiKP7EsXEbVSf5uVM+FBSyOkxsl
0JneYR21Iv6XDY9LBgaMfvZ67QHr7Q6CaLf0A4jWvmSiCW7Gdhz5FrHvxQwci1/x
88Q7jE/1UotvKxF0bsLgxybTy6KZMPgoIvX4Mb1ZRRO774qRX0OYCK7DKCOphmLu
Y3ulFP8irRejnc14xFAo+Qx0DjZO8Wiz8neQl+j/8+dftoUtHnIXaL+RawEDSjyu
Ax/OgXAZWOm7veqvH49okQzAZQgzmOXCPxjAkNXeemGzcWphA05gix6yr2GQH2jU
JufLPO3Ku3o5P8w/9S0ZjtMbP0Gn2p42vyJ5x41HPcdUoPqrVc2LLJtxd7CFAcur
4q5v711lTW4bXksyBP9/qDiznLzQ4z6tESLUt76mHqh9VWgXO7gceUGQDbZ+USnM
Esdv22wGiJNQmTty0CGMb0PZbJOIxXjbbEjFarcCe/JK39TK4madcv2Hs8lA6aRM
HDlM08dBVpXOQHSDsDcqVhM8BLFoibpNjbES0sEY1FWAFMINwMJzwzGLIlL+n0ib
JKiqYtqOzuMO2j02mhiFRsusmos5z8fUyYXiHahgJu8oPWSiVMFV4O0BmonAptE0
fI0457vj3sqhvvFjlqvzQm/L/eu/9VaRpb6CQ8lnrY4eb4Zk8vAZSP4LfiZPLtXj
ST8qv4C3bb6DhZaUscalnfp/ZWJGmhtQJGsE1dpg+IZI7sB4k9qBT1PiM8BzQITf
ByL73bGL3FusYAlvmMX6sPulo/nGGvRoOUKjzxlPK8pdnGg/s8rmqRXJDOfjt2zK
xk+fjy+7ytOnCS/tQUEVCbaf1RHw1xmrW6uDJY+TYU7LnY+4IAbrSe+PGNky2AbF
KQbi0xnRRrpe73rB6DxDUqZPqJLzqKOaYtimQOvyLiMDtFn2d8n0iPK4K8PwIYGh
dVRw8977i/v0y5mSEfh8MnP8gbKc95wJlhQ4iBjhKXPdndoecAKmspAyan5hzfN6
/bKW63I0wbVshuwrRyQWk1c0DjX8h7eSeMySWY7HatCpMCzDp3Fq5976LKQOR2PA
7RxGZ4oxXq55kK6nE5fWxLa7Nco8bqlD4jRZlR4cr53qFGQTy3NdQyVd5/a/I1Rr
GHPeVJHSSpLLXXggENLhROp/T7UKHBvylFWBF22HgQg5n/+zt6IimSyzmgsKTaKo
gfTbfmixGNeFmcR9NOfcbJDtLMlEtV7siSsswxamcekO56hgJe66ZrtEArhGE3Wn
qMTeEbdjOSxz9ip+YLw/JmRvUEqsqcNXR8P1V8h3wvrYJN+5rGnz9YcR+rSbreaS
FBtL3o4nH5igRNk8jjIU+Q8b57zCJTG38ER+TLLg0o8krWRqG88Art6XStMQ3jTq
Ifn2jdXVrnIJ5KfYBf8d3cC81OCpIv7KL+pKok6Ps0ZSBjsX430cUsoaza8+w1wn
MnBqSRWSK4X2p0rPOfQZSkNSZa4R2GyoFn7qe7tJFB+IQ+kO1je+0G9h83MN78xO
1XxMihYcP6gdl3i4flzL2WiWGINTkV1udnKtnuNeKKK/1bt3yLhyWSPuSVqEJmuu
emjKvlLhnkENh1aECF227diN0CVq/Im5rMST0YktyXwvwQkTfQQyi2YUU5IIftKh
jvMRbxkQsD+cEzdBJVATZxKL9GMTi4ROldlCe2YjsxVxL9ecCKeIPs22YYskte5H
wabL/+R3TT+ANOs0byBI/s8Ptr7wIRGpqcW+93l7b/Hw3TXRJuVjekG8Wf012LSy
Pm8aaJE92lpGLhM+QRja7t8LQjZCuiSZkdN3crfxOh6q49ALJaQ8UkCnIqKK4/a8
PINC0LP6X3NHisMSClQNDoyEUb4KRSWVSfShI6QtXheUM+NtvR/sDfosYBbVkatP
2Qg7uMAFA6W5pVj5ED18u6FOJ2rlUmHwnKzOVX0D9FtvLrtnrsgP3wo4+4l8hijO
KiEfBtmqGCkFkKJudw8vpKHnO7xn5t1OVtmLDHKnw7NgYjDgpxh+2QGKAZscaVQp
tBjgq82wTnDTFEeAux+5weUmgYZIkfHPL1/cDJUp3pjHotgZ9TBgs6/0FhIyeCPL
G+4r0nQb9fHKIRhYHXUEkR75CMkSwq9NWtBh1qJUiMSKqDnMEABxzaiXkI/P7hw0
fvIqAWCLx1bObU8oPyHYfozN4Qicl19+SqZG8bNKxDoych0QzvN0CmIbl2Ly6K3K
SRVUIrXuJ6YCP029OkbLW65wrd5AmqRS6maG/CErO0CY6+4eXa2j5x89mVXL2gvu
REY+hjgxVSguZUmn1gK+ESoccOoUSrR5S3VBNgQj5E1cbh6yIMkvzDmhJOP65Wih
NWLXpuKgk71J7TrxK/pd5xzpRhnn8sGFCoif79DCqTQXzGtNynk0IlPvlppHTHaK
DEgBGq8vMqpjIWvT3zbgeEI6tYdqjTm0BdGUL9NtoStLrZr543DxSJw0HLXn6PN5
W2fGTdVm08yGo5/yov3xmFDqE3Nn6jk7+fo7Etao/qQqNIN2CBjbPZZvHRgGPFgz
RjjhxHzkOz2IqGRVaM2NUKCZfBB7O9OfGEjOpzt29CQ0FJztMluwliCKPKmT4iFp
eTEhnW423w3eKGaZhYzBo3ht3SHG26oex9FY8/QUTxznaoeJ3cFAOLXNtLN1KuI6
bBd1yRVtwuyRhZ4/8ReS18+iYiFzxSpSKw586kYgIFMZLAgftna8fBjjgJ4UpFC1
pknA5Rr7iI20n7CcojDXabGwVzBRNQwnGhQSYzl0+F+d1VHcJQd71swB11l/Sntk
INtf2sd8TKamA+xAm5ZAYfKVsNw4KmrDkJpkm+ggqFZC3rTrd0VJt32Gz6Bbr/sF
jxGCSfqp9ZjZwaXGNLC+BIkT3ZIaLuq6V6d5U6m178lh3VKu6exFc6xnc1YkOoLK
CtUlirDetMx6D8XjWWxyn4tikdTwmXwerOS0DGHl1SD8mHJumXP4d1BhQZ61QwQD
0ShhoF5RPiOwefXlIn12dkHShUo1vpnKosTXuPJmI7OBYdluyrfnVZl1qmr3kXRY
g1hWbhFCDkMZ405/vMhXKjVn97pLN0bGTr8w88Z883lPGG9XZwfOblQIs6hvIMz1
pf9+FSaFPGxuAx6M2Wis0a7/0RI2qLb/HmDIrSGA8TAyROifrFDHUBHxuMPH+F8/
h5oU+DB3OjYCvF4dmdvj7lb6n9NJAyofQCFyYSsaMefS/zw/11WgoM/dZ7TKgqyu
IO7VKPXgkXAQb/iqr0O9op2akDgO6qOYrfttuuIMi2IinyQ3UCi8AJDXJZQs0uM9
dErK4HS/ia3N6wMfj6IeB5RNeLhuUSSESILYBZiQK08Oo1wdZdqB2z9nBQ99KAGD
fyaRqSxkC2+fbu3CRz0nM6t1QsQvOI8SlB7exkIhbRJ4oEgNG9au5GlMdazdBPOn
6crWekZ8LWH4JZg3JJ4DwI1R5EuffGjl0fciE7YCEoDukKrIwKMHwA/GmUgxoLq4
mC/X+AynyJ/H4cPouUckwniUXNXbBI71BGShV1DqVqTgGvN8r2R810LbTu1L8m4F
BSOEd4NGasJ04ymRUTL5Dm9OPiSjV1YLnr2jzmllh+X4VW+dohowQALNNfTGYb0q
eQ0uM5FAU5pwfvPWkmaUccsMn2X3bkDos0HB8l4cXv296ze2zNhJ++7CIrH+8MU6
mG4uS5kEE2ZMUx+DlrZvWpmy0QrxbPz4lUcepqJma5Ncw2a3j6TM27zLvmj6Phwn
2XdHcOPigC74DW2c2yDMWhLa5htk4Yz8LfSzyZ3+iBPvIkbfYVuOhRY9GvzmLesF
KlYU7T5U1Iiduuy4tbdb5cej4wHxZXBBQNKcjQbTOgkloPKnS2/ak+gEBYp/TCQX
8oxsW2yn2DD1t/Zqc7Fk1zybi0Pg9NGBQyo1MNjHwgepFBXIWM7UreOuVKFstrO8
A0uzN/IXfJvLFqGQmunz4vqA02kd9kboKEWCXZA1bvQic7OWj7DPqzxG9lc/XL7F
aEiFBZtWjlWhdcgIE6DDsRAFwQsx8vCLUdGm+lYLqHd1x/WynnC1k5SuFmHusRMk
nHAhpwBRJgc1qjzO+eQqUPWS8yZdp/fEXPXccu5D40+vt+KhVHOosHtrF+msz7Jh
o/0OHfveypP1366U0pTgLd9ua4zNrOGevPj1hE67sugTrl44o5jhz4gAA4EH85to
dhzKu6/20lLcNVb7reXSWdOfyzwTKZtwJE98iepZzCX5HFhyJDnIjS8a7HiRSSCe
bDtMK3UljnWLeyGbIJkKjAvehb2oY4lYdZaJBs/rcysS4eLTOWrlR2GwRYI6e84P
LC6FbJNjkVRSXUmJocjEtBeJrcRF6hYHl9rsyil2UJpA4rLWevb+F1bE+65NRTEc
1MGW/il8ggDST82sgHc8nvcrreXP6VDrGYgBqzsKI4EuNBVNLGra5GFnahh4ScZ9
dxN+eqXgFHeP2snBMD+YTRg5NHiomXHFNNb0LExJIZFyGe59umTLQ3jWhmWnz8/2
PiGkpZUW5EYLDo2zPanKXYmp/+pInXIvEkGgWYpCDQ2mhWlOZ6WfLnwZg8t2GBem
FBBnkMiyB6tCbfR2gYJCeURUdGU5XXjeGr1irFh4WooEKcZj173qJJroVufI3NUo
LefipvYzDokhgogQ2nfREAOnBwt77w+8AGEnI2hzFP6RXC0chLigCMsdjfemytMi
HY9zEMGkPArAEBjEub3j3wSnMWkWv57+YVeDj0gSWDyku0wsX8SGaVk7BUYmJ2+X
K5AGZSXpCh9y+M830CBi4sCpwac7NE2sEG5QujqEaQWdWi299ulR7N2sDl5pP2/r
L1+AMQNiDdv/FIL6tCVyX8mC4g7WTsNP2RAoYKT1n+9WRE+vCbx7ujDpemAzA1YQ
V0RwfgVVMd6SC91s5DfO9obaQzmdJ7+xgn51q5gS5kHzHRG4P27k39+gMF9XhD8Q
kQ6S0svnT0jhjdfBfZ3ln1NZ78C7048WSCQ+m1zwaqp1eWUwNGhPglVra+oKjfdH
1bxIKT/VE2s0kJEJ5QWhOB06x72vtiI+bglH3E/xDwwUEGtIkLSCxSjyRUAV8zan
i7wjpguTYBp0zIZ9vXju3x5uTfkGuGoe5O9kRu+ZKfx3hjObB8vu5p/PxJk5hbbf
wwxAkkrrw3LIkGFT3Nv6gL/jvRX5pGlT/G25o9RndPbHWO9M4z3xcORnpEiaUR3h
cCx8pLxNmuEktAceSTwqSPBoTuYdT1xQ7Z68goKFbvvCfCt2VTxfzPMJUlzTWm55
KoWw11RHEdQUcWfOH5msf3PJvfrAhn3GAs6y2jPf1iXeqPrl4vvbzAtg6q423lmY
JN+zLjV0fX3iS8tr2uWgwB75Zuh5pcTGXCfIauiPLdjjNwOZ5V3K5kEEfahCvLVM
OOhmQTBgfZge4+7Dz5i9T5CBoYLe2dSraPP8PhM1Z2z6HZllDHDBQCeibm+RRClB
+neK8o3ueIs/pHzbTNCdzvCOPzZbE5DIz+dmPYRKGZrxexvMn3jhtsP/h2VnGWTB
PHIQMD0PCNMQJe47exrY0HaNz81iKe/nKqHlIMT/UUnuGBmaT8G06L4mB6bfwvKT
/ezUhye+17JRvF5upvE1kp3ZtU1GSKLGAwdPE86yhEXYP6VPVt+eX5Ap7MbrWQ1t
0OufvEvNnEIrsOW4aGd4Gm32f6a+MESOSuRklnO6OtavsDPYnW/WIvod8s06Iuy8
uyg6o2lkvxbvO8dGIDWaXMgmgWngdvvefW5UxFX088DslJ6jAqmtJxpqSFcBjISL
VcRrOqBkaWFGtc7nm2uhFvKW/ra38CvsCyyvY4jjGdOD89xjHCkh70i1WvumrkSv
EiveOYYU/FljwAoRr7/U2HnzRFH3/xyLj519C13lWnmRfVY9K8k2Na6NdZCc1zD+
4n4txO2CUvRvxIiNFi7Ryo0dvHlgl9+XoqWIMOVpg8EyOBgMDnBtDavWX3UUczJQ
m7OHI4TVu06yeZ88CG3t65gNVlLYtjPYSxbiSqc7JqLTDgU0yhtKIJgVcM54BjfS
W1cqCW/JxgC9p4rGPdM7cxuUBBdRbiGVBqLW+cFpdX6bikr43sxG/ffdB4Z8klAv
bHR1GjuBuytvGnSaR0QzcAQZHyp+nSZXdAhXI/ZXWfp8bXED2MOefj/or+O0Aexb
QUlTCRUcFEvQY9aQsSuFgTDEq5iEeMCi64JnM8VBks5uzIHUeLDrzbty8gyzGFq/
rzhQgu4zYGal6h/GQ8w9ocUW1a3ih4kj7hVtuCqGIRgixkFwi20vbMgKhslzidPm
1EA4VRFBDcq/vuyOZty3G1K1SF9uPkvrOEEsEjeqmZhjmwu1YMqvG2ffgWNB8ZJo
oZEXQ798UNDi1jKn4ej7Ot/kKGCVGioaC9j9ucuLg3LjtXQsRDrr6murFwpEQLo9
K9sdLybC/Zp96NIU5i6TndSPwFrJ/uxxJO2QZ0XUSnbUR5rGmGsa7/0b6B2V2d5V
2mPAxkKQR1Juoe8OUL2ac5POPXj3gPFWZBArBLGqxsz4WoqEAbbj7ueMg1uDMtCS
/U2yNUIBVWsust1+JvvUD1z6FWLArOi1U80W6EV0U8+u/BDK2tTnjBEvBCYxgmr4
h1pMwmm4LeAJ55wLzW3TXuwfB+rjH+DQeMQXqNOSP3KlJ3osl42ANfi1TuNBjr1j
BEqlLAzqLnJKibudOMEXHEL4Dpa1PN/xDeFQxuTh+OpBhkrPX6Eb1gW6VsL/mMWW
4f7yKlNCAq2HkJUgON3em6WNpTnBUOIjvFNsYspG5vGp4Lh+VQw2FN1b60JgRz+f
u2iMrrL+Bhlk5KMZ4WdJIC6qGoCM+MTYJKmcXetAwGL4Ylv2Kc4lCmmo6SyOF1vI
HmBDDrPktjxLVcXTBaBvte2QxjoEzBXN6hCArVPyRmJjXFJAPMIBScPo3UX9eAjW
6wLMRJgLZw0585ze3qtFnkyy+h4P1frUQMko8cV+nAqCrZlNJnBznzqOZeJxnajU
Oft2XRVf1oIUjtpxTlVJn1KVIyhjayKg2XLaIjTP8ZIZT05mnjmNOjxKbelTEQ72
ACW/lk5q9q9yhyuVeAQLxbCF9PT7BUp2UWWd1cX+J2FHEuyjcjF1al8Ew9hg+Xvk
qqDbc3e3mReejxHlgYYljy7EilfGMHeKtesR6KSpJOApUcHkQmr5TaitFWl6SH4n
KtbvGJlTqr6mO9KJ/gTWCfrzttfaN5GvAWOGUP+0qphYSpALhcUlQnNvjkWJddb5
Yxwy7ZXvzOJNddkd5BKQsRuz5USva/uVCMqoyj363uyyQts8/Bg1Y+hyy5kUm+NR
9uaGzadrsY4xFL/WW6u8PCnDTW+Yhr/u9Ab0M8cCCZFIkwylSdCz/nybvrg9720Z
E2/aUsi2Jfnu7YpQ7rThbvhcqk+D/RXL/VxBaxt1Ba6q62Pjlq5QkWRHe/LPY+fl
x0/wNFjIE07V+sNhl+bZ9Ykcdmi6TCQ6ccxJNYb8sHQ1iOo89tDcXLc/W4BEWdlG
AreATAe0N6iwPY7LOUArOU606YetZ4fs+fzV1XiAEdkcMsjZ06RYRIEa2+M2Kt1b
KZLQJPkn9ANfZ1+yhuGFee04A561Pr92/hoGgGVuoyXUWOL93tJY94AK/3tzCPBJ
HWHqhViplthr4SsTzsqizmVS3Nyki2jK+ptsIvxip3r7GdcG1LqxvFoG+q7f9WyG
9d/Ze9LHkCXrqufv95/29ewwyfxs43N98WtpHehXPfJzHuCduWVqFWOgWCbIpP1I
5Zh/Xko/HcXucMgb5r+XaNG5V/1PmnwAb2bk8F0YtFLBDH7W2nOj7w+tsdeci+SO
fnVQxbYtbHDyWK4wJpSpGLBuquELU9VSZotTGSRSeYWfs16iWvK1nVjb1Q0cA5Tx
UOb7ZyhS+7d16z2zK2e988f2AUgPPhsXaMhjwH8H9IvjOaMouA8Ice8/j6iUa6Z0
d0swifHB0w/+h///L0Aq+T25WApCk08R+lN90Tv2L5sTpL+jZQRbNhlm0tZQ/rfU
PdOrgizLx+bG4ztyajCPTjagupfcD9OvALUjck11zVcjoHnHt7mkwiMmqdq5kf7h
aADiEEHB+fFNk7R4GOONzEQoH4D18fPIqU1chtherjDaI7lWi9oz0wVshBzwCjkC
vHSDPrNsRrmZDlTNO+PI+fES/e6IRsxa0l1nztmWMQtmHF32hHKdMXAo840MkvBt
QlR3WfzFQLcyblFXoYcuAFbqNdfwvpEmO5emvXREq/2xImAq9+LpBqjixkIlCs68
ngsC1/ElpMOcXijHjfCcbzxklakLyQhQQ74TB1xFdfAj43qZRrdXm04DLwXyH3Os
AdLCglqAtQqDc7Edee7wS2tx9RZXTlZaHKfqhDF0pNHKPy8jd3eVaK2q4hIB8Y3H
WDF1J9qC72m2lQNVef6MpvLV7C0IcM8PFjsVRgQfDZogBGyrU+rAcYZPwA7zw6X0
+iMdmKXrgzPydddkGC0id65a3huHsGpcykhxcM5ypq2yMOuJmupOvUlZY3L0pg90
dNa5qk7qD1dQymH+x/Te1vrvKEHXGBIo+urPAlV4rZBTrzhruqggDwQ3wunBuj4k
wfs1QNsSi2fI2/XcAeNXk77WhmsWHk1z7IRLSgWrWVASYyue7btQNaxmZCKDs7sw
FIb/HfZ6NQdI/YV4BpHjQTmls2GAaqUeSoiHHSsJmdSaNULMCbBnscuDGfXX5nJA
cbtsJjXvba4tRWmEusFINy28R7fsUEQAQxAaDV745uWYsCCL8S5CzobbAElNE/Tl
a0shJxfcFpFaL72Sn3+9uwl45ElWFcoJRaHTdJ6/f3tAZjLObx/Fw4f/lEflBEuD
ajiG/1jhiw9HNuemV+T6fuS2zt+vNfp+cx5SBVNRPnTBVd4hht5TRjF1SP64aY7Y
vYS+ID+xYnFavHPv3PKQ3V3W4Ki0/NYTVBiAJ+rxm0fWfnK0E6VB7P9UgNToEg6S
/zXj/UZDVsiv1BWQp1g8H+eg/61pEvHNO0YcmdCqzTecQiZrFqgTbeleW2fNgUlk
BfBQL0/eKzl2mdPeYrVMvoXgAeoCkOeg0vF7i1K8s84hVgBBVZZcKial/5Wc/MPO
OgH47N074PRJ51dScbNjkwK5rKdmwLb4knA0dXhqH/AZEmvWuSZZMl4vI/46YyKS
cS/5rGdIV4N27c2BKtrgsoL3qShYVpILew/M1caRIHk9fUbRrG/lxqE45vhqqGKm
/yrPnpiYA++xQZU7QUpf9pBXoVkc98KyH+0WJIF7c10UyR9fcVskJReqn8EwtANw
L031Kq1WvK5Cbz0HGI0BCG6fTKtseTykN+axvebY46SiiLN52rGpRaZCb89PmpY3
9IajXJxrMKegeiKqhWzDQLcqOF2BaIOgAnjOR/oH3ARPdKxpcV8pNydBcaAJB1g9
q/NURKYV4a6XgFc19aKf05y1t4vNNJqbfqoTI3S3inN74yzLJI85BWwcnVAxO2M5
biXxtvSNCu4xL7apK/V8hUkXqREgqcOZABnpIVG6tM2s3wIqakJXyJJyoUGC5Hn4
7pWERDVZrP/ys7Ae8TDQr1nq/twJAV5ASxjSJoDTtWt8+ruOQhoU8xoyOUVILgq2
Bk4PnIOgEMATjU/+StCTaB+DWB4fplDSguLGstDTF5aW7WPQgXLi5Q7fsanWLEgj
mv3oRuzVbfvVyUQcxtMAdAsN1nRLWru6bPZNza8whNAtZ3mnV8y/4+Uu2pgr60xe
ZMTDtSonVc3AXmMRBTNh3/n/qQ9hdB1gAHNgzwDGv5lxxz1M6trlkibFaXd9JdmE
BWoZrVla7Os4l+tBEpWKR8INbIKywUeziwkzucD6t2HxyGLeojdlWTac8J4B2GQN
PyFCo276ZWi5wpS1y6HDXl6VTzzvHxIb83/x4AB0cU9Y+wyjRKrDK3O/EkhjyKHb
V+ejk3D/+eq2LTCB2tpIuaSwMIR0x2jRVX6pl63VrHavuZIh+IknR2q+mJWjk+Wp
KFAhFsJcqAjbEhJ/zoPVpuY0/Xz3WmcHgCNRv98GNdB6bGTcPMZtXybVgVtgKQGC
C2WEhN/jTTsQhysF88V5e1Qke/n9Fk7xqDzzPAzjB66Aah8KY5cDj0gfNPbz/wpM
z1o0Yr5KJyOvJfRhx0mDYOJHUgOw3twhh0u+Rr+GDFBD07hyJoe71RAR3xFCYmqX
AdwE9kSn5Y2jix/8prFYueS2y6Y/89u446sguYJG5H4i9nhj8lRLPH9pYppj6ZiM
NQCoH80YQ3koCDP39HS+PAzusyErKyzmCPQ5UujgtUuqgPtjm6BV0fkIuVssULne
jClXiMpgfOuc4whmJjt0jI9citItvj0l/6aTjSUs4GL1R/X13GoECQCgWbh+kbbB
V5vh1XWoGH96D8uuKztLHi7YctX5HabsWPGT3C4NJmKAfDcIswjr0eiDaCD0RWTe
+Pmd3poAJNnPhfZ88UcbO4PdzHPd6Pyp7iJOP+AeH+WZHOCTR2TPUl7MaPK6WlQK
Fecz3YZfX3AtpB3N0nb1ysxb4gQEVUZoTAVC5FGj5lm4lfdKae/aHy9RGe6YH0Fp
5GD+oiUiD/N1nFz2RYJs2RBtjWvy+KCIoEu9HITnguyWFLHTRTafmrzoeAVWAnq8
cQ83vbeQDPj/+kwbUdVaGdkcXSol3llnhoNwHufl/e0W5uFd/uwykgpJQ+ZO9AZQ
ETghVn1CQVOPp9RuC2uNQJTAnasYbbNiyUVcR2OryW5SmBGOZljWAl7iDCF7sZXo
AKNoLcC16kI9+32Jzb5s4pR55r+NJgBByzPO4InPZfLsaLXNcoMm2/TbPyNCScYA
POHmbtGk998LQfnx9d2fgAv7Cf9VVkEU2PVThTHI7zEvvGYEi6hqcouPJYk4Vfby
BjK22k5pHEqVSYz7QM/f9ER+5GyxYLwyZcxc79K5eCjFqqG1Q1RvskjGA6HnvI8P
nGgbvaNhe3OCxDiiITsStScEnMfiSHEuHRCWyglMCs7r73F/Y1Wy+kqudcOacpju
G/8V2k3vRWxeZCzWJgJioNpYG50g37C7IzS86kI5IYJbW/CKHuOAPUZNjuKbrGHL
q4PqBEyudd2nEUhIb+HtCwinLyPnbnCkkfwyr7XqRPoRuU1al8J3Frn0Cm1oDoDY
0A/riErLAbRhhtyKvwK9o68S7LG3PAnst18Q1cvA6fQZYnCoczrFNNOFFMzvnFKc
S+TZLaaQ35kXXHYPhcfoBsDacI9ymPDNFLndQ5K4a7/AYWeTV+KmwNhBWVGsx2Oc
XzPmdoyteqGcrJXn8O68A1b//3hdUrzquzj6uGujGjHlfKr7eqUDTjmaF/LqFD8v
ZXnG5Qg+qWcpMIlsfaPR5JNbYgaS1WP0hrgGbsLyOic+fY+qWU4xZLZqHNWNGI/Z
UDaeM59Vp8EwTicpbn3HY2s6IUIttavyPAbNJS5WoShOX9UB7ICbU41O2ACvFhCd
5/WQxp3wy/T+FnznXOIfXdEtRO0Rb/fVvvLDWTOctqaXnv9q/o4Cd1sktDlOzgdU
YkL34+OUnLBSGRSZsok6MYc6y5tJ6mCLaxgrg7TFOkWcNHKLRajhB1hj9gX4TWH+
YibZhRYv06sArReqIeSnh9roAiy9EpSwvvoATLB/pW93wN1VC2a+C7wMPNF+EP6f
f6l5c8SlqvmcJG5Z9962EoGHPFY4w13gBuLzy3Eqv2J/R9CVMn/Zc6khTDBcbQTA
pgg3ObDJ9/Lqwq8pn2pR7wEf3qZ6ZpaWBYDqV29CH1SVpxUqXVqvoUQUFCoVotbG
9/2Vb16xrDiZLWuqFkrx2+rxIS92tcrIBUMxuUm7OA98NEQNEWSghGjvBr+rI6fu
uzqJDH088JXAfgkK/uNrxmwYNQoiAQYtg6HEY1efPbcDD3upExL51VM5Dk8ul8iW
0HP+VquteXcWQTt3nPFG/2ZKEQe7sJ2GXHlp6QXJOKQDggOjOPYmFTQOlKtbFGSP
R4pXP+zC5INK91wFGuVuQKX9LgV2a1W42XHrgqms5D04yxPsHLjweBwwYcdmC9la
WhkFMOYZYnjR7P6okZ2P8iub8+Kfuk8WQGTQuYRWPgH/JHlqQfTI26WQk6Y3jRBa
xWaVJLnNGus988WCkXdASeXjny9k+9rW6fyz4Tac1qP54nAfJ9frOGktUI56y9d4
RU9zGZEdgt2MGaJX8WHtmPd2xBirIvKeIFHnBXkrTk0lA69jI0aTkQQ2/4+BNOxS
CakRDoo+wsubWNJUwcPcyz9KNV+fsBiRKpaKF0Ra23kT9egeGD06oELNfQyU5Knd
DxR48aJARiDmIp9ikBhajrvWHZGBPTdLJBmnAs3jO5G8Mhr46GMo+nIljt3iKLeg
aCyEa5DrK7DsK9dhP7LybZvreLIaiEJdTATMz/6HFyjaCOxIeFU0K3z77M7Y6Z81
lCNLsXzATTf9tytXrpeS5/yVpybR9zoyTdUpeVMaBwg6eRSNwJGdtJTaq9lZiKFZ
aAd5F7F6Ncy4e1H/qjvSPjYr3PqUpy8hqYBV6ZycKjAmHKT3CCVu5VkpibbzWFKH
fAXF3xP8ixcEPQSXFCL7b/rVcW3sbJs6s178rA/oKsU7mvzSnmol6O9bmTPX5Idv
8q+UspS2I21u1wr+7ON6rTu4PpLgSAiEF3WC3S3R86f2oMh2mS0xKzwf6idwBSJf
Vyyunicvmpi+fnmI5jtxYHVAn3MnUVe22EHJKSl0eBzl4zoDScb0ugM5UX4ohkJg
v+LLvHW1t/CffvxflTo6oC/I5WPiTnaB/OPJ7tha0SNlDFsPyfE0MZ4CrMnocoGQ
rv/bJXEVF1tV2UqEc+/arm+8Au0yFVkCJ83eq/0a9/rg9hO17TwvgjteMonMtycA
cE2HQeYPm6Qws/FuOFW8tXYFV6pwsAH53KLNWadPO4a+BdnLU9XL2cy6vCv8xyo7
OZD7nFSOdQif90+wo/+c7zdJrthdmAT+I50zsqmEAKVxlkbhfw8kzK4Bsc415llF
ALf5qsxGxQf2yR5T5LldDoRfAMxFMsLPF94+vlwLaAAna92qaN2n1g8FFx0HmL57
0AcPNbB7iedXErbgEnCdPd6eScci/lJ7VUO/EgaEpFFbMrHgo/hhOsoYrhQkj/ww
smoTNOKkjGHHNG4yB9AKBKHzeW9/jn81p+E6yVEbTxf6u5pProjEHsHFu5n8yn0l
oWYyOqGj1Nhzc5T1GdlGKVKnuMjQMLfdmiNdTkj4qT8pseTtVf1SvrOGTwJkxVJ3
ymerWUrVNnKc36Db6yA+r/DYFFZspPymsXkGF6uoq2QhobkksY0h4A6pzC2eehdB
cUIlZ3ghP9e2SuekwEEzNx8RILxIiW+QbS5485UOkzQ2Y+y5NHmYAIb7v8yVJFRN
/6YwsvddyMpXHUKJWoKhwnebdO7B+zyXq+Z6ddlExDbC+KGB9+4Df/7QlQRFspje
1lASv5vDfMvEI+ceq8h06PtlT5iLQ2HcO707w38ORu4MAHhVyChiZoX+9K9MPxCx
1j9XpDKQJNYXJl2Dj+mboqkht9cid7JcN66N3rhTN+mibZnYICMYseXAz7vmp+xT
d4/bPL2Hr8nkY6FPlfEseMBgn2PuI2pgjMwpCpeyD7HybP2VIYqsAGzMN9Xnd8im
aI4uWRMG7qICntvrWjsdNgKMeDGcJko6jC3++99Pc5vSi4gNHkChH+x7FMh7AxXY
PpQFFBS1tmLzjrrG8+1jLalAAo5tDffZKWnhwXebvQesg+acbc9dJsE/s2xVnG68
qEAtgIMXwCxnkKhruq9+OhAL592OQ8rL0JTeCbUY+Lz9sq49q87/14tjZ4Y7Qnuk
Wl40tPp5Y1aL8J351ummyWnvq80EFTksoK+gA22kejTdLOxLYR8KbG4WCYTMTow0
vu+HMyR+WsWNVrkyUhgfOVhKq4Mo22Ebw996vev/2LE9cDNyabL8/eKNaUbclhko
DUoIoEN5L5CFQvlLFN15A3XOTrCOZanvCDDEK0deXYSutbTW2H3EYpx6CDnpOG3K
ChEQyO7zjBRivIwvM6I86Jvu2r02vfaKA1OxZhOK4qlGvTi6JXYu+xdvI1043ki9
IfFIUpWQBcZEzodKKITbmktaBhfAP0KL7z14uHfSx50Qg993XpFrIdezKWMja/HX
S1zVsMLR3RpzrxtJXhZzH5m2YD62Pja7IMIcQrnjOIEkcYqKiBl+DSH//26pSxLr
4syHMwxw7bxhUG3VrzyzLrvqaX8dFlEu+0+E5u6cktUqj5ytB8MyN3npbWKWJWjn
YMr5wFLPMlC52yHqeMVTuTlfFI9mHPktNfHi7PlSkg7OPW2Nw/wDvWqlzLusZEUx
bfwXelgBRjW6sxuEXyigB4GAxLYhAzzYXPIxy7TRALPU3+e7Y+hhOsEOcZEKBrx+
l+jjFnoFrTzz7i/agybGzsE1dNct7C3YoEW84eBXIhbn+uUSebnZ7aveQZnKeS+N
w2lQj3HvO2Ol6aNkJT58QHjjN1/g6nVTO7bV0H6d5Ef0oQ6Q/NJrZW0PbEU2Fg51
FEKKrFUGPGBNMQx4CIxSiavspzCm7qnyc5nNZSOI3QekO5eZSmVCeJ5f+suOwTry
24znATXZmdibxJrwB8iE1sjtJDM51U6DZWEPB+dEcEqQjUIiJvtGuVjie2vGm57G
auxQ6VDdAdqVa6solzcoVYAT6yWHQtDACeODfkAnj6lbSQpkxFqq2EaLr5YYgtmI
iQjd1xVLlu04zT8MKeqGpi5hoCVW0iSQiKEPLdxYjkRpOOacZVlV1NA65H7LsXWd
Ahw92dUeyVtLyTvc+PjsVaeLBo8NYaT4/yMzw9O+Op0huUN253xEZeryMMeeOaLT
1DlbW3+NPgn/h88NsJLJ8Ri3rYkHx0gIFtpEAb8MAJgCoouVRwCD6fUL63ZjUfAO
u25aUv7e9c74JkI5a3+12k9vnE39c8BIJq4epBOmBrdWQ+uYpF7d83GaSUKLJ46B
fLBHKHH/XC952+5dlQhzR8rXgBsKGO83LP4ngaunvt5+8JCI/23o9cSrwUPpoyHi
ej1H4VqA3BVFNFGLnLy1l7A11Ra7EbUWwfuMs6mXytTjLFLaAgm7ny29KB7U5dJN
Qd8SSyLHL04EQcy+KCAONh2Ui7UnVKjUBSSUWaEO69z5TaS6P+hWzoTP0iWz5l6u
9eiADWEUEfw5u9xt4vJplslHLb9B8SNUnpPKtGZihDWjOLabV+1WMylkGzdnRyyz
MrM6bPn2PX8ETcE4d1IqQtexkkoy+67NuJWP8IDnpBP6ere0IpyI/O0ZKTf0/+oA
nUKKGAgdwOchkoy5rufWeqHqL8JvHq7ViVpNGf5xJ7aelEbY7cNEYxUE2vzlpxbw
5GZZk/jZXdRd1cZITnt7sgftjlqGxvAu4ITYYMj7pZ0eKWWJERI80b/j0/nGHnq2
LsgSmQ64TXSW09cTLkhOnIW6bGEiZKluY2KR+5el+Mb7+uWKXNTdFNp6d6JIURoW
Z21R6z9YdOFCYZrxXkwfQ7/YiYht/NTg78mA3rfNNWyt9uz1Fz7lWbvoU6nQWf6L
tbxUZtEeIzxbPZFwc7q33q3k7qm2DL7i/9tAHIJ52e+AUpIWotm1v1vxx2YsYNmg
CsLTIYI8I0kqcYfdERd4QT+7IlyKwbjGUS6XR8VkHDY/b3a0L9yPMcDkmdeQmoRM
3a0pyua3viN2L2wu3YQY7gtUwN0bQKfKpzLAoyYxHt7SZvkwxwFhyM26hQHj5tK7
jCqTkC6aJF7OpShj7BBljd2nhRS6VKfijsitMDiZWy2E7h70AQsllBJGXUOaSKuV
Ha7W7YA6oNFEaTHukuQ28sEo3sRts77sp+dDtXrVTkBuGPQPAlxiGDvtDO1jvP3B
SbQd1G/slxqsHfqqlOHFCkbDMLq8og52LuMN4GPjDX2fMW7SZe0lamkVWd34gmxB
85F0Bs4taeAfNCFQ9jGoQN1TeZ8+ZejoxoDVJty8pKXJkJ9abEZOhVPNt7LZUhW9
ngQYaH6cVLmSXPOMc6rjTaFfdVjLCC/0fISgPrx55BZIwMcwI+pV8YjA+0maudas
DUaN+T93FF++jLKykLKAc1A7gOPtWGkXwvau00c9kiwCJt2314YUfxQBwvnHIlDO
oOJbu5yZPC18uyxNuLdjWGTvzrmMnjJLKkBNOo4P+URLuHMbCBEKrExGlEJuMw/g
fEIVNWoeYar8s9YHB7Jc7t8UoXrdUXfKR+HckY32gLUcAldXrKrE0CB22OoUUXoc
bsJqih6hglwmXLnv5mko+AtqGtIcMf7cKQyLlfghD5xSTUK2s51ye8fHuOuzzD1f
ZnfulP2bvI5Lju0KCktFfMH1Sdk5b0fhbt4U29VlyleHmi9P86Hf0T1ZwJ4eeYj0
RO+GkNDaqk8awEZYefPmOtQM63Sn4Ot5LWtkB7dbpMkjZh0urHN3Mm8xaEo68aY0
QjFul0/CsFWGh8RaUSoPXy/kQjeG9SAMU6YB0QMkkqlkwsFF3XZ7azirj70NooFL
Fc2vZ5DR1k47mGa8aGwCkPhCo3w4MY81pe7F1YHhFMThh2dLFf6Fadu8N6PMipBr
d5y/8QWpqoGM6yk5jzLaeolEaqe4vmo/Oavm4nFt8wBB5auqM1pZX2CPJHvmx7oH
PPZbfmByTvA3u09p+/Ddu53mNUeWzc0ofLO6Ta3UmIh3VB4YYOs+9z7SJCNodqJD
NhCcGCdjv//rjReeNjxI9KzjMUHCdc9WAyGFCFkMnNKegcA1OOYqL2tybuNhg1eE
GAcoOscczkNFxtjZUFNEs0nJGIi3IaH2Oo6okft8vSn6ZAAtRjpbquVgfKWfKQHK
HxNuLMHpmfnNrPGAME7lnGxf8+jwYq56w9PxE49aZ5mOEBcTSfsYzG7FQnJedics
WIsabCANmyyi7cTzDur/Q5CBrYr9OS/No7UOgWwNgXyKFKhuH2+xI4g4HIqT4Tzg
qi2CwuPwH09iJ7+ox6fafNQ5tKplsqWfRRNy0utvcQoDPvwiMZ2R6faIG86WnO2e
jTKr2nkJCdMvbUcfCH/rHjZOMYJabkzEHnBNqpD87EqU6vH8hXZWtTjGnPOP6QIa
NvfyII/V8nVga0Qw1QJT10d1ZFlfBRxTCfeP4vUjgypgjloGmdaWBcnCCxITDYFR
/XZSBP5pIZvU7b+e9sxc3y5GAhxbA8RHaUT8wzMySPnqmr6xiZbp7mgM8w/FfO3P
jWBcZIHrYjjbVDs+PUydoDEu94XFVSqdwWt8ENeVyLSNAQxTOb7g8BBDO3NtSkMS
UmURfciTIeVNkkXW1dG/3dptkbx+LWmYGxxoQOB6rJJobBw6x70K6/t1dwa030Ow
V+ZA09rt+N+viX1JBzyIy9ukTovayCGKLnW0SuTkyd9COx7PYUbvd8uZv+um907Z
IfD4q3mN5P7fJULfzowlqfQmyukPnrojO7DJeBBZfYmHoC2vGOWUx+4+tSGU+xMG
BIG2mFRtrBr62Nc6/LpLVB1KuUZH41aFivYGMntE4cjsjL/vUtbSNyL66cKQok0C
FUwp0fZqGaFmcy4W2SnnppglZdG3x0+8LsgAJWMrbg7d3dEB9cNqy4VvhGqeVX8a
M31TYzq20h7DHo/NJNlM6EotyzJxqR1bTVzEd5PPB8QOFE8YF1gHXk1IcxIa5lkB
LFVxQajYjXKhaa7jEJFsLg2hmOxqJApwVoBWtRjVRBCfYbupvpjmvmHoFA5+tMgL
RFBwAGBe9KeV9UGImQooUvN4kKcujI1BSrzyc0goYGPTpJRobtclxsorVERen2UH
hRITr/3UjDMbbNvpPlHfAZ8wgulf3QpvpQ03cydJOeHAX5CqkOLvzujSPCDMwXuu
lyRGHPhJk9TaaaYIq/01W/G4YvDGit2HU+VU2emapxhSe1qO2bJxS486P4OEwa7a
3Tj4mT69ngkR/lgeqFxHoRmKZ9WYYhy2Pixh1/YNgpLcRAshOiyK9n998oNYvpJe
sUr0G7ZYH/5TeLCwV4roGXHOMQzldtzT3WXvKSKCwmtNCAiZmKnkHcQ6zXAJTPhw
5fT7FCofxqDJNyin607SS/YvxVaIA1IMLGAY0XwI65+F2zv67Yfs+UjK6CixQwtE
5FKMmkoHMZw+7xc4x6eQE8McCyFS/Vg50mvZC4Iu7cbcai0kirqq9//CADdMDesf
uyRbRJa4FpZWxj/MWRi8JtVLfDrIzjf5OobWefow9q65yIGngHPQB1KDahcsOUms
EXsgZBgIHerpsro2AVn7/FIIbprh4oQM+a4TmcgPgRHIhKcopb9aLTvt6uq5WAc3
VWm9bzGs+YGRKTaDAoOSCmVK7zvJ24SsoLc4XfkXw+Kvc0skv5Z///Kzxsze0A40
NQpfw/a82QRZCLrruVjN8ao2hkKwWQTIYCwICoBXm8itZL05K/paEjqYpVjhG0re
4FxmlMaccDD1hQh2ZKMTM7XvNvCPOYaiCsdUcb6o4RpEMPnBs47/07G5INXeMSZ9
7ioiPNh34toVEA/XniUlWVk9kptPDm2znibG2cSuqrVYqZXGrQOHNSCIiCKwt2tI
6kQIVGLaTFGg3BaEz+9ozdwkKMmAmivIZHCuuITa6JQp5vQNcd0bMvNkpVUT4y+D
oaakhqhrRBuCr7eEuWQBUWd/H6CDsRvOUpbIpNaxxU+twgFiP+2VonvwcOzykgXL
RtZIiWZ44NUrBFsoZx4/N5E4+kbUVRoiAOMX3wLN8hlpSAszQ+ha1C5BEVlk7s0e
SRi5PP+JYin9ZBaqqpOBWMara8TScc/fqYLWbho2P6PCqQV43hyT1r0/Xou3FEy4
7BqDPbsa7haxe8kQEITU9QPFmVbUZlxahd0I32FKtts6cjIkNAfNa9HSyqDPjKCG
O/BE0vD7UCJGlALlR+zpx+QqDTKKy/wJzyedL/sI6o6PFEzv0YXbVBlply50C7xq
vW6pXcGXFgl6c18uZPc+RdmE5Dzt2XsEHaxkvpwQ3GvXyJ3UYsrWf+ESXDuGLIL5
ksh9G5Dtlv3N86+NcNIOqGSGvzZWy9rkxr+aHqngN+lCwxko5dsNV/R4v95R53lS
FrdIO29FBicYybiuCeH7tW09geienraozvTdBLkhYl5vbn8lLRbEhbCVSpI86n01
YphhpyqXQ/bjEqwdZK3qMw+N8ptSWL+fq/C5FFv0RNWFCXcggHLvNvz+9Id2n3aX
PtFb6vLNqgs5MDpq2gOhAjdAgjLVhF4YpgZTD3OJ/JlGtG09KKHdJtV2EqIpfHY1
GophIhSsD5yvkJVJRmquTKTzXgXcgw77MOSbzHPEkVRRGuKklSTqNvQeWCb2fEtI
gCF6NXnErTpspcG3azjMT9A6D74af/HSOXETWoE2I45OwitE0Bxc/x344cPy822W
nRXleO2hFoTXN1XDKDg8I/PHSAEfAbnXoRtCl2JsSTCvgU1kRoVEuD07C011YgPb
3u5o6/1SKZGr6bQiZSTJEX4SF250gJGzICMKvE9EUb389UtwNUnhvF5kA2O33WaI
XzdFAKPaNjJK1LOLJLA8nhWcHVq/XbGG3J/KNCrSXE+CRvkxdRx7sXQnpyHShMk/
vYgqUY69EXtgrpW9L/kKYpKbUc6ASZByhdDgm/NYCsOGJHrVVak9eHa/8Ha31Vzl
sVLVinn4MTPRxQWYoqvHYsdrjTsrXZ8r+eFL2DyNOo9psuflWB2VbZVANHe/oAgY
13CWLlH4+AlRce3cmAoQ9n8GstD3X+Wwve7ktL3hwKYuHyPcIa0MdXPuvmN/g2n5
sc6dzCfS74Vd/1gI40FyKBWE+E5KpklyVk7xaKZ67Qin1dedavv48XM16tGWrJ0e
xWyRjAtQX6fAG0hfYxHj0/oOU3e5lotgTrTuEYuA0UZxkpUjWR2P9NQY1by4oAJq
Ho4frJbraSl5YSgBj8TUJSAubgoRoJclTcqBAJ3BXqXlGDhbbdIBFKWhcXcCydIm
2HU31iF7neL47sWZSP9P5sMXCfgGuRtL5R7Jf32KXcmIJPWnozrk3AZwfMXtLr5S
/0FJDF70U6lZepmspEIm3NsU3BZ0K5l3Z/3St9sMuKwWkQmNNrB5G1fvgRRjCi6A
wJGdX0cC2Q+nXqid3r3lM7rxSheLRExsWJhckmohEBHaKoqf+RBPKTVLSlqT3OnD
HePDtalliGwyU/Sf6Ar4Kr13K2mpyk02xy7j+5kifM+X5m9q+YkKbhSl8X1qeQ5E
pAsxmgU+867zHu/+0/UKYxIIjnxEXMibuU23mE2jyqNoOmRIBYxgicG36L3Nzdy2
FKcZP2roo4FjtBui8yQ6OY4K5o8wgq+Ox4gSLDimcqRysOGfgC7CoYpZ7sK4cZ6B
IN4vOSrkza6GpIRH8X4NrThB8p3/qUgQBUXxzvFpsc9LxMqIYELcfaDFm7CpBbD+
xoXn8o945ejNaZs7spBsTqLAoGuBiy7lLCYkadrOl/j69t3Gof20VtdM5V7LMasE
4BsKADE/gbd+fjmeXExGe1dD40B/lAOD+dN4zjIkdyCPh0gxTOAOjiMy2lStGOhD
Nkzb6EcVRLphjoD2U0hevrU9BCon1yZytGiE0YdhJkAiGkD4e2zavtAtQezSQDqI
JosOR4PWyumIL45HliS+H6z1+xRVRFckuCM/pxO+Z4cpB1E4c31I/paQsp06VhsD
HPhDjMEO0JKzxnImy09me5Sgik9d9ybP/bpBSJ5f/Hm2brB4hg1sBhUI72/eUuHR
XMfe62T4KlA7GBJYCsJKv3ZyBDxH/aNUCpdSSZI5f8BRxTlcqrAdcJ59fiSpadJB
cU4blaYuNeSSNDzF+EFEwc6/SvjsPTVlUbrtgXXG0F3qcJjeDVfGPNLBI/xFlvAk
yfRh+bgifbS2aVPoZxUm6SdgIs+S0+EWu3hTZ9qDR47EV4EZFdptEflSn/g57r8q
hBi8vXt2SrjV+oJXj8UMbtX972qZoUdtUjejT8UVqaQtiogVHGWngHDSs9WIgbo6
v+ixj2tscka1vChFSTor5xzYqy1szFM1W/nLUPK545K9ywVJbYR/EM4dgylNRh76
oI8FXRZ/FRjpNPUxFqascARUcdJqBaJufx8IGl2R5AqJ/imY8ZOGKQAXP3OltAWu
GRxGtiQ95ZsBFGKAsemMJXx4/lrJryfLZBtQEWdyvFqBNaeNR9785Ffv5CvEXgzy
u0UI150x8i/ClK6guW0/wlckDoMxXBnRSpUIS87fbrFE5w1WQ9ebLwq87XNsvYpT
koGUK8WYq//pvH4A9UPfUauaGbCZDs0NPpnGhsS3/wNK5fpWtztJ+ojMgeSTBKio
spI6/z2CIXSZvPC7rZ6kGJeTjBILyLlIaR1Ed2Ox72ZP5TWnest9pUAYhO5CxS8y
Nb5JJCBhyk/UdhbEmdidaUbm+fT+Us8OrZzv+csT6cQbtEyUCF+bWrTgGwRZjpak
3nvaji7SPlYakKFTvPDkr1gvFp277PmGi1VwlrnxmNqnebeIBxjRqvIPc+ATjnSe
C8ZkYpdHeKrcv8RFauIM10KrhD0FYyonsdNhEO2IgkbZXh7RJlazHG2NRWLy5ycl
tcy3vcuXxH6w8LPrBIpRFxEyHfj+O3+n0SFTGPCeZHZOguXMFikAeRA9PRZS/+kG
9xsb/5C0XgFz4bW9APSATitD0F+u5fQVJZt9kLlTS1I6FJ0JiQQYoDDIA+fqTIn5
lUgfWs6iJqx05yZxiNkuiXIL0Z5Ga1uLccGMIRF26gzzaU7JDeqpGnawg5s+JBlc
Er7qiWVx/b+Ycmip0pg2zl864io+gwDyGSa4agGstiUwoJYIwllc6HKDAVa9aH6v
QGE/ndJyUo6qaQpi5eQDUFbiTSGc8wJpH66MY3uJZZIXohQeG3Rlzwca2g/wLqyq
1oPIQjJtk5SOfNWoEUjDyfW0MsITfeV7Vb+p15riq1Vr2N/TUVoN8fCQ5RFrkDvp
of887CTwkH3OcVscKa7dD+zpv3dPYLNtGaa04HKdDArh+gR1v8u03jjBT2+Dmceo
kZgH6swBiK3IwfN/YkV1hikd32e/bEXsws0Tt4IaNfbh1FV7omT4lhQ/aBwyk9vl
E9ZQKaYaLzDVr9RcRVnJE5HFhMPnYR8VHWIcOuyWdsntaXyOT4d5WO9ozhtqTY4F
sJEZxwNzfVqL0b1rvk5/lbQ9mth8x55kqWsdnjBqPQk5SNGn1xwNK4/V3CZRxlQU
H4VgM3PiAJPd5tBoweUlFDFtpQIYAooIxaeQhApUEZfNh6oatnBDhbkOQIX3hH8V
SSaU0rbGn5FQtc2Fg0WSBxXm15E0c0QRKt4fVry735GGCGrCfLZ1jlG4YWsS4sW7
zqS+rNKjqXZ/zubQJaBrBXUFsFA47R2dFq4lvYSzxg2SXEgJTQfXBRYy6dzf6x+4
pTRpvm6W8BGjomfHCN7ClIPIfCdiFuZ3KLJv3coNbmTTrDKDkM/ecr1LAgehn+wX
VofM+a8f47ISC/AV87DekyXJTUuI8B+7CdYsCBUn2q6lU4YEmM5TT0XPSQMaxRh3
/OyRSrdvUH2o7ejMU+xmXVZkMG64zUlf559ABncnnf6HRooYrDXAlSoyA4NdbtVB
LwYuka5DHa6KVCMD6hVdQdMp/JEw0mzyGcZF7mhuHM7GqR5VWRsg2xgDhqr0UGzv
KKYybel+Emn4KicUJIr4/Qza9dq89YfLgdh6XU7T9X3o5lV+jVOHsyr70mXZNacv
p+ZMrP5PJjDPbnCCMZ+K/3ovnlRN9Fc2qLMHqJypfhUwy9kJQtDTQU9cGTydX8Id
p135bT06IcgpnOqNOfDmkfqT1bN6qd0MmmHn9GgVXqJR3YWU9oSJyg0+d/ltQQ8S
t+H7TRr5TSj6aIN3mAg0rOaZD7/5AO0hoshWYYJFAdCa5B7eaLy/+F1inB43+dOg
Yqbsl/4cm5f5kzkVn9FzZ/Yt7bcmdYtHuGWrcyYBRt8fAAI4tHCbzGqBqSjEQL6B
E9Nor67dU7YoBp4qf0W3RNGZ6xUG9GDP5/WYlovBYuWKUAjAuyGAqZS0E0QSjfb1
RlFNy/u9L9fGjaKcLbNsMU8OWl7n2HMrzu9bbkMZxoadj3z1DHRsmqJ1fc8dlVIu
etDp7JwMs3PI3zFkRbmkdqypaXSps9x2900XTwSSC1lXrzbOTqsnvIFh5TmUxGSX
FGZotkONH1QHU5Oq1AS3JZn1baOI23OuO2yJ8oQWTZIvgPfxut7mPJEMh5XvUzMI
2dRuXvHp0YPP15moo5kJcC1jyjxNQLoRngR9dnvN6l1f50GdDXeSUAX5ZXF2Uh1i
d8InGt3KRBIyOncgqrRGJSEakN72Y5iw59Rnxw5FtmqZIcvr5ihh5LtFK6YZ5ZCu
/n+2FDpbWKA0nzaCfvpKxTOqnIqrYAQCYvuKXiGbopRCkXW5KvlY6kzuwsmxJoqE
+xbjjxoiCAim0GZLpCw0NtMcUUvmFeAWqyaEeXVP0QcRxpdIPvO2WEaI3BJ8jE1G
gdDjoRj9kfGbMUTWpAqjabbZ/hGSO/BXoPPn9mt1HHixoF7VCjRPQI76rjzhGXq3
msGGQvw9UDCOBKjBWWafzLkBDLG3pTKDXIfXTIG/xu+9XRd5+DCvSeKPsOqCBwVe
PJM1RrVA61PM/UBV/b9RSQkmarQX9060i24khFnUdRZleBxP+kH0qfkNzvboNtyN
bA3MW4m+9FiWyh82+Hbk1KPAWzc28Gh+srv/aCCvzT90d1pj9nQaHBhjcBKOFcBv
9T4DGIbuM0/W85nCRRAuN55k7p3D5ggqHboSwcy8h0lpW8Ljbh4qsB38LdEKMO2R
QLOiU6WgHkBHCP049OwsxmUtTkDovuE3eyEBhDNt4tLZaf3cauph0+ydZbu3b8dx
WQsUCZ7dLyOQfYGUSvosmXhnPAFxhqDeNFEw1JVzzlmGZqmCs9c29wgSL32kIX/H
n0ovwZwOXP/UQCuCZ47P4LhHbBbzOczbQSXd/VfqtNsr/SrXSgL3oCCSCj8D67II
oPhNZcKU4yAJX965M4bovCzcn5Ga/TO3YAa2z597jtQ5ond2/xObOKWEwsr3JGjy
OLLhapDUMuKg68DVEJOsR0HA9rrEUWiXNW+g93OjZQoru+Xir/EycAe4CfyQiT7M
Arqn15KjnTtNITgYHtyfUGIjogNCFr/yIjEF+av5F8EbFV1lO0mWfK/ma6d93R+0
R909gBVxfdl6fGsWhtWJgqywq0att+GaaR+XtPu3fx545aVol2Lm9ztY/9G6GQrE
uE2Yh7OgOR+1r2DhZcg68x9rCdTsD6+9/Y1gMx1RVoRSfqWgzPeDsgxke92aIMzg
+duCSUtviLnmYZ1XemxU6AwXLqnDznpMZhbPzu1axuHKBgojkE4ncqQzohdWJ+Zk
4PHBNg7Ime2fv9i5bA54XA5uWR6Jz6YYnHZVt3mqOQOgrcsWgzMi9Kc1PzFXu0gU
rNH7YjNQMBUlFlggazWzcZ3gUaSnCwwtwq1wZj1bwXKVfvlCB0RdZYnjagfRrKHj
rn25qJ3caEdBynP/OWqOFzbMGyw+Pxkvvz6UGZyLh66IVrAOlW4iOZiwx/y1AZvT
X7+zAQ9G93VL6tyr7baPFXLQvrFswrdjNjfjjcRM3BCCPLesOBZIpFLKmSS/DzsY
lzbXIP1gq+2o4T+cIWY2DXlPuM1AoQKfizuYZv9NLWaP1l+3ZC+BBLi0W5dR7bia
yXrYGl9qx87W0MQdgYD7rDwLdVLsRhmxx24TMQUZEntlO+oauTI9+wmccuIPhHtS
RPrVfx1eAO+ACry9kOwKsmhETqBfQnFjbIwUsnW3McYzHnICQEp4H2JFavRWpit4
v6VLew7NtKhdEDdwQN212i8mBPdtyIsgNfq7kGgVOj2Zi3ID0aHBOeHfqGGXA/IS
VzILz++kfT7NfTlGe/klPNo/stMW+V8rcYYMLAKGoz81qU4Q9zxzcVqOXPa5Ao90
+uwPwJKTfBw7F8koXO4V/zxaiNwbYhUDpbQbOw48uaNUvDmrnxyJji/aZRS4apsh
/VqZwQd+UOtYnOSCgTGtgivY1DWZMBYMkICYZXyH9JKkDG19K6Bv/gF4+Sray9Cu
fR4NrNPeg2tyzEhG7lBK99dZuQHuFpjsKv19U3ViDbRUhNlYFpzrpmPmjRp16LAS
j5p1nl+yr5xJ3j9fEF9fYnCKdNSMw5DPEKQoyavajpUacunkw9V580meF+75xxKy
LzHIAh5xAt6guSi4gyhAd6Te+JhQ/UBZhyNzppGjYSKhZLmBLzbBe3OxjzCKIQ3/
GZE6UFxCID+nuubL8FnUCLDMA1ICZkGbzBmg9menQI7jPKp7aFq93P8FK+ihgbKM
re0XCIAetaLE1cKuBVw4KIoQEHB+WunPtQombLI2KEUY4oTvaRxcoNHzBVdG42Fy
L8y0BrXFzKe60T+kl8t3XmBi2+4lrjX+nGUvTafeRUn8K82CfKaNVvWswdTiTtc6
kep6AjYxXfE+l8BV8Z0PVRKTmWa4Jinf63GMkWDQGBBv0UZS2rc45HIBUbem7G5k
Vgm5Y14BwEI/azzbCtWdM8AVZxOqWt67pRxqvufDpgN8tjRIKUZLP9C6A0uTaBWc
DQyK46o/icdzsIBbW23CSFspF9Bsi18HsyOVsSx1T1d2u6hlyh+bzTrtrAynbRrT
tyimhmA2PUwnYSw/EkO8mUja088zuN1cUmqqLy1VLlci6xhqkZXg/fv8krQQIWB4
ETOfgTOAO67/YbgztsP8tTdh3tiSJW+1M62cYyY/JQUWY8GPakMURhPIsS55hrA4
T/aZR0fsigjUaYoiyYRPg6RZnLVFTMtJ88KeT0muRFuSWNwlqQVBK3ZtVYkEhiB4
3rHSrtC33Z7TwrcSQbywLdtOqOEUwakclGHRsk+f7tK9K/uAQR/jT4YT/bQXnZys
trO0MiUmZ8kB8PyovMHY30mM9syqSQubT/gRQdl/TPql8GBzBO1awfKK6njH9e2x
FiC1KcNKMWSkDVKy4g9s/lTvDGqjLOQJX8jMwu7o4gd8r0pfuBgjaT2n7j8xpoyP
LI9n9MALHS3yMXKgD5qzkpXwNKfsw8ZcWBpMogjMMJmPnvksL9irJaVR52ObDlQE
YlZ6vh6FJ4IbjTM66fMRnZ6MpVqmBzl2yaNhMxbmc/zHT6jBzAwkbySUYJg/WObm
5ixxp1xRcAFd4c+oI0PRDEWsqGvZVQ5+HyVnYlx1FT0338jv+pbrIc2FNRyUXaaP
cMekgC+bEGBLnEEwm9S0A/uok5Wk9WzioUHkPSCYrXUkzmc69NjFmKfAPlut4qp8
dENG1058SbAB67iBTI1OIa1Ibm2GPaF7Xn029bnSYF9aySEZ8DJAQlVQtz80Lxos
EHC+vvgUWbWVKSPRXHG4n9QTs1fmsJYHGHlQn15kMd6cNe3o6uyurnc01fXGSSsY
Nj34ihnwztvukZ6CcrFO+NO4apNkg/spPlEdOt3tykGJvULJcOF8Q/wxuDFq6r2E
htldRMiZVCkWMJ41YVywM0IRYQ9k0Mx59xHjMaL6ib+PchJM0mDk1yj22Jbwlgpw
aWeY6msj2XVbtnJLCT0WR2gWJ/y2fa/uda55ur5xDzme65dW+sCp5biu3pq3Hb3T
YqMyncF260eZ4+aYOvclsYT1G9BrSG5R21l+8nF1PPsgKS2g5O6U40iEeviXluMz
2gpn63TmmjbWtVZq3F/VZ/O5fStbzI+kFOy0Y2cUQHhAiKd1Wio8PinwYGppmavv
JBB7izlKHdLw2W/WSLvb92rxK5apEhuB2+3A6U5rk0iEDZpJ9Y7EsRyCIJYzU7La
qBWmk+dMAil6rJRuqqZO6/+gdHat3IRiKpteHecyTqLay6QAcS69zkJ+Z0PV8gAK
LGlNDToE6FS9e1I2VNtwUuK5yiQ982Cj/uYtP3C0C4Ts9wP2iub9ZIH9A+MpTm1a
fIt4K/sgi9e8oJo8c3sB3FRjCagPLGUSYzNUUOwFjyvKNbGXNo0rOzeZ18qx/ww5
ueSbcwYrifv+9ykXBk2oFGGpS5gHoi6XWJNda9DHEhOoUbJ2m+qPy89GstCMejsd
vWtfkS5i4roCDS2k5vz63O7SiG1NI1ervAGEAAUUxAAHsWxLyVYZCKVuGQo92roO
cCnb3UX39k2n5ywNWB+zWluzHAmIOvjNfmVjwKq/EvSFgUROjxqC6NcqA5O/oFMH
mylShASH5D3I/NwR8iqX0pdgV91qplsydhumspEWlKsNFInfyzUG+AyjlScFu2pa
CNvtrs3oEeh7qEOoqGApVHFePTYW4NfmHIonTgUHoEVH142avbSNW412maUhcSEF
MdTpmrRe/r82KXceBL0CH0+/Z+4dC3ItsK7cfQHXa13ajERsXCOpavRqX6pMVM3J
tL7Nw4HYgIKgOlYUwvHPYubaDSYu48rRjGz+2qSRu5VrKJFowUvlTw9QFeww4wdJ
sI1VkuUrFaMNQjMBgPjBB41RiyP63JvP+0fiNYltxCIhz1Lj/6bkjX5EW85dQ1/I
/LuUGheE+ZwJTpM8zbkjvS5Y0K2YN0wzf3OhAXa8mwLcgn4IZ6xzimJBUV/4SS2o
Y4FsnJ35VSZ6drwoWcNO3HufdAWfeaou1eM+tHIaDlbtPyHjGseIARZR2izjgUnQ
4ulCUjQpMpepO6s9luhkfj8H2OI3HgEmx0AB/SVF4EpXsbyPUFc6K7FFxyphAhQf
3qXH+PHASkOe5NpKKwoALE10F7lspTlKTSE6isZh5vrz8q6p8fjO2/WaMZ5jeq1m
zFWIrN1xhkUcec/Dr44thvcJuhrSX0EUmza5/RjhlMnY0ZK2AL+tD1njJECv0jXB
Uya5Yp7aGvhRtX6o0ql2gKDqQc2qhCl++VbM9f3E6XEiMuXYnRG5Sg190FCvaWhh
LawvvB1SzG0uKCSHj8x959jBT7vwISBwHY5Hn33hgRLqx8Kn9LGiCdu1ihqqxS2g
phqaKPTyDR3bIsQ7kyur/Iuf6HaQydtvu5wsUgfffGntdatNRTuXbEc2aqDciEDU
1xt8Zzdmsv7YaliUXzNaFsC7O0qRg6HqfO28EMXgh1DAk0des9CzMXe1De8Eyl/d
3OZT5ge7bnMpx5g6P8J879ih/eI/7jHXLDJLHfpI+UCPZDhjhqj7Vmghj7NX0cK4
GfegMHJCBh61omwp8ANgJEDCpVPUb24eKynhCuZaUcGxzpyLOAosBOiBC7PVjfCy
ZMho1fVqlbE1zIslz9oTzjh6pgocUq2wF9Rpq7egS9EagmL3cJyJQ4ZQLDCoBFTS
wRqwGr7gNE4TOaX2btB7hdslOjO705uAu7kthr75CATDPk0Ak05tuhkz/GfuSZLo
+2LuKF9eB/o6ur7A3If6VxwwSD+MJ0wU9EQ7QsFjky2ebPk0STyUbHbWjtuPbg9v
ix10l6aPXC1nPn0+E7O9Ibwptono6lsqj+Sv8P8N0LOsqL2shVI522x/ygQKPgWz
8aDEa9lzk/Htu2sr26Vpmcm1aaZpZyIXZT691O8x3b//oJL3zGuyOg/o1Arhf/Ap
DdzBYxKagh4c2Uwn3qq8S7d5lK1uhLFFrURPHuBJnzQONiWPvvFTxsxbLKJq0ZNb
Sy7bhvRd/y2TzyPJj4Bw4aR4kvVm6feEFTTDR9xXlbd8sk7TlXZPDhV10dbGm91K
2dCIoT5k4BJ72e2+DeUnM9DzMFpZkDWCzS8TOMtfHGXj51ccuSMeAkky3jNkVxHd
7Aw1bzp3R8SRzae6S1HnYB6lfq++z1zBNgdXAFH/CfK2in6ZigZ82jVXdcBEJZpM
HgK6kwI7jqGFOna8bTIKb6/Anjb3+1pWAq3ZiJ1g1qtSPVP6XFM9C4iH0k7hEpoZ
TE2Mv8swvbceXzbRxdqjyGsPiy28RZ22C5yLNf1rNxCo+l7x8P+fufPmg9L3BD48
LLHSHMgEc+bkFFvhYtl025HIsCZdDag+FLY1v35t0iZpEMndW/rP3SIwzIEzMKMr
T40x52e/NssHFL2rSRRh71vSfpmhKev5zAznj4k1m02/bliUCl0m3mvTMji8nQ4f
N6gQ+3g35UD1udnfhSpfLUdOeacYs7fiYyzwZM2sR3tgEIgzCABJDhKrFFPA6rHW
eGgB9+tBXAQD2DXKzlyhf9tGlyidmzlJtM35BzquH3GydnQaV23jIq2t1GJi+OTu
nufZqUGbr80WHBhwDJJUANtcH7Z4yCi6eFrbCW9yz0MQ4QMf6C46XVRQ7JqIBSbT
cVy4LUzptfFZ1DjSQPA5Wr9CwqxpPktcGOahFTVqc/IOxUhEz4588mbmsg5/l9ne
o042Wi0c7RYDQ5aVpKJAwd2J1ZA6UFicxId+qpeNK1OLgIATkcDNlofWeDXfcpiN
53mZ+tGI4KUI/A2+bfi61p+qS9TfbfXVw8Hkwhuq0zWHQjfScQWvzwoUMgE0hdgS
k6W/G4KnrpFvUqOkIMwZzwT9GOTePU2LQvqM+1y9lOa61cRMFGebi/L6guSehpz8
js53Sy/7guKyYzBckwZRpcR+ePGVd2A9cJWdBzh7tMaZKR9RRN1XWn+r+kWWLMlh
8FOmaOLIPdzEVm09XWR4X8yIUz7XCd1wv/fiZhsnaPTB11VhWzAp7RNeTYFRnw8e
x1HhQShFH1tIOov/pMOQw5uMq3YyX4KsA33wb6bZ47KB54WkQDs6fOG2Ns6aAguN
j+qZhqc47IdfX+mcxWCF+R2pZh7Zt2ABs2lR8MLcX+ckNZ02TMG3rnf8a0hCAop0
Bpas9puUkxAdh0O6YqgT7mytmVq2JzYYtJM8f3tseNzK0ab5pP6xDCObrpFZFJ68
ou7l9SHNnFs0+IFls1xc5XKnJ9Y9Iu6n5fZiEVto9m0V3urxRECIbbEIBmMEZE2C
2CbjwJB8DQHTNr3NXZp0NCMP0BRRSm6M6i3yZM6SkXvZU38XJwAlWLpz8kSfZ+vD
F+U7pGJqwrSIAxEpQ0GPWMB4BDH7iwBGi71ABXFnk0j+Xx0UqcW/16K5XOgYnh0o
HCjoUnMIzoEgz6yaQ7d9EO8L9ngeKcJljAIqOaJAHMLcsDTB6OdVN/m1JotudLva
OdKiJwcoDc80w4upB4wjZtozqKh749CfflOFtcVP3gOljm5XFzKLc1ulusPCGkVf
EzvAA7Jx7ZxDjnqBYE+pWKUCsieLmaQuxhLYaaLyvmO9xzV6Wm2AlXMhEYIukNm5
d+pI+UnBX7q/u9bMUg0puCapZaM0eD6ugTir8kFep20QOiHglu7iPBQ8EDXRAjI7
V40CwjrVhYoaygZq76T3aNMWzgscyF34V2qSk3qaLHzwBoI0aXeS7z2B6UPRIwiA
iHcPhARGwpxDTNQKStTbxbht1JE3e2VDxmuRBB7Hk+tVnHrotLnas6w1En8Hoxwn
dw2Dsl/U5WPDqykGOjK7PLCcDqtfePOy9rtrQHyJclZ8JarOlMU+HiaUM37T0zk8
wZoceD4cvjggfiDQs3dRHNG1gBYS53hNSPpZElTTdI6om4QMOyuSteiEO1C4M4td
WESi6OOqRkCvONZOTTOvO8whKYW7hiYYbRzedDAVEdSyUn/oP0R+xI9gpRLG/4Yb
u9kY8CqCaIIMjI/newKpOl2QmimeU1ZN88B7UFY4c+WxnGRZilMry5Dc2v3zWrMh
jXYzB/lrg6T/Pf8/BkGIkaY4UQOrTesAxE5N6HY8P2qTlcy49EW4c43e2th07/+M
9GKsOUlqFhP0eNtmAwHjNKYLNS4PXcxXTzh7DD6NoNmLQFELF98KeNCrTXJoTicX
Y0TpDL1GUHm9ZJZ6ktx+yd4+ciH+8d21Hqu9P2E6lWb0dCC/HcIAZpIHFCYI0fWs
D+z+r5xHmKc+fjOnnbOSk1lHwEWw8u9SCz5HxGgbAKGc83O6eLSfHoqjMgjx1wQl
MEZzMCL2gahRkaYJIQ17AnZNLzjmSahbMBSvdNx7v0KYYfUY8VYzh23J1Fvt4AB0
6BQGr48lBD+VvgiLKuVSg1Ffh5vE+FJXMqdXAPMlOVStt/RwWOyAaFxG5UdO19Nb
5FFdR8jb3uixnVvpX1t1dCpHV2FDtpvQKZLaGPNY8Q50We/f15FXFx+wxAQd8Zcf
I0DcJUemtpvduWQB+N2xSzzST04xv/ssO/mYNxzSVuJcAPOjAI+VHs3orUaAVM5O
sFWI3u2XoqDS8IrppgBr9s11dVKqaIos/QkdFaVtVuK7PU/AUGeSkH53w9DQe/Vc
V6zYeBGebHcNCGkvXO3DfN0YKC8fLo7QPqj7hWtyJSO7OvI200t8Sj5TczXBCa4J
Lfbc/PQ3YcHUCrtm1d7D1+yAYBToMaMLg+2uvocRLccMvECALHRXkQKd0MLwpUoZ
VkdocWGP/GokmWA+nYwn+X17IrED8H70jTtcGQcFW6BENomD9xsMTK+wkq+hxMoE
pzxRzsEqEzNaNWLYcP7SsbUMzhiKL2eViNcXNHeDmXiLrP0qcbnVs03HUPawAczO
ANuBdglaN2Uj15+K7AWacwf3MzD/pWcsCl2g9CsPLhwX+Pq3W3Ep/2pYEstMgrD1
dqngMVGbDZnt7o3BurqMYFoUpnRK9UXRZ6SNm6EpHgnuUapkhHSgaLi2Meenr1en
8lNLmZvOyQHe6QpQVN3b1KJgUX2vaCAOdhUBR8CQPjcggRIPQSfIMO2J1Wj7xXsZ
Lf2E5dKPtJnkehlhzJk8URhBrUZ0UiEcMh9DcN4QQtOieQR8TFEVkAsFzFHJuCKM
lCWnc4Wxp5MX9ghO89xTkMg94BSbAKrSf63IUJ8dxmaNZAReBkZYyPO47iMeBMSS
+RQY0/tOJ3RuvZx9Oed37xFMX/0BeBv8FYgs27xMwdDdifluLUmGW/BUvRiQJYOq
uMp7H7iQSioI/zA/lX9hjnWF0Rx5ar1S3Dbkha+lYTYT64C7Osw3/6TGhceX5AaQ
DYjHZRykyqcTbgsfzt2Vj9udtYDyEkw7eTPj6D1YC8uL4e7u767H535ovuvqxvOc
pMJzQCs2+q6F0ZbHlq0PLuV+ukl4opMz+7AqCI8pGJCZv0QyAZh+mPO7DdBq+kjZ
XpVxOXuF7r8g3K36xE2C9VV+9AzR7N8Gqrt5pAlOBQTOKcywfkCfoZcDJRbHBWXk
8FZZLswHVH/llxqypnfftA0Bxq5lgp1x7HcL3VimTlF5c9NK3QH+XXcTLOuJ+YkW
gesCZyyMqvkuaqTmgf/JK0e0gOoc47GHaJ8kn5hJ8JHYOrTp5HBPakbh52/oXsWA
DYPDY1q06OZ/QlHK59+baU3NGdPxblgXgSYS9lrSlHWx0SEPxUxQecln3SgexB14
BvB2gFBK6dTldK/zh82DdHSHnDN/eJOSLtAioylzofVRRysvz1fPtFKUl2Jsto8/
kSwrVM8/U+j1ai6B9Lm/B/RCdspi3cGI487jmCVbjwdVf5Gn6tJ6nTN71nMfgXU5
0O6YPQEl5jGWkKVtk3ssbgUw1JI6X2cR4+xatb8j+dhWPEA/kudBy9W3rH56dPQ2
rS424dOxfnIQWvlqMHqNdfDSqQi12KKpYhX5t6ymmpPB+kUsiqqATQyjyrt4pmlj
UedG30h/Ddp6osZznK+qCHVgBCzKNIPnBSskPs4VPiKJ21uUpVJdF8jZgUXDuvKW
6AWSCJOYXQ7ZtDEo7sgY90fJ9QR4DQbRR8ZCII8h/VxTD4PCPentjhXfuCkPLn5D
BPgvEwgDTIHcPNyq4e8+UupS99b8n6hBSOYD1vYO41zOTdyFPIfomqbFV57N5D3E
bC5fOe+DbgCxy6thQphrx2LgUUN0Y3C5q3k3tkI4iWJ0cEC2dV8hQyYqpumI3Fd3
aBtCLB4q5Tdlv4siSSkX6gaWEhlyjAqBUpsCQ6U47sbRjv71tYEB0cTM0hmVREdC
T1LppKDMf6hzWkVWyVW9mmnCwUAMeplK9EY+0kgSGuQQEIIqyjlqxyFblCPd8V9p
OfAXtEXnrvVt5SDauTzlwAMvdVC8TTzhrNkQpos3CtnuKoPsY2bahSmamL+h8dek
URIP46ol+N8lCQjxCNUyVmEuVWmOTsNgDoDzHcfUWvvJ10CmSDIZSvNqn2Kx1b9r
mWrFxTc2aOi7esV/HtkP6FznxA9gQz+ApEiDfk52iIJBWeHcq0CAsGQ0vKgKiPhp
m0+fbZFcRb5vN6gpzS4AhHaDFyCSsvolt3axFm/W/p8qU0a8qCcC0Y59PE6dzgOy
RNBQCC4TC+ef7aHq+jpOTjEEx6SUhKuSNun9tULuxtk/xwS/5zsrSWeBPCSvIG4X
C2n+xnxFK1pxtxVT6iACGpJ7y8NDiKAAFQarWXaURNeoz8FYXb3hlPa4yv9VPLci
lR7TrDruFgFZ4fyWnFH+OU9v3J0y8HrHOPYfy1S5scu6z1JYKIGvjyUIEURUHoht
4NQyg2hAWQcZwtO8uPZGzKyrr+Eo557xn3gJp/yMYGW3OmaKOhn/QJ/9z/ZkFmXT
UozrOYLRLNJ582m/mzr+CE9pdXS9dHih48laIJsr9A5Fc8dKEoIjT0ux10y/QZyW
HMXvCSOlQ/0dZ6SgubbRqVySDvVv1ZeD06cASvJUtcqc4mef5fz0d3QUeQXyZoj3
kLkEwmd/AOKq16iPnX9EddjEroo8rQy5CgUn2LOpXxkweNEpKWhJ6MVMYNIEOCd3
aUSjoeF1JcNspBuwWxYBtzEkPSGNBxN0XB9UZRYnU0IqiOSkP2LBpTURraUwEB98
qNEQHI7+30x8EsscVRj79IEBrA5dDwiEUsBwOL9d9Q9cOQphiskZmh/MJRmT+0GQ
596suKrlYVdHOirHk7+Kk90mnbIlu9QhNd4Hc4BZkWBv7JwFDHdCKXHvWdiUh+ld
fW7bbapKa9hptDqKKqm62xvqi7MydZk/QRwoLQ+1MrEYLMkVgURvdsdVXNkmKfUl
ED5IPQvdE3aH+EX8XEpleYTF/fgNYiWlkxUh5CBSUj9gRLWfCk7svoG3fl3OY5j7
10B2ptCPveaJst02ReqkBjeYrhDerdZBZVcvpt9JX/DI0YEbgdWPcpyRTRTWQH3i
c4cmEjw7MqqwX9WZTJPiJdE5RAnvBxhTQO5YTPVlMLsSLd+11SgICGQYrMr1sP/Y
KttdzL9m1ilT9WnjBEtP8d2AlHf831Hr5KXJScifikWtRsNsrowlQWixmdTizyxC
98ybUL0cG7h89J+zSe5MMKk6hRfWJ3h7fJfnGA1gko2dZrxUaxXQSXr36KkpBUSA
Nkj2b/+ShvjFjNmasxQr2QdDwyX0cacUxTxt/VgIvRIWpe8BaIObpEgph596wLPS
iKEmZmuvQiJWBaAWmt/XMSUPvahoQCaVUrefLoFBm/h3i1403TNQNy/GhKtLFlhp
I9wmj5iQhLADcoIvumothSFMM1M/xR9d6h2sde6K1RgbN+RGGS1asa2tNecp9G/2
iPLy1MZA1IWJWUzbwi5zDcBgg5tLZBWiStsxoj6QYcREv3EI5aD7dBvnQtt1g5ho
yl5ltwW9y5q6P1VWzOgxMVvAp635h7E9INMdkdZqxLTJ77nGdSc3JODPMiJ/RvwP
mcG2WOlRIlHuULhNRiK4yNkdyPYeUHEkwYH6Nj7lMZeRXjTxQ3pwg1uSY43SSex6
aajf22P+pennqwGhPVdKQLIm4f42epjm830yP1ZT/v84cuR82vzBuOEe/bPaIu2n
nJ01GMal3gEAZUgl7x90rG+IA0zvPhayaaIkbcOHa03xgOuPSKlNG0OooDy53afl
CxeyAxVv5uUDuPrawcd56ObsP7dJZlKskEjJsbOt/LnFDNbqJDNWhLhYeIBoRFHs
/br7RQPbNuUR0XSbNBjV3Ok6O1DQSs2hx8qw4HOujQb4pxQmTAKyVnCIUYsHdlBE
2upK09gD3yqkaFjslx6pOieKlNux3QyQkSqnyPVCjFRXlGh/xx+/lLKOiJn44qiN
dP96XqOb+gqxm7RYrU9Byo988NmuuXl+mgivB4+Gr7hCNfOTfepGEijLhgh63NQX
EHM/QN0AHusmv1lJOpbUnZ7KlCGq+TmJsdfD7raHbItYsn1CxFU8yI/VRKZr+YFv
cWgvnme7dYFw0Of9gNFOf7dHrU9EVCcIOwibI3BS3CuExq3RDyFi+hvfPe0XefaC
XTHuYWYXDXVZNSnfj/rLnmpMwaSphA7Ydd5/kcThXB+9A31fwj86aGwUBnKPiwj0
i8NoW6d5Y6CCZP3Ofu+82tIwAcyiPXUZq7qQFs/daIej1sRsQxl9YciWHbCztklU
UDHl33HHI/Z3hKfOoP1n5bH3lWJs/pW5sT1JXvMmiqg+W1PUUN8W8uWEjgy0fTcg
v/cTmMjhbHAnB1h8J6M/GhyxacQrLM2FAK/SakzUZfnmNeW7LH6JrAQCD0CUb33a
0HXbsd5xTB4Nsf8ySBSUtOudcUbyLCDWlhm+NKd4kLvIcFQxSHBKp7e61tSH3LJC
iAUq2DcN1QSuHXwS1ksrY0l/N309MC4iURLsTFrEvvPRU9pcA9rBcQemzk5BKjIw
NigzL94AhuR2u1vGaEZR+Gy3nM9rOMT4M77OlYlHl8o8q+7qWTvfDJINK1PB8bX1
d3rRlZ0SG4psFckw9Iny1T3H+E1KIE+069a7lBeWv6DhiJvWjU74I3bSazpGz4HB
YawbS9+oJtMClNHFcNWYviKCYPFaITQAjRSfDCrbObGLKRVsE6XRGIM4EWykDohL
IpzJ6DX7gFskAawlwBT/ZsmbBqxCfIkiRoeaQ/juT+8pnBcPeB2p8o5gr7/TOvm1
id5C4ILftbFwt45PP9wH9uX6fjmCSuCiGXj9oOf+PLTQNNUTWanGf0uXvpbXT7h5
4bissshzUNp0abHOSGtKrbiWw8UUTuxKNwkywC4PnDb34vTRFdmo7LcSkJhBW3pc
Z83lkKn3TNT0h/PTfNGvnkrXtPaqHHcw8bnN5D4/X0vp2FlXmo9MbE6Brful533Y
0wR1/GCvKoHLFzjuquPks5BuxIVXwPhVDIC8vcOjwc9GzNVEvTJJO/8c7ULxhjGM
f6x95xuWMIfSstoN8DQq64XoC0X/ooBkdtnQEByqabVVvj75j3qTntsZvAvmva6V
YjXCw14PiW1QqbR/HT93G+VSXmFQfR2aSNgq0IzosnyfSaxaWb5I4C/djwx3Wikx
RiHc0dxpLFlNvcrt2D8RaZb9OPanS302V/rjO9f4sb8GFwnSiQL4lHCir1GQt2V2
mVVpVUM6FwfM0LFNG+pZMsgRx5SjgWjHyCp8CMoC7Keq9oiTMFeskq+cHP+t89ek
H45Kk6sXoZPnWUYpzN8Ku/hEKQuL7APo5STz/UcYQ5jkloC0iuVLLYt6CLvMFNgF
GQuOdhwjljq0EqQuTYCV2HqU//vsGC7tkeNnWhL19lF3i5nQ7+SeaSX/KCirC5/4
GL+Jw9CG+8tCg/06Itnf2zhiGWAV/zoUA1M4dUhRyOVUE5Vdt336BvcDJpg55xec
lwZ4HTcPnEIQJq+eEnVjr9/gNv9P5TNv6qJFK0veCA9QZM+Het2ZFKKJUgzklj0F
ATSzz+AO2O7Ag1jNzDaVtAaj4wUsT5XvyLQcc7NnPu7NBWLVh8RN+lVw2ZiNrnnm
zMWLAPnPKpyURvqL1mmVSc6ebR1iGY5nCVHBdahAQojFUzcVJWfbWu3cp/S5O/L1
FDqIbK6Yvzp5xGoyBBi8zHm2IGQ1KLqqKFQbNRIFRV8ADSrwEwJEwyx/upAc8MIL
MK1saR1H1clqUh7z1VbMv7LHs3rJaw1TnMtnR436svj5NTc28TSXQqxdTfnWLOac
T2wTbhPGszNxDifEta9oZA1Fb9XRbhTIAOJfgqSVfVremNBMvBA0YhvSF06E4d+S
PR57APfuiIsSNkmfDEyV0CKWConQXeOQMaHZrPTDmp3GcetSn7Ql8SsXky8x7cbp
2Nf/UScz6S5AYWgK3rS2qJWoTYOtGyj98PLexZrpl+WmZKig9x9HpCWAN1S2t5lM
nqusj/H+2ipiaSv/oXtBRi6FNpKBsAIqxkwu+cLOuR8+7P30ed9AMz2Lzr2T/F7r
W0r7eTerlq1LgZJAaF+FSFZWMyBQxlRKrkqQGH9knUS4+TsyDdugYXNzUylq/xrJ
CbsWlLtIwP3RuO3DAA9iSXLn5Ng/JOUUMAeh/g3KnxGI8KTblifjm9xK0eclNAje
cGcV8cXIo/GN/jKgH73dyu3R1oDksRwC8w7fIrTXrWfybFPu+n+CPNNMcKV2qewy
lXlcn73yY27Q6ms40fGUe5AqpFAxeGUvKujKjkLYBK0cjUZmjlsyOsCiudOnQukJ
zF7txKip1yWKFewo3TTrwgbYTO42diwUfVybKhIsgGxD5hHZMGIDe1UQYAXA1bNP
Jzw2v+wk6k00+LK0SlF46ZqVaaY0oB/XAOzm5ApGjuIs5YSR/S8at3N1ghu0HIxx
hBxp8a1IubsGgC1eOEkw0mSzAgrYk9ZL3iWhB/5lXPX8QoHbsu/wjKK6NlbVqiAI
QC9Ny9esB7TBwELUyeXs0aEvXbraiYCJ+OZF4WHU++2RTTdnIf5Vv20LcXeifH5i
/x3rCFDzLIIkG2b4XCkjGdFR7VNzdeRh8VsuqMUCNsoTZvqepg1yS1sXZDIsRjjR
julEoErrLdfOmF8Q3wfG60tIpaV1LZJ5wP06h9LDh7iS1sqvte0k0Nx0Hncq+LPK
U4PKVSiJjvRBrJruGJpTgAumUXUyrRZITXh6/hINddchdujVtfVwZt0mNHIMrm6o
7FBKk6EDBMz3pKE9QeVbdKya5+KV9C4Cy2BCMj/qECdavIQsclFRTHBWQu3pJ3j7
cHNgbyUkmH3nFrG2huqvph2jaRbujgrLnR3Q8MGvPpIU/HUjuoKdYiY2Dmz8dHEO
q9iolNzPw+tlDcRibpr8zfRl6LK8KdINW2ULHi0u+1ii13mlghbhJsIaNgQZHW5B
dm4cGPOARJppMv9MogVAqeynG5tJTDHvJSc1H2ufGMaxELQphhDbul6asO7vtEk2
hDOdhKZX0kZSq6mpO0jAeY7CwN0VQ+NUNg/xgD1Mo+8v0eWs/lbiCEOxGzxxj7vS
JcE9mqegPb3DRUCfbUqKN0cXFuIVccQ8hvXqPxeTAmktbV51H0ZgHswZQ1NqZ4K/
7lLh/X9sGy6C7AZhmkGTMAM3qqF/TRs32CZENlv2qWfXHm991z5UiY7/gLrsSsHC
IjLU6uLMyJsfkF7EfYsZfKY4EQpYVj7l4Kuxw/vzPi17Y8hqr3RC/FJGyXKVJ4/n
qXf+kHEaHfgYvPI/KnMqvlG0uxzSEoL1eSJ2daTDnTiOX+PnjliInRx8g2gVwJsF
GPsk1li4O/qrTMHM56nDgbqxOgEVA2EmwTg3IqghRiCwaG8cgdP+Ez90K28ivKkr
4GPv1DUXlFxH39XiV8LHk1rAk9SivsWNaAub/nEKaQSQ4xvK14saStv2L/5WIDI6
oqYR1eeGZ+swluPgHe5MzwT4JfeLxQjA8qeVmzS4qSNHEMUTwgSR/doete/ZXUUR
2rnDAnCcnqhFYsCb7bdeXyYPJ4owt5FrukIt0HoqEqWkEkUDgOBfLY+VrcmiYGMw
xnfqB+WCyLDSgDHbirDjV/GrMgy+wTR/bsUuc+zyvl8zPw0Gg/KeptCv7bxIvgBi
j09Tz9QEfLBoV2GLvJFn+k4+5vaa9Rv80C2wT8B07z3f34UTI6PO6KbQr2Li/SyX
DEAjlQXEcKTe8/nRjPToBpXuce62LZ0Q7uQN3RLyeG5J8HM4gqM13T32FN1zLNDp
iTT5tuPlMYyioIaV+atxgsnOXlY+/1hNxPkpIWgWU+PT2XOZjMzZKatSLK74EReZ
up9pRabYgJUVFbKUWhu0pVeC3cKWTDoC3posBWpNDu+Gc+cQzZP6iU+67H7cnWzS
Iuq5xecsC34pTMwSNYQPe4YSP8D4mrh/hSF26R8Gwh2HI9+J96vOjim3l8JDwVLw
r+WvPWZ1hQFInlI/jHC5A7Iy2SLDl+Tvr9YXeAnP7G0yTt6pTjs7m18m4Z+D4oY4
Iey1YXMyq9Bdgvo6qWtv3idVI3e9sssz807lXR5Ssnjivo+ztmjpehb7omJQU71T
7QQQVlZPhDwtDYXNv9oX5Tk1eqyoIIQeuko5Q5h0nyizVHvZu7ArG0nZ8HSb+jXz
cVq8vgWozhNBtV3iYz+sOFNx0NUu04Zk9HHyg8c4IKdwNILzSOaetAU+hq9/+Aov
BXlY9BYlVlJBZtN7aowqjibjr7iMe59pGmU9OKoG7xuAQvNr/jN1roBNdszINpf6
WiRG90pGrIXBPyjs/+Q0BqqzNm7rJdPDb3zt2RTII2oT1dJHAthz5hzqlLLb9TmS
HeaE6L7qSs466/3xp+7n9cLI124yauuDU+baZmMntDjEmHSG204zQ5Oo1KZrdYdr
jC41b2wu7e+7rzcLqDyGpsU0RRHPukUUldJM+e5ELH20XXVe/Xm3Nm1e70bTMCZ3
fDQPhiXBgct3NCWGQzYi9vBEhBhDRzUqQkvT4s7/rv7P+X8bvS16Gf/fFvqfpLU+
hgveCrN2ZzOzRKtZqcW4kcFgUBF0pqkYSBeK+kRlGpBhAtpgnHqIqCuF27CvGcVF
aQMZ+BPh4AKERe8AulETBmtUJf9XqWiOSdxoU4N1HFJ/LjZePTcPGyUroaIgO/Zz
qPgwzt8EZLYfmjKthvedgGwF1oi4WYY2zCwhtSuLNnFyuaKJGUElX3lmMPe7G6To
l5oQJ5pgVmO6pBkuu0a0MjRYD5An+chhtLBbOSOFbzEONoUHMR6qQ8aah0MW2rnI
OssfaPnjN9Xy3zQeLPqY37324nIfqDF3JqvVUHpU67Z3D5ZgpJKlQGlRcOjWq5zs
SCMmYJYRbiLsXh1tbUkE5wzHw9ExIbxtLyDpaFv2qGJUn+fzI89muOAtYG5Oro99
sK9NMuGeOK2nuTINVWWOASVoyDdEsNTRghviuOyxLaQmD+guq91hBz9AQAVmA8VZ
1NYsFW/XhesrODSJawgJr8DOtR6VEne01so4IiCjyMwYAgT6mS1WgaY217wasak4
bnaiyLAhQwK3hgCOtiqCV/MdP7t8I1tTgfon8v2znGaXoHbswVzpBULrZs5q26JE
J9rFiqK0loQFGbIycbK2BN2cRvIMp9BluF4dUrMERk0Zg/OgUV43ogm4w/kbVMaX
bydytOk//xEx+Re0uzeTdE6RhYhxLdUQ5fkkCp05Vu97MbzVCziZdUJ5OX21K1Nj
LS/PXYgix6ZCj2DgR9qwg6Kk+nqmPesi7d7OyG7raFWj3OFAkstRMORaj/+gjxy0
2NTiKFjLGDnVs1dxlJzXGPeMg4g98vHEpiCvp6S5Zf4jC8w1CcDGwvXGWELve1w4
Bmk/+wpPFIwTDV5uMPfUs3X/nRRathQEtgFYeZYlfU3EpYQs1JgTsVtaNHxUetZY
bDsAjSJIUrScrDfrfqk1Lw+ldj8XSuzqk100XyxzPhsNp6cD7hqcSLDzVOj+cIaj
UZ3lwGaWjYhZJ4q5OV2K/V2zq08iIGgabX/dLE9Rvy7yRpOUoQVPqDNorlpruyb8
VEdqJDRssyyanOiWrvLe3f/PDfLSoN96EEhpk9Ygk/rcPVUgqIjKxTYyXoB7Z3tG
+IKi0J7+sG328sFJsReZVDMcR5B1+pqjT9op7yMp4l0AvQJAQgqM9FOaBqr48LKJ
h6nfvcgDUtGNyaxPSmgWaYxIQhVyMRSph9/hTvSW37xyq1UF5rMyFQ9EM8uhWpto
3pz4EButAp/w3uakNJ0dqdWWZ5AADRfwFrMbEplTClyxT03al+melcZku/yrt1Gk
0lLfD9s/h3TZbbhVuKqKFO7li8YXRkjXjydo5l2mk8sMDxQ59cK+UiTqB2Mut/wn
XHxpmHh0BC+UYKeeF3DDTfuvFtV0KmBq8A0/tQUDF0iUf84actWhpJAqb7+vkf5Q
Jv5DopTQMQG4lSDMYgBk56v63xc9no+ThrduBkVOutJdcvHRHx8Qo8C+CoG7JXq3
mbmcfZVta8wPyWQa36gM4hixNEOPOWA8UD6nbmtWDH7d4GGei00oRXlMFRTdNIn0
pNk0A//V8bmPMEa6IYOigyI5JKE+zkuibhdS2Mc4nrVvstJAZUEg2qp99txPNQbS
mYU+3BoTuA4hCj+xNR5CYy4J5IRgQ2FA47bwy8dx9LLeBTOJmy+nIyeyHo+2dLnW
ojodvgLJ1krG/mJaBH0sPxiLeVJ+ftBV22LAEpYeWyFFfgREhXxJpAp1baKZl1/1
Rbf0iXduLtFbottNPxz4s3bZ5+4dvsfpl+7L5iZxi8GJH2TyoN6r8Nqc5Z7Eb8/5
6oL65hqbsEriPgYlJbOHrf07C1M+yYOj3a0K7PgqjUW0ha7ecwouS1mKLWz1i5Og
Ruq8NH39NQzPMyvQK9c0ERZ7yomHSpefw+6ewQgSUEnw6z9XHTnHK8id1mFyKuRn
x211CcYZL18rmg1uIcpx+tzwoTvEg18AEgnJvuoKGCT1iE0ZEukEoiluUrLMvPI9
MWtxQ44t1eJb/6ZMANEe17/Ui+BJ7jv5/SKsKto9SCZeEYveLg59ueVIQ92P080i
MumBBtso1MURa1ounUDMzzNNbHeYmx2e7rUHDovJ23WtbJ/koVYEPMSaiHgq69Rm
UiEso+W0ABaUnPjhbYUavggdLx63ZR4/MmOzaqzkrV7ZsgwRPc/SbBsCBLF1OOAP
hYHGnnykqJ+fM6eIo6825mDQG2NHW9BNUwFa5HqbenG6X2Zb0zg5haeVpNY0lTZW
8jYyW+cLmDoYhop0hUAJ7YpQdZAzAT4PPMCM6n8umBjwk7+mb8cJ2fFX/zXqEu1t
qtJj36bCCLgjzfbss9Rr42OlBy/ybakjCZ7YCX1v1rvPY+71ZEugLOVHiwv11AGE
tmdfMv1rm/u2HKlJ9ytOR/c72Ba/KLrm3Kt0qwNkaf/X7mB4/SP/QfUX3uNfc2Bt
8SLUH0lWEeAlujQZUzxn5C3fQbB6lPKdESiTD1jP6pSNMPtZWLe7G5CyMU7zrc3W
8Jv+M2lQYhUvoE33hcHe7JA4IErsIsSgorF9yvd3132fqvygjEae/lFqjKJNVf7K
qJvAsOUtYNa1SBgiVeyIIM9VRLp1zlg81pqrvjMdxJVpVNK9EbYBDkR2eJcttAzu
JZ6AkvcHb4x8dUxNFFRJdaXhFEhmYEMdF3WVX1t/f/xRx1R0n8ssOweV4K4uiJ+V
WAzDKCLPNhmjcAY8IpWLvjvGFKzgEMX9k41qMHDpA7K4XL1HKkC2F72fxa8Yycwa
61QE/hBz9wDt9q0JCZhpPegBAeve/Yo6O6ecdDP0bO8uQzaJcnyAwUaVHRUwhsPL
48CpVSkIJSaWUociAilHFlyHJtLkMjmpFShxIj+H5Oom6bK6uxRG9U3BDiri9HKi
EAhbhyjb/36r5aLNqzbrKb4zIqGqvSfgw0RWQ7rD7cZXAPEpqfXHxghorQPd83ch
EctI3rXSk4Icd/Sq1bjJUlx6W9eDYwObUZplWt2IN4TylZQZ//UyGrRr9SCW14fY
3E/pMKtcjuRqmpEK1dLiEVMhXkj3D7xw9i60paJmUm6ruY8ZiOmvXIswmSIDSndD
ivWkckiDScGS/eethoUg9ZEtxdN4berkrzfrAmCV8iYUlDjn5eUmiXIHcfJWmcEg
DgDXpCMXPK5m1UQfn/OEmeLjaedanITzhOem6Mq1sczByQtDDjJbiRoy0dPbRnWu
Wmo0uO3Ik0H9w3TvKJPa7lpg58DQ+99zTX0i4y05mLXg4TRascKhVoimq5/262nb
WySLkxK9mowOrV+6USGsGP/gTqYZAX4/EZ3Nxnp2xmmR47bwx0gqlpJWE/khI2H7
lfBHoN2l2XVDkfM3ZoKSHL2EacfI5MCpwXEiVUPB1JYaheHXDWimJI6dOWH5ik+E
ybfLJ4x8UyCxQjlXqQ55Mh38gXH90yagg0+WkCt2XUYvSFgwciNGv5FDbDwm35Tq
SIle5irWFv/9mnlrSFYNMATmypW8dTlq2h5C75iHF8Ykq8l1ed+Nw9IZrDchJQ42
tZC2tCDiGx6UaM3OtUYueTjTFEJ4jqiRTKCaLPfM3z+8R7a2QIyv22qcUHD22LbH
ygzEQNv7wtopOaLVExkEAnAyonFoLS4mwoAJsvEZDFX10IhlisnaRLWYT1PQwObt
0LuNp7CRFy+uA+OKYq2+c81SUE/j3UxTz2PSNRHkA2q7yrCjePaa4YESi+VyLHC8
WE665wOvxK2AH70l2CMq9ejvifGHVgHx3+/jyZVFzUrX4HNw0OsxlfYirNUrj9Q1
6T10NvA2f9Vmi+WxnnO/JtrCK48i25Uy1xTybmssUDvqtpZI4kDeU6h4efnBWEXd
ThHXYDebqwBQ/PuqJ1zmxXwTG/ApphkqpF6Zfo9oMA6m/DjLpkyiSLdif+tC62ld
pIY3bcCir4FxxoSkItYu7dT7mYHUgweEqaaXgUn7t8vRLu8sK9J5RauVRRGzTClm
dSwCm8RL5sx96YiDzeXPlsDCxmgPAuriCRaHMjUqGPpK1orI4w3bKPmaLZFoHc4S
DyTcd/1N9W5wiEIFTjOhaf/A6UR8RVcRhLHVOUY6fg+Wh8NA2fw1YAx/Pq0+iGAF
NRvgkDiQJ8j/bNXHZygaejYsDiJWXDHbIijkW12ho5ol3LQYu5nHrXvg/GKA29hT
RAWPvIZQ16nhRlKRk6fFcmVe5TGklfbwnag4ukU2ujAdODNOF1lkNenhMurS4pc0
EsDUbMXOUOZeR9Ke/HVDuZXzMNFgOUORXpM9KNtOBg8lLHe0Ph5ZLWOw7V0RKD/S
OtNt3VOdgTZKI9lKQIao1UY2n5s2xXjCS0vyK369zWaJ4EWAMqVF2ZltKq0vVS8d
FEPQH4vACMkhN+tPXzyiboLv6kD0XEOQpgbmaNtruQoAb0bsK7JknC6VW/gI2mTn
UdbPXEy0asUjHwUIBCL2s1TO5TTFpXxMSBeUgBfhlo9dtZxitYlgudbvCHGgmNsv
e1pt1TJ6g4Hn66QGlXQXyGTcCLQMM6EtM0UFGL7MFu/rpT4unUSQWWqSmV80UXv4
NBWPk4kAiDyx7lOL8yRR9vyUcNuIjpRsNZrnViNkVNTPMqoaX6CDEvRr6P3/86HK
gSZgkzNYjwCeIfqo9aW8oUKalOh0PwtJIu+a8SndyAAtKDKm/EEMjYV34pOC6Wit
Zn3Z5N8kAWmTKE5JiMgo6cEyc3OoCqk8GN1tLPgisqiKYLrO7FhJuBbRNK8nlOny
BqZmtaUCFtEQw1s4RSZ5fm5fC2O74J6Ki5ZeZR+69+qEf7/QndvijduBKVLKZjUX
/LBQTo1Ig2gctImbA066kyTSm1Wsqtw6GCTQLF3ulrH3BzvfarLeARkjw1IqdwU/
shIbd4UfDda55v4F+rXTHgGEwz2eBX3drr9IaIkWlN9YNuQlGpv10p1kRdrFFisw
Q25Ikvg1J9RRsisem0jF16L9dNwUf3cbbOcVXibLzlnFUNugfc/4DX8rJ/RIvi7b
OzGJZDNnTxj+xyiDCIaDnNWtXbei/FoyalPykKUPyvSb1PG+ehOky9fRv8rHZgDA
tVP1EAo9Eewx71MZa1b8Bak4P7ZmUZK4t/ykKPI2TlEXK0GzUn2yp7IpLHBnh3J0
2Ork4jSOGG/YhNObzDR5hGVGg0NPKPIm31+KR7p/96G+jsqn0+VPW3f8q2qgvM7G
k1s9uylOzith3p/7wsT5c8N/hASPft98NcLkxJNrBFOGOk6iK/X9vpRRPs8AeUKx
oyscx9p8U4CgtAh4YsnKc5bHWm0ynN8Dx0Y+/Zvw3RJ/dxS4bQ6O57cQ4/O18Pl/
4pvMMeiWBIpHlHLU+/Vi0PNekX6AjEvuEvVFFZlmQQ5WKSOgO0exEpcJMcU9D0pc
GR76VZ/Mc5SF1FKMAgFWhgkUAU/dnDgtKgMvDJeBJtKP0LkJzQmN6yAw0GDgzjj9
w8Q1HXuFYD0+uZNNvNAjT4Dxas8X/oZ8IB2RIzVrxkxACg801Wr1HdWp8Hu+Af27
6BH6S42EsRjFrn/UgIwJZIfNHY3WhS5ZolDzDanCqVoo60RyNYC+wZtKnwEfcvSQ
x61sUUwJWDT0hPbLHvKPN/1jRMjU+aYJSFjSmia0IL6UfU+vaPD97IytxsziubeR
bC8S9Om1xnIvcfJooypMk5ah7kA7Bh8Dtk6U4DQ1bNuXAkcK85reXwlJwyKJrYP/
erPAKLrHY3xJsGIU4mLRFlDnQzd7M6cdej7eRXL0ws6+oc31NN5mnYqg1E4dLO7p
iUjSNjz3V3XGO+lz8TpeUrO+rb4EDj1Gm2PLrHD5aZJBMXv7pMyz0HO/yWNJaChh
9+/uGDJXq+SjZD095fKbRty7m4DH5rqOSL14wawRftYDnGgyP9wbsm2MPbnwO5+E
6CKVRxqokNH311MEBD2UbmlrHIs/zi+u1keg9Js7zO6jCbyTq+UrRKvqjh8Gxlv5
5exJEwinCJfFDr6yu3ASoyqCsI8c600N5m0lLmnXPAl9lKAU45ANhMq5ftbZK5sB
8tIxmUh+TAs1rzN32C5giY5nj3uxFJPlfn7j+xr1hHWNthKkXCeoeJW/jgoBxuNJ
SQMlD9qTuvrdPhuD0qmebNO+TOxJ+ggSdcE6LbSCeelr7vUsv9TjlLEOOYsrOUK0
sDH1vkJdR+64aIkIAY3jEtZezRNoIh8eaLVmT9koHJNao2jemGApXGDwxbIe4Cif
X/tF8tfUcaDM2zeoMXWQe8HMTvOViVR6XmhAii7R21xngR5DMG79sEjr7jKSNbic
4zO7cNFd7i5Mowu+ZG3KmZNTaA1YGHKJDJ6HWmXJnvkUVv8IlYRcKKMNn1mPVJdC
tQS4kyoRAgwGjQyFBDBnkzfZTsQhI+o0NYjpcUANgr4qqieSBHJiA2RfegW57Akd
N5O0wHxlS6VcYBCrPDVfHW4qjg7fxDA03knz7kOUqHr7ESjLetxDaUXd4rtAdLax
djP+Mqc5kqIPW7ACuCc5xRkOOepEUIesPEQtUIFREOktTXt3O2lWSdozgNk+DziY
jDVuMC0h042GeCZ5Jr2DE6uSk+Lhgazk3qmyV3wDEQKOd64r9L1o2ZxOHMDRGEDw
uaQ6PyvVunN50zpNySqegp1UZSUXSCsdK9b1vC4vF403Hgivu12vhw+P6WzH0LtM
3ELnsli8GxPr/Z1nSuuVhUqdwEo5AldZkjCubN0fpG1X/u6fd5qKCiy50HGVA7Ms
qRg0O/Ht8I5sK2MWxntiFBUDPo/tpPhdjJf8wHsL11Zq3vQxoM4uYmBDPF+Jhygw
yhfNX3pCOwh1zOzdRESaCSktAiazrMRRBz72s/65ZImXwEpGtdZbh7l1a8nvUYg1
lD3VdjqRYOe6it2WMHM8WfOLVyvF6mFtjQZKZ1SxyguESat9j/HMNd2r9J20V77P
XgIYWmM+wpTa//oOMiyaclTwAoFPqwOlV5lFF6ZZtuiVBRwpvVwk9BEt/KH/fxPw
F5MAYiomOEiK62YvSKp4HpRsn5iNDeZUFZB7zvg4NqOAo4eC3anTguixR9ADgE8Y
DuEBGl6SS+QDZojDMyO6+cfTpbiz15p/CWtxiwsu1fuBwfNOKNhr37D+gcNmY/5e
CRk0b6n0bBFWF93tUHEv/siWvOLbvyPaRCIvjE+abAB0z2s/1QH/NZ8MDBAjaRTx
i/k9r/b45AzZc3JLju2dFUe6Cw8crr8f3MZuMF1J76rIziDiqq2fOw2wQg74gTMD
B356WFw+HxpnCzOTkFHgtFJQ+QQAywHGOZbYUSTuXz1knvrnP++OOApk/Sd2e9ha
Yu2gVkzVJ1MZdV1dL4C6nVMpaatm1AW82feNUWC7dNfJ8szYnktPddFqsOFo1jja
C0hQFPNZN3ZFc+79nZunfE9Qu/bDWOivlqTGQej8LjiR81L6L0tXFrnuf+L3ftoC
wYL+P6uiJ+/3vPGgwIBBZtUEn/1fCpnTN9KqBExGvsxnOWJ8RvEkLFBc2+dl2pgT
NssgVWtIkRjLBjkbTwMSF0ydbb/gVNC2k9ne3c8VuqyaEREomxfIH1aO7AmusyJb
ypMSnPChObjCWKfpmXCPThd0iDqke9EFRWJn6/QRIDAPx/TvcC1w9h9eZCZP8BvL
WEC+IVhQEqQSO1FzztD8sBSxEei1ssiwXFpEwq/oR3jtT85CHdxev6FLG4uST7Vt
zuv+fCIZfa7knrJ5YV+dZ3EVwYWSQ844E1S9UhqyE2zQfPz3V23ue51jpziMLe3s
Zl4f2DD9Me1eM6WkGtSPGpnPAIc/UxMHmKel/CB6pERRl5tZezZh8+UquXhfjNCo
zXQEyvOG1+wlan5tR7f8LI12MNITK+TZgt1sqNLUcJeLyEXmTCWX/Pl+e8TofmuP
fBtSL7VVYRY2+kPeTVV659B89reWtl8k2wb7pP71Y+gr/MgAEtoZAeTwSLtRCIOr
a+OsqSxWTVALkBr4wpmJEY3KeQTxDjP8QasElc4r5+PBWZX9/Dj8+o8oG1czPWkm
mFPMTw7o36VU2rs66xSXLBQgDIm+ZnDlmhDHd/KcK32wXpNCl2xKnlCOy40nN5av
K6/1vlytnzYBup29Iuf1gjAu01JzOUYdtzP/ed45ppExOgwmKELiNmL1HpIgeW6m
fk1AhYsQTJJ9aM4M58xJB5De1dFovEMWGBn8TEb2THW6L79VbMdDkTwPOgZwpEjs
GROezHWUELE1wDY6GD7IDIbd7fQe+B8EQ+a8/3FHwRdjJGUJBhM8JNjlzlI/rDWj
+wGCfVSQcc21sdgx6/7nRJgvzX6nh3XpgIfuIcvhpMDqai9ImQoHvjyVLCluoY67
J4gRLf+Ij+ffBOBHBHaGuo/GwUNbyRnAbirWjazEBMtU2ZUjwBi/F/VB2aKE9RB2
jn//88jyfncpVpkQaGGT+w2IzNKD/oKFX3FltrMlPfY67zv52R1xZbTkXmChAZoX
bBwKyiF1I1s7cwTIeVD3dqyNfYssjYXLSD4SDEtrs7zqknHmXKjqWbn6exbL63Eh
ltX4tDHlAos6hE4ZzEIFu+hxSHx3B1qppN5zvlbWZa8FulviayVo/oI8oEDICd1q
Op+smOOuoR4PfducU6bzBQ2uPjvbvTTKcWJ/KNjw8STiY3EUtb7N1vl0/nf5LhHp
Vsr7qkx4Tf0Go9vxbyg17BX5klCx+RgTflNYvyfVZ7yUeCKMAw4WpNzPGaP/rG12
2yYZIJa0WPRlC2sdkVSy7LQEdgordT7WG9spgDGtGRxofuC5xnzK/Tl+O7YHCpV6
B7/wY3yWwStHi3S+oyLRaKQmOBYg7hBBFjhrG5f5AvZ5717w+J3okBn1QTDvBleo
0hMHSkwguw+RJyn8EXZhp6SXGdpWvurDVG+uIoxf/PL6bOzqhXJiumKVbybyu2hm
ahY9YYEq3gUyIaOKHOXDh5V6ukX2Xk10TyMxbxjBdOmqUMnoyFXjtVRp74JvtBZ7
gh7kL3dDAsGCxnWlr0QK2tjauOCh0N/al9FmOgTGMEZq7Qx4jmNTaoqWEsdhvWrE
cuj2DpHiqeZCgaTDzeLeJqHOpi/MXbtsCIVqhBNQGajdn81pjkPX6+7Cg4MgNIYM
jSrFBNhaH1EoxGXMEeLSD0PEIdx8/u8QBW0YY+gXb4/ZwH+jQWgBDGkn5cP7hoF3
iw5OFioJ3ze7W33IYSljjv0mn243aoV+qqOSRI8R0b12iqEfO547s28fjLRtFblu
txxX5DmRdSEJmMXxet2i2fMeOf7jgPXRi/xYpRmROeizv+MPL6zT+quxQuoOlu3w
sojFpnejTRJf1T02kF5n5ZF6fBZUhghSekbBUthJVXBCQCSeBmyF1aQkOIekwKVf
pYWED1zfrv9nPbgCdcmYJulG3/hNfs7vzX9da+5kPMKKS8gfee64O1LIDvik751K
6xDw/axHWdjWQ+9pq6cxroQ3tnsmYBbEKtZjwZHREQA+p7eqo8kjXn6qPG3v4c3A
6dqWpQhBJK5lgfCGmYvW++g/oR26XSI+WYY56avekRc69mMPF21zAoGxjxPAxvp0
OjpLb9GyV+iOokTsijBGjefsNZedtZ90Jbj3DmlBRGE1l3A2e3wYSqpW64fEOpRB
D2PhUkVV4iezUBy6kBpEHy1xg8RHgDTarDGfokLo00DyLR79dtNVPvZtmijI1Nel
vk9D8lXt17Ou0mxTGZNARpne2w0IIsn7HG6379E/S3UEr4cVBxmNfEEz8aqkHy4/
XjnvOylegok41oH15AGX8jzSWcDTBhE9ykg8RRU/+YCcR1GKqbfGahwMsBJK3/1/
jl/Zhqgnu4yWaS4UonfcyN6K+y5jxX1tMEUVZ0ltw1/szWjxKToo50HzXzZftTE+
EYGWSfQIuxbDpRHC7G4dm6HkJyjvQysjRzsMaSytp0/hGAhcO5UyEvDp/D/dz7t0
kfBDYd1MjeNOsgszScuYA8Ug8LezmW2I9fK/l1znl4DCf+f+4SzthyMs8KJH1cYG
R6Tp2xPx60AZ+f7FW0VrZfDpjuXnySfuviVG6XgH+D7ph85swM1x442e8dOtjYx+
wxM23MGg8a6VrnLKadNu0CXD7NP1jsh6sUNgL1TLBpr6AE6A9Fa5WyfLjr954y3k
Wby90K6S99Y/JUpL0YMUGIs5CmvZf0t/c2qgACU9jTV5dcNx2+6GI899AA0BdYHb
UIUZXnPhpIV0CIIVpYGqoKyswcW4RaLrCYGopMjeTnma02fknn7Q84IoqpFsSt83
3McdFRvW1MLJb1sxJp4nbCxu+y27a6x/O1Ekp5HO9j5G5hLmgoBTVE7g+QS/v0QE
zAX5AUqiGeIUkrcSVLMw44RWozWj0Oa8AMWFl9h6gsR/3rdY1IIwNQM5Xh/EGujN
pGLqNzmixygNJgnbWCACGy/O90cbq25OtchKB2aGA/qZmyjcSHRK6Rf203xFp6z9
8QmOs5KmI5xhqRd1I1OKDVaNEDeGfNMnyQpK9KFbI7fl3HqpkzMARl+Kv9oh2vec
toKcrAkgc3qNIX0N96aTcwvrsJWLRhO6lrv+Rm9f1sO/aKD2uRTK6kBVwPUh/CDf
cHvb+mrdXi9hkxLvrDAyRQ5dr6CZCZG4KPawOyCn5h7nQW6ujy0K8S1miRFu+kJU
9Sri8KBT+5FdRxFbE+egXkMVHwmEZ2XQeKIy6MVnZDpepGjqSz9UREMJIwXzBQwW
4vYUzqj7ZLvu2fgsnHd0B54o/KHKCy06d3ahdKlVfJFPbv3Pe1hcH6Pw1trUeT3/
s3WmSSyuFwySrqaKZH/TjyNlvZCdTLm2V0BwksKdUslID3hYzS6CaT5QXWhRyDz/
WYkUpirIPz18OxEDLxs1s96YEDBvMMVOu7ofD1lfNEXN5GMkMb4IkBLvXxmWDVgj
y92ceFTp9Zcrn5NpdaoAUKum4PAZCemcH2n+6iT88H/2akovcJiFmDgXEV6Ya7qN
rxEhIs1a4JwSkFEGKAJNanzVazGrApgIkYl+kzQbtkrpkltHgmELJfwH2f99Wx2L
UuNkhyU0idJBe6RFSSGOSRXw/Puomlk6xZt5m5ZLHnq954KahnWmEeaXU5ytc2Ch
1zIaon64LOoKc7Rc+dzNBdgS7WoF+L1O4IKj+wJlS0EVuOdXkuiWHGE8+8GOPBIi
WCBhWhXxvdy47k60CaI1B7LRzUBLxKKuNzZM81U6AxIqWaBZ+9FZUkyLJPTFhdrG
6u/TWPzqSXRSfK3WIkeM9pp3jhv+Vq9Wd7dO1WUeT6t0CXEPE1cC7b/UQiTQ6p+Y
9NiI9boDc1fq8KkChSvyrOig8JL8ohawLbKW4ctqOqz85dfbNutHx2qvzi3oqD0Z
Y81GsO+iI7MHE8OgbbE9LzKS6qUmFdNLbRENkS0bJO73EAV31+DVXVid/dccRcgl
E1YpkMlQ85afRfkCUfmsJfiCDySSyslieYone4Efu3834xUJ5BtUfMphnAilqDzw
hzzAns61nk6ZZtjwklkgLbJoeAnHax5eRH/17mDJiYm1qdZp8SLjG0n3SvIphUha
ljIAci79p55Rrh15jvNTlgFhzukhpyYyzpxz7sp+L4JBWpLFnKsdMrLmTZwF5olk
fIVN82roEA7HON7qJMuvKeLyS5D9r8ZFnj95w44CH5fbbbKn+aVPIP5NBmOY9QKg
vfPs1AAcOIa6PJCp2xcjSWApwVYcCSifFqo/pF1DCIx6rmTfoGQsao/dhSTFie44
VZQp2HE0IVgH40TROaUEt+/sJ15GYyqOqbMbD2Lj4iruQ6h9YdAjeZJBjq02YnIR
TwR7jPm2Ck/IONV6o6BbWfySlSxTmeoFgmeFggdsUxd4Ippjvg1U7tms+30X95RE
sU/vtu7066H3K0voHEbV5I2kOqVZT5SdPGcw+0ZkT0IJZa31NbTvt2e+2WL2Nu0L
As7Vzw8r33SAcEWtXfzO41ga3MPU1SqjFo794VAzjDzzGSugZQopv7g5A5z+2yFX
ABv8AnZA+m6/8EfULfpCsVNB4wXysxZUtlUhoZBKIxOm/iSJ2boMCIkp3tGQPLkA
wDzy9x5MCFitf4A0ng4FNbZc81orNzF1YxLXKpvghdWu4Ecd4A9SmkFnJNRFxS+U
zMUqeG7EmD0gKkMqY1xe3QOGJOlQYyY4FHzvcPyrlQnmCCvlswnWJaYKjmiRRdOI
9tj/jDyKGgNg53OdpQbQkwh/6CN6QBVXAyDev0Q5gr8hhRffaaPUUXIxw8lbTJG9
+6gMbYLSRckERSjy20TTGJrdC+FtEXv55+U9nggG2gYj++q3LdSi/iE74SXHwWOy
o6Po9m+6BJZLZPDxvRWiSsBIgIiFmccoOuegRX2KKGEhyAIKPdX9P5IQ64VFYhFw
r8ZrZFoJ8gKZu7pnxvtN/7riP7rFN7g+GTSKbkkbtlfTjynjUCnK3O7Mx0fS5dlB
QY6N1xXanQ9AkZORNBllBareziMyQul/P///ZGxycX+OpV4VkJ41sBh47yG8LIab
jRI2Jlj3mBh294S5gq49uGCd0fSOmAlhf2tC0eLcc26W9EE2tvDZXcdFBksJQSur
MwyOI7wD5g0CnHVB7fSoQa5dxEnI2XdFFr+M5bUiNZNUg0BLEPHLvAZ4ZP+R7ba5
gyz5ujFjudm7rNoD3Uf1iCbq9TNp5VlGdN/kqphkn0RJOpkEwSf8Cfe7heN2eTJa
M5aWhFlMLv/w3nQ7i/DtfrnCoV92Ag5a1JLKX4V40MozI3KExgUXXfByTu+P+ZPM
/od85oyA++pLmADFHLX4WSk2Si2v6dXAlI9aeaTjyBhfFgjW5l3bkkE6bmJbB61c
WV3EOwh2a8pcQlel9yrXAOMrcDqaoxK6S1wrAHCvN2qhwXYRuqCib0xsGq1yNwdu
BFZUeV2uPr42Y7kNaa3VXs+Lm22vTYp0aYI9HrusYUZkqctVTPZCIPMDLrbqWBoJ
sitBxBRZzSM1uw4mm8v/zQ2qRQ1JcukPi5e9MzlEDbt7dtu7V4Ag1LwisUvXv4GU
nwjLpvPZ1tmVoysgSqF1AE/9nPAN+Ra/UdiGX3LJ8Zk0yLiCahsWNju2W3kFLzLr
nzrPwebqbVyTU7qJpwiMs9D44/UPM8rY4kb550QEWvNFIATFW+druXS1sOddtTIe
nHOSS5+udmtKn6eXnwcDKOvgo+y5MxpzoHX1XYqghygj7NATX5GUeuQDFK16Wx9s
rTu0ZXoupHSnvXTek4+Y3Au3LPN+Okdwkouhcz4zHUAF0mvw+EatvWTyBQzksMMh
RJplzEyqOUT56p1ExF3Cz1KJmhhDG0LruupIJtZxZyGIIO4ierFfc7c5HZfAkjnL
+L31tJKrTsdFggofaNu/xEBpL2Tui2asQt1nGACNytklSwI4sKPwh5TRLtnqhYW3
n5xpj6uA2d8iwi/apK50ktd5zz2Ufsht1obEXO82g1tmtmgG1wkSuTfa3Yio+ypr
wVXcE7WnI1gVvgoo0ZZKuk4PnAs7v5x1OqQ6AzypFA4Unoat5L5LcTIB4nuV2Z0e
OtTjkJeUzfOEU4gqhYdtEvyeszVi9PMlde2tAdtXdZAJ4Sy1R3L7XZ3Slc7x7cV0
IGmmq/EgqcNu8Xrt1ijWvl4wqJKE/MebMuqTh6cBLsD6rwdQ1BNoM0w3Rp5szH0d
WGmYo/yAgkxFrOrUpRU0tKtN71hMcguUMzAThlc7non2t/ayP2W9RlCwWmAPYazj
5PUzl02iIqcG8PW/j6pJNZXfeoqMtqkkSvOISm0PsZFeoQRqjoD9/X2HeoxHaqLj
jhoNufG2Ot7BBgifmRL9wB9mCOJ17gIDpOhQs9UpOX5rc3W/Va1t1aePgeSoWzTE
Mm3R15twmuXvma1y+D4Ds0x74tEap03Xz6AfojsYA65DN1YDWRlz6RoIEuxqGCGk
Syv76TH7Do5amT4uchOceSDqQibt0g3oGRFqPtRksjmb3ZknOlDT6LdC4dogc5Pn
909KXT9GYWGVbpSA9Td6fmachzUBILo8aQsL4pW/pDkOjFwTt9Vmv5z3KIxfE3Ic
1ffbxK+EfoE2r5Eaqy6qnuC5WoRpKIXOx3z7X5sZ+k2Zy6zLu/n8mfhXMMIHmsXF
aaXh6m9ciTTvCdBU0QtcIJcX5wFeEiWLqczqHLEcQYmm09blOzF0H9VzXf00ZPZP
Eze+z7+Q35e5qjb26U5jOBHLTzpj/jIy4UOCY6dvq9Pv2Fga8jOrFGP5nMsIhSRD
D7jCYxJ3W8TIhE6HIMxLC5R26ySnKPvhurtVwWN/nXF+o3j7Xthfic8Z4lzp9DZ6
3Sl500ULw8xqv4R7Wo8hWQil2SL5CnEpFeDfiP0FKraoqynerhfHM4vhWs39eCrA
qyY2aEhLTNeAm2952VNZWImsgQIN9q21TwPka6KmFMCqs79HbhtGT7rwZ9HZ6/tx
cYH7Jvw+/qdvWjA0upH0T956H7BhJaVzKMiyhdZ2b2dZXmh0XXtr3hc1ldQBr5yk
9Xv5rINU0acrRZX/Xwt/6BkvAzdxabkS4nO9qCY6LeBWLDmAnj/FpzO3SkU3docJ
PcH7Dx+T1imyjIcPETRrRlY8OqhXLV7PpckQJpd3RipF4fzfK3nDthEE0E/aGPVS
e1A7rpe+h5Sf6FfQ6P+X6QyuQVoKYt/IARTsrafEc+a7yA1+lVp4aci8I7cN7i+q
EgJHeCB+Kl8aMyBQwDgpfLwqwCbMQjey4BeyDSxk0hTTmvoyRGpn8HM+jcDTAZLN
HzA5iMojaDatOz7J/tWvmjn5zrTIG2javc20QrEQHZOE0l9EvCLAaeVadm62B/NG
jlIpbqv2BMX5whdynJiCBFclPgreXxghW7xU2mPFxlxY2C2eVV7MwcOKCFJxG1Iq
CoewKyC/XrcWxcvkUwHp5jvKfBWE86DvKzx4yakFXlGksueHJH3cy0pe+jpyB0CE
VIIyjweglkwMXa1S+jr3ajXkjwa4cqCEqUxr3/apualGG3AfN6l69Bic/PNshna4
85Lh7yv58kPCt9D2skUSW2rbHLicOOYTrQ7/K5uDSznZuSky6U1q0TVIFRvq3L7y
GmIaaHQpK0MF+PzsfHJCdlIwxeyaiBxHj0fffypXsldErgtboqMir6M34Frm0vwV
fn8mIGnTdqNVyErIIRUEcS2wub0uTQzkoEXJzXJJPgBmmxtsnScvW90h6df59CL4
zVGq84ZmeDdT+9P7+F6707Em0lKQv+OlUM+4lvTTknYjnZ0lToxaHi3oRxNGug2l
FG1HJXBhjo39EKYl9MpswrRnbIzHMdNXHfSayTAuS2YY6lb1gmMVYIe3m9f7lhiO
o+mbGzT0YYNW5jz+HZaCSIs3tG9S2DF7rkt90VdqLZEGwpOCUIxs/gUdv0dlbe8O
3OpQoF8V8EdWB6Iqpj9TJd8TaSba5JIPhXs3Lei2VQJXl+sGCLVB2Cc8q9b4E5vO
7WjWtQSja58lPyPCe4aaSrPK2wcSF8QDncNt27PbBVqSJeG4vc+XH4mRy3VhNj0g
+AAEaxfw71PlMHz10UYTPCP93zrxa7FCXYE8CuxPiHPi1jeFIxqCYPVcniBzAH5o
BBAVmE6KLEdPZvqBvHdXV4Mr+8LtdPhxQNIvUP0aBjYocund/j6tOSdsirmqzVUI
o7EL9sfpLR7P7VFqYitPEYiELLJ4ei3PVFFOuU01ugSw0z7Cd87UiJFLAOmRvWCt
wxhrYWTUqGITRZqmkZTLAvW5tRZ//vprtT9VLBbaKcMs2lQqeQ87NW1q9HPPwwYI
CBkAc4WKBm2XVMkG6YqNNjjiOsWmmQPFXRXMvW6QQyVUqpQJcYxIpQWpedPwEtTb
GXXGE0VKCvsVSqW7XzCoKUo/UjlpI1yQao/GNy4TdoD138k3/UEPYPZPGZYP2vIf
+ro891FC1rX0meugmesnNydIBv3KxeBHP2L+M3EjJbMY4759tqkhA22+InvjVGWN
vR6DuZLf6cs5OiBY8ecT6KTCYPsPWF2pKL3KrLbezk42Ba2OerMU85d0HGOPCmdO
xiwwWqsQ2gQnOizTb6HAiKv+5Z5wUMGQFud2n6qiAbud83cBNBpwofDwHpkl/UlA
bTop9bXRwptkYVUI87fnZhcQujkNvcEWxq8HwogP9rHwZspsBK0jMC52Bgff/izk
STGNqfhebuA7P0QMDlpR+Ub85F9p03CocNxTMe/1VRgFingHqSZZYXdKZ8rMyvbn
BkYWljsuYVITAOUCqHzDRgL4W8osHCrdU8V0mjOsyUerqzBvS51XhXo28zwTIuD2
AgoV8/TEITcywQgcJ5+4mWb3iYWRU2b9fJ8xPQ4eNxn4UOUVipY1cfGazf2CkklF
lC5TlnKLKNIQ2dpNKkFGRtQY6dj/Ex4S/Z7iJPdenzq2hIquzSDR08wyaFUs5YYZ
W9fTkJUmxCZhbglCNIBHQMlkJuZ7ufFAZBNGwIuBP3Z1pdJ1cTOt1sK1VFiA8/Tv
2LNIq0RSWEuCW3J+g9y51Smn0CMODhnwah7m4L3G8txUfl2ZwvMFYf4Qy2KHd7VO
IeMfsSXxPEF5P69G3+jApVHPfqbwxfPhMLMi2umhVo1KBlfWMFpOkkEhl01MnFtM
ubQRfYLhpgTmqJzsrFvCTbriOoKUWB1HkA0JDzGaTDmSFIed22aPlN0oFIDXltD7
B/A74SNLJUmh/TOXR3rggg4I/Eh9BGClU1OQ9sm41LptBwvACNHEvX4GsWfny6cl
0Zl2cKX9J6C4bMlNM9sh6U+NvyU0lKCdcNQO6ZtzBzHIwsksUyyDf7X8d1yj5uAX
SBCKISfC0CsMVPihFkbhCuPgxH+475LVYrVroFJfBi09Yd41x3NTEBPbxaIidDaf
hFFtBp9nluoRJxUPE8l8xHbM3nS9iU8yRD3Y+4+027tPI9gFbFO+CLpnbeS50I1G
ZdLHeez7XJ65Ij0oalgYjyRu4Cr9Bvi4sIxPxWDYpzY1rcachdyogUMsUD6kWfku
sizDh5czPczc73moRZuhgSgh6v744sVo1bnxnLubZLUQNntiE+rBlTYn6L3k/LOa
LOf3aQtBiByHnaZXm1mCnz/7KPLQELIOgiPYlUAkvEUDNAhR10sMwJK0hY1Gpcxd
/uxMyjc1819e+XSy24Hrujjbj18X0qAb5zBtjTDZQunkV7JbgdvFUu8OVbZlTTkh
YVPshN00PqgQkL95giPlrWDHdMaftibHpTjE5yQxBbe+EGJKfTpLOpWpqx7OSJ2y
fEB6N/9ZMrCwgrYGiO0DW6elcu3QvegS8OEm/ZSscfnjIVCEHuKzy7NOL+h38Yzh
0gsSxMLSca0n6AiW1rfsh0zD7wQfI+0XGzxfHYKaLNh5vHtgxLErJyHc8SOZLoef
re9HT7bx9egFqV9OqcWwhjWDrlsaADHnpOdVOq5tu85Qto0Ux9jAgAFpKqGSgRtn
m/ox4xtVv4HpI3WM+Awol4zhK2V8O6nHSj4A1qqyTgzjdVZplsTDJWMBi+LYiu33
xVve8OZUcVYD4XmyaMwenCmEa3+c3FCkGBxivzetyr9JP1bg1cyiumyBpbZEPMTD
mkDf+A6HWGSnCD1nnZs1rrHapdBMaHAvvPKoUHCzk4XS8fBL7sYZ2jDJ4By/5VXY
rKjwyT6tuRAc4NPiau40gzGK8cZM18LGTOwYvEWPiM9nhakhGt43auhRipRIzq2B
Kt+XjRf35nehz2ayh5GcBZE6HOxTPCgkLWZnOtEueZqSlcKg2xnp+hRNvRRJx3za
NPCYhbK5O3Ve3smkxvWFkobNJd4h4ceOfFheCcD17kG3ktmHV9492JLmHc9NohNP
OMYad4WQOGIEguiO3sWEym4pyjj5auygq098y6MMWmPIiMA77PM0/6avzrkUOI96
upcte0uqqtMNw5XAtMWJjf44/wv9EDnLPQPs5sCTWG0Dosn7M5gqYx3bpkE4CG17
Wcv9MPB3fXGhLm/3XkgH7nW0z6/r04PPq0A2hFOmeiXz8ol6dEw6KUmXkNYc/n+T
Sjc3IBfXP3y7qfy49t7kG7esrkSMZVz98cq6PR4EkCzJuLqbZgLAvvKX+CeGoBlZ
QbYluVO35kHoBHVeTHPzrdFlH6lzDx3OvyvzNU4J/ISNRHOm8djY/iHlUi+/BbXB
ecvuMmXUaOLo3m2WSXh6iVXqSCPBVlvZw3s0sGWCwmXv8/HO5Su6ICL2DQSzAhvl
BDwki+/aukzNRmq5GZejEI6v/HcAiKhIKk1X25uerAyiZZfgHPWc3yhkO6VSF3t+
5IYKFG7krBQ9U5E2bAJ5SYDlfnQ99neg0vhMEdkMFEMIn98i8J9G/sR+k5HRNjBm
IyzvvIO+OQspPsFo5DTiCNNo5f3YmEDLOsI/Vzl/EwC+LvGduce+0hG8v2Mt0qjw
oyEWmbrjEXnimDTl7Ce4Kacq74IIL15bQugG0is4WOBnJibI1ADCjy/XZFpvms0G
35+UrZFYxTMznJsHibUqfIRMUngb4qMqXsud9HyDzU0bXotzSVcPqe5fSUZoE6MF
Lxx+He+dmijpjqRBjGM1fnVmui8JqiQg9zb5svZFtzGuSoq+hmJhf34cPP9NnjLY
7KMiECWJPDgAcDl2BPs/xBJ2MsV5uG0wYStPWCIcuioP05ybySi94cDfOXd7Xmru
L+8UOuJWwniSvwMs044pL2Ny0TyogJsMrgGnUmqOg3WI6J9SA6y/ROgFajprCbFC
iTHMEJPXpCdCQWdEYsvcf9svIJz2ZSBQ9kSxsakgJlWCi4Un85kV1fIQIaKHcpWc
nDDq7YywOHaXVQBtbIB4JUW/RcTnsJgXlnkq1E58W6DwPQxuBw6jr/N+DM0khnNI
pf/LwklG/bM7e43KwNMdVz6sypt6dkCCTRz6qPbQNAcAfPW22MtE/ksdWB+P6K1+
TAKbhbGp4reG+rNGlzQvGwT8+/E9xLnyPrrWVCwmUpNIZJmqZrzMrfpl6IV5AaQS
Ky2++EzMWektCrEjFjHFABKTaN1Xjan/ln9rCFSvO03sW9YEh1igusmi8CVzP9E7
DJjQu2TpszDZpbEnc4/3KqXkNXHlY/Uzh7gCjzWkWgij5b6TZw2vEjYs/y8les7g
ATvJBdARGKFWz9DoyzPI/w1zRvGrOnisUT1E+MIVGvAb/q0xQqxVOPUdP927sdlu
jqL+hLC/0uqt3ZvwXqM/98SYNVxlbMGk3egzsNGdRbIdTUBmKxFuMq8Hx7FzOsVs
5OrHNFCvsUc9cKKNSJyTjvLTiWogxue6yroN1lczlW/bs0coIPWdqNIr17Pe2uut
29Ccyc38JJz45aiA/VtH3oczFNKKA4seOwX0oXJNEy1iqHDA7oKW4AX9s3FdBhYy
wjp1/2VQ6az6fqHrqvFaboa6HCE2J+99zQo835310nB57qGF0nZF28p3Tge0rIgK
O+Xv1pgUe8tuq0UP9aoWOLwTH1clLNJ7jsIofB5/g6Ej+VdXaEShUkLvZ3rjgbvJ
2drQufIJHPsHCf+RaFy1XI93cT9gLUBQVHcEuBjsaqYkolcWwqAxNpNHOM1DW5f4
FrECdZoGYGzEhjvUEtkAIhaQki6izZwR1bQ26JH1u8pFt7g3xvK/m4uue3mwY9gm
HIn3Fph3/eSlCNLZYZ6/0/FJFdU0h+zIvbpfOw/BfECFx2yy+h5f+/w+3kKTwG9O
bl8styjGU9Zt02G3hChxYF7vlhsdcy9KgUG7MzAQZOPK1qAF2+QX1SBxxKdZ/qmO
XW8PvrUgfsazscZ9ZEZXysqun5SK7UY9ro5vTeC7CXxWniTFJy3zSkQoYf+MlFX7
kYprRXNvX8fJkKshz5oQaIV5PDP4SqEa313i3S8i9eXC6RXjS59YA9QaeA5zR8+v
cTBqt9Ygzisb9ipPKcxF+7W6YKAI+JuQcRiVQjocLm2fIfe5cytxOWH8WzmoyHAZ
bCjKWF/wML0OOP+6eCDvW7VQ1gtCCRymcOVdAkqQqjIsQCZX5YYWIgOqAfDBMCe5
TMYUM2KjvLPKGbqKpfgqtyQ1M/GMJENwbYqj++FTktbafFRUUXkN9uDjSqWpYo5j
L8dZWVGhmMUgZaPnuZKlkZdTxnAilK9Zbhb0pfQeOqdWAUFKGjmDh99Y08s9h3K9
x3uAVmHSKvEhSt0FenVdnbNlWBPJuVnmt0JBuvebqWTdW3xGRkWWCmDl1JdP1LDZ
lqWQ8uiX3dy5z/fsMbJs+5F4inKzZn9fVmJ8VMAEkf109fNuq6dPUuNZijJwA+ZB
DgD8/Y6iF5YYkuPUZXETPETpAsMVjRpTLxu/ZNmkTTqCQ2gArVrUebe+hethX8V0
7MKOyoTRwmM+1EifeSRWViSSjHvExzkHHm9vV/ddl8LwutCQYTLfNYFZeQkOyNCT
Y0hyLjdnMTpz7QrZ/7nBGTmDgT5KPjc2DYB9vRa0h6jPf3tmrHWZ9EzBzGvyMhIK
Fr7kZ7XaUYNBJqjolMmgdkmE51QPH+NJVDMDENbF/tAb2RjLSGjlNQckgFJabxLS
Xz+97VTtIVjNjgOZF9CPUTB1dnwDi78rY0MpOLcrcn4unEh9uZKV8SysPwj2NqPX
GbPGxkfeY2CfRDS7y9M01hJSD0wTPG40PCr9ZIunPJ25GFRP4cTFnhMcZMDjNxA0
cUtZZdcG1Bvom2IgRLnDKzCDnt0A6sH0W/uhQ4xhhODpI1lVr8GMUy3/MoJqF9JV
28djaK9W7QGnuqrPOIqi7slqN0Kc3PJs8ulGA8XjeUAVH6FW9xrBxYGFC2U9+zGG
5q8fGVxnFvm4Kiq+dUj91O3Uyzm+kwCm4T9U0kjsw5+Ey6gnKpPq0JduLXFqXdxh
fOeDgw/7BMICJVf/fq15HorSTBa4CUoiak6bEnveCzveD0TqrcDGyUek/8YeBhVD
x+8ncYyh6pHt89bjRezCbm6LdiEBnbpjbNGvF5eCepUYlvIW4F7p8KqAPqC4hM6Y
hTcyFrpBK3xn/MLCdFatl5z2HX9cpPK413FQvZ6qaTYPstDzHFBJU3/HUrO08mGI
FQk+fs5OZS0ZNsKpzAkYxpUMIYe4bt5QuVinX60oyvdm/QZjEHyqQIkT2vYNUVc2
LRA2lGveHEmvVEQiBxjyUj6rDrd3k/qYBAusJSt4ZtOStV1oXXy6JGVkp3vIoqH7
wUiajbEbtcqSBSQMz5Ij3kS4JXi/bMe5VYuPqfhGJAW/nhYS9XO9PXagg+rZhFpF
zhcpikwlSrac0V2vaX5ntaA/UckOIGR6K+zMuNxtuwRnyk93MyimHe1KhQ3WgtnP
6YkXfI5gdL5y5OoTftiLpd9Yyj1K7UMaSC7t0phIQu04ESmoGS1HUbR+MN0fUxvg
4n0/aXqPNnGPj7DeSJtdo5Mu0BVXpvbXSYbkWKI0stVryxcewReT8m0tj0b2uSfO
kEN2+WT/INGseNtDvVU2O+vstWJ5fkKg7DHkSfqXOsQsbHBvk/iWBKDBI6pF67lx
1uUelEI34wb9Js8kv422GvYz7ZgIO5pMKRMHsbBoW9Z74LlM4HNu9vuXQ1cRM+u+
ZHloA0yYu8+i19YT29YljAj0roU2G9/94pJulB1vJ7Of2lmiiEzIjTBtqak8+puq
17xG/v4juihrl2sax2VIH/vkQ8oltQAkvQNuFV2sl3Pn5vA70byWhCq9rVsZEYc2
PI/hc7kNLcz1YtnFzQAmwhhpJ/K/7xWFTGb9x2ZD4J5+IiHW3dtpLhUKrRnwrW1B
Q4/ZV0iHvZcyp+HJiuUDMTOCLhSEIiKSmX8piiJsJYBW2sSY43RhGcgLP/Ch/WP7
149W+rMocz2z4XFlsBDIo5fB5glJmsHP1OcPoZ7Ygbb9fWHAJ4OoI0aMQODA51YG
sPXHambLqfAPkM8zYYeV/9VbjI5Z9gnX6Rz3LlcqDqyBDHOaLCWbWFHTuv+yltP2
/9t6HTADaR2jR/KCcYT0rwyD4j6FFMOdVB/x+lPdbIf7TSRgd3DOJFsOA9zz7dcz
iHHhJDWDagW+Ua0K0t0vdddWZJ3+lY+2YAx7jY5KuQ7RayyyzKt+BiFzA4JKRojT
Qvz1tdYXdmPHBAgyItGULlrauSftmEcfxy3Kk4JC0h7n6RTup7rziyuKcFI0NWO8
0oVSvybMtkSZvgKAXOIK831XO+wSl+AlHzccPHKidFnmWINhJDIn+zTFMZNU7KDq
DQ1v2RmAYtSAZcDqW0upgEWanCdAhChnl6/keucQkJ8gsAVC0GLbB06lqQJiO3Mo
eLqKPACPqMXo3ZY872ZPFqGIMOOgVpuW+rtI8n16rk+kCl3r5/WPOUHeBNxAb6Ml
bRI9zqXT3D8xBerFmptycDHWukj1xedeizRch/az0UmG9gUMIt/kgdlCZxPVqza7
1/WDY2XP6xjt+/C9z6aw4af7VhVW2RSOFNBaNAs51Nno2u/oYXulHPH0hYiyloya
FyJkNNycJ8WZFxeQGo/WM7j1XLSmwfp+kDICZk7nHtA5sZVYxyw0ZY09FOW29CPK
tlFj1B0jH9dW6QUhFk+IHMPMwJcxe6a3NNeOmBwrJ6gwz7Pf4sxZ9VZFDQPy6wl5
HIodr6pBg+FMhUq0FZS7qG1hYprs1fqunf1XYu60ocjrBmYFO38VaYQED0VbH1w2
LURi4Rv+3V87X/u7qAefa8ZsqF1pMfC6KFDF6FO2qDjjgydT2Nnl4E/AybirMK8B
O0ZpilOyGdaONSTFMm0bfOcqzVjLlfmYxYJJybhGLfu7aXkCpO++HgDzTWyrw2sx
FYY1BTbAL5OeXaY5Gs9MF7JlPFAsPmNmKZ9A1RH0mWE5D1MJJ9wbBGiZ5COrUfq/
SWkMhaJ6epk8TFZiBJlDYImWwFZSN//mBa5Rxd1umlXXfTpD6I9wtLO/BqoTcZj6
xNhnNY3r30W8GKRaB2pk4XBmbF9IgzTancappg+NbS56pvvPxuC/HL8Sv0oWJ/O1
nBCl6pk2tg1fNKSBKPbhcQqxYWsesHpwlrWfuE0T6Vn1oUt+WMd3HB/MzAd54fO1
guVZ59pjujLM4/8ncJM/cLFX9CLKWZL69MCGdE5Sf1OYxjZVqGKaZdhQHoyEInl/
RSqAJetXn/j6iBXp/kIZ7yCD0c5luhcvXktNJNdXPr9A3gt/QPgz5I8bqaJiElNC
WylC2+sh2JqOnnEFS0H5+wERu0vk0vey6PlHf/cNp3Lu/siVaxbA8Ywsk54nYffH
Q32ujSZPhQq2r5w79ah3BpqjBtbIYjyd0VSuHLa2oKyAHirq46wSh2Df4kKNHBkn
bFMGdF7SHB0G93iLmDwloDzTO/H+rrR+k1tDr7MTrGkZadqTtJIvF7LTxvDLur3t
ST4xANtPE6M813udz4gZz5my8HMOUeWTSr8R27FdBo8FsQYEHyE6XLW1xwq8ahzc
z3Li8IJP7ioK+nqQJ7xXdrrGQiejstjxu45tfO+fgjat5jSb5ru4O2Bd/FJCCvo3
tVW2Nky6tPJ9wz2kU9/KH81m2j0i/ewBGueBA3Znxq9H2sl5S/1+qIqjewxfkTxG
7EUR4X4J7OElBKexJRAvFri9bkjtrPnxNZy5rj16ShZE52p8xXnxrqzJCHayIxzm
3Y7OjZ9KSfIh/xEzIC0nsPFi0s6VeCLF/mL7zsm4hqmUPXh5YyRDW2i5ClvbhUlr
oa5Pe5AP/KTO249JoSz9rOLMZCrFehBJ7Hn3SDBZL1VNl+R4kaNwqygoJzV/YzSF
O7l2UsvmHcqeu3ZbWRjy00eLCAVvcpNYT8/q/2nzZAiazw84t1U5+42ILlUQtapW
lf448wtiSZcouK2vHqk9mXn2dTSBerSUA7CMsm/njnfrkp7916NmC6hKLTjRUaeP
pHaq+S9Gfh9YhLZ3GrAqCF1o/JKHTps6heL112G4G4wwoWJHz//pn7OpsQ6gqNw9
2mtneVFk8JBHK59wW+J28/Sjr73eS1NsVnxKRzYRF13mqY3CvrGIjkhC612tOmJQ
Ges6PG2IyIRXUIxoifv/7D6/DqtSr1YrCC5WsN84j8uabbsW1Az/uroe48ANGDRw
wxPeBK9uYTbjdwX9b65CBj4lxOOp8W/YF6YNeuUKrNb0f+q9T9Tpr0WQdEqW124d
54DnbIkIgVeHntKTo8f3LQyo1sO1C6hNpdLlYKbf0s4wY9pNMKGmAt9jhaS/zKHX
woxrjT0XJUtTJZD5u34YCwio8Rs5jncuCbgIsL3uguKsc2aIh8PB3sWaZHkaDAzL
kAFV3NLFXi8xW/nsdffx3oSDdVc1lhHProxQAXp5W8grE6vLpnEd2es33yRQFSqA
fsti1X5hh22I1Xh4oujLiYkvlHLDFzmwGi7Du9dUG5Mz/znl4HdoZ9Y9Xl+GFZbJ
4qsbPsIxzSzbFfNWCYy7Nq2kas19RJwc3ZBZKCIvVzZ4kUwIKWHgeIauHBfNjave
MSexP6T6e1/g67wfUO0hxZOcNTQz33FBznZYpshNquUbt6yeCBfeBrpFICHKdbKd
t0Ons4DvZqMRSNuOCiyDj7nD8NJBn/WXgRHIdKsxSprQ6yJZSgXpm7wfB3zQrjO9
VE9uobuxVFQiw/dTvc289O+Pm6VsnLtcGFBGgU6Boq3y8/KvDUZOMmYfW+UNyXue
Wo8lfgKmO5ZSiEvE3NlraYIJLXgekA4vktVTuta/Dco9bqc5qeFZwd0Iczd1Coob
nYz0b5jb+IDKyNZbMXErYrdF3aYuskCDEcN+L88nJPOruLr0sSZ9tLgV4Rj4rdK8
eaXBXUF0cDzFjAnZfNLWr6gsk/J+HE5ZqkZRBCZofs9D7i/6FZtIt6y61vaaV1MS
/Dq9bVBH7YkrNOmAotOwBfiF17DZIslRQKrEyS6VGc2000O4dCHmicPleEnrE3hd
fIofp53ddt33wevPtZOrpUPsnZ9g+QZUcPcjbQ8LVuQPRqTiqO5MTNE1jUny8KIC
+FS/0eN7mhRNglHs2hYcDWqxeO0ME8HRqe4z+BtnK1hKNArU7TUuWSf78R5a9n6+
e0h1vhBo925nt63ZfypbRXQslOaXBVO72dkmIIQ5oj5bgq54YQxC7rq6/dvdQ51P
C0vc9oOA+aosp9FP7aHnHms6h8sfTo1IC7AQd1oW+4aoqqVLxboq1HYrbxdoL7tP
tlS9hh7LbVx6NA5Z39T1oG4T/f8NkrSmVGNq5befubNdxdseUUlnEbUHsMXhl3Su
7hxguyMpmGJjhEWisVpDFGwGGmWxZnfhNzO+qLb1a28Ar54cTXChae9RNfTSDu0r
Uf/qaemlGqUg0w/+N2AdSm15wh8HPJ6MnLw4GM8W0cK+wVKhbDvV05BZ/AJqKFQ8
sWeW36a0xHtS+vadJsvfY1XzA4Vwpo27btQE/IWGHqvbs9gIlvGE5l5snIWeicaT
p2J036YAQ7pD+wB7JZBy5Bcx+4HiEdMZAaVcdCKE7icR4vdITjPNHJXGsUXPr391
ZRMTdsiKyBf1/L7LJhZNMz1YrnH4/8im/8W0U7R71EdNv3dCQUb/Y00P2dYqJ+Et
VXZzCfKNAh4P0SLa0wWYEdvpu3MbYXlbOwDSy2Xpqg4GE7QruAszedN/EIMS8o0R
zONW5QojGp0Df6t16vV7NG2y8h/BsH3/RC1maP0mRFHPNOSUAchN/QtvRclEMcKe
QgNfl7XOI687fcwOJJqgV7Bq0JQHssgGjHifOIhdNNTkpRkT3syigeTZtIQngUYs
y0Pwzbl4gFEflIkK9ByIE1megPWIcIRydBs5scJx0TIFj943dPLTaNYhC+W3ie14
kZn7eURG9GDDvOWqtBGv7VVwAEjriET5G2S+WkGGZc0hmjPfb5EAi0qC+0nBJWFd
vgFAnlnNjgu6tC7f51VrzBWK6ezknqoheBlnRtzi2LwdqTm8Wvaha4okUs50KIp3
BjC+h5fzsnyGFKPUHck0kNGBPJr0ZG/+eJmeWsD6j8oeQRpFQIiuibGAyqhBAgCL
BJYg7asEL1j5u0uM2vNs1gm7l50O0bfvXrUsHmwrpK6gZpl+2XABwWxK12IXYdIe
OajA/bucyG4EDixpEpQKsavaEUXpxlLxHzUJ0bHnWpDR6UixU5Irdvkwe9EstfXC
T2sb0jT67iHQqWQdfngsxji7FyZzSFYZd+I2b8Uzx8xnv+PUmbRkHLMNkgLWLzX0
rUjaBVCEeJMWCwIc5qXS/I+f0j0H7TGAHG+ngBoH4NSPnqZclSoRjZExis5Lmo3T
OZp1A5blZnK5RBjJHnfTVsnn+gy/kp5sSbKYJYM/PTLhXiOVaQXpl7ukddKz1XSb
w4i3YK31eQO1nbxsCF7tlEZeQW6+95Qh6MBusHPtBfdIb7ZimDCUE2GHfzj/HprJ
P7suNd456W+jdJGd2sAvlF//DWjiiU7lgnZ7f1fm0ifYxRzdBJrg8CGynOHXvMGF
tNfyL3z77iCXVMp5BJbQIweBkzEfMGfljA4MGkoTHmnTz+CSCFNhX4GUkjOeNY+T
jDeqH0uMSPxiVGywgyuPVyx/xb5CYLHXLBfo8G63QEdrH9iEvmTWZe/Z5UhkJ23K
rBkjU2nJCsuopca0Ds1u5x8Jobb9dnHHg8SVpwW1zHOe0FQPzlz7FDC4V4tgdThr
fs0zSS63Y7nlHlmHFr1QaubfxcSDV00IxifYgEWU7dnmDuTeaH/2aCUFheib+o4G
IT7FelJDCQTrxh3I120QyV2z/CZFtdw8ewlUPHVQZyjS/7EODlX1TgoPpKRdqPUi
rAxO2e0kuDgk+3J82DCV8gu9MkzqqSOIB2BkNjleETBvRH5HNnJlqiPadNPSS3lT
rZm2/3wBubzRDLy0LKoQ7pxznR8dx4pxJf+WLi58S++DyVi8T+Uq3bSl0IleOI6Z
JaiHeeQ8OERLSNPZxf7wpaTAB1o3MTQd/BXrWvkZUXufLqZHHf+/Kxn/2dl9Lne6
Z1p8L6krKdO12+Kmz2F0DLh1W33YWyOApZ/Z/BwayyT9nfksnxIYN8WAd5s/dWfY
wbAkASHhmoGV3fyoCA5ZcbPiTgLiIz/mNA1UsKcBQDMM5wlb4V0FFd7QiVY18LQ3
Bs2IfacTGBK1JrJWxY0PkY9VWf6Fqswe3wDOdlk/ZosLjXHX7KUrVKhxpS9dDMzV
VjbCXNaZE3cQ4NtlcZh9rYJEfAOaQ2858xdj2tFQ9658jbp5Imydo+oj3ZvpIc/N
pIQXLQAiG+2wn/AkmXK2nbJR8kdDR/fLn50YpWtgLSzH6Orq4Z0+yt4RTiqcqMzb
g3aPqnVk2rYVH025R7V4J2shvUrTv5B1u0932EjwnzCnnPRX7QqvGIslFf6q0iJ0
OT/Iz9mXD+soIniccjUsni+zFiI2Q4t5rfYkVtaBxFHTPk8hMOsEmrncVAy/+tkj
0UyloZDRlaXeShv9avWabiSa8XZsF3NnopNL9yv6o7cqmuyRp/CfLilxsKyNUuOS
ERaIj7gkSmH++2BMGPegSFb9n1XlAQyEjFCv08oRhsp4Wc0OqV3F2rMvL+Xpk6kr
ciMic4HbcFbNLoI1aNm+wPVN1etQBjNDbzfQO9lGqmHGt/xQGcXB/6HWjHSh+bBT
lBciJJEQtq0r5SzDxxuK+O8NrOQ8fTxnBnASZ8YLS8qBXHWzustRwkltR8BX3CqH
8+DivNalNNSr3j/iwEJLrg/Vfvmtb+SaiS6ZxRVKPBGGJ8+JhKFZTPT1rJZFViuv
Ll3CNR5lKhNivzZAl2i8B6e2vLpzpxomWOxOGEuN309KSmiK1p8cPYlHpaRYtCOb
8wsWFT1oSWOt3ryJQwgmVGdA4hi3ESl2qcmP+iZw6BPn4oQxSPO57kGH6dCynGMe
/b36uqfR0vNZONcJF5NXEd56er4tIVT9jrSA8HmKJ/fs6ZOtMNIgda55G9mvgF5+
OJflJfZTVmCeJTkacqfK+y0cdGLpNLuX3fe0AJ6/W+mJVauZd3i7uOtfFAgqKkfI
QmOOekFGr8nUj2IBtyHiKpV+XUKVVh+LUdwrvdpV0FNxdNVetHRXBYYyQ2KpsB7t
dUtVUJ4RAZgUYN7NvDd9YksvqSKFgEgPZ6GUatxfymARjFcqTK1Xv5Q6N2ylY/3P
talmFjzBrJMaiHzn3TVbmkCnymqlDzjOWuJy9RvkmCKPq50Nkg7O/UVMqUD5/tu+
HTCoO9eYJ/vxig//9cFROfjesLLZdrgJ6H05nKEs0ZMwyTz/EwYB0qm9mTLLI5bB
LrTeGRqc/EntJgUcoG8BidhYiwKrZvqZjAGx1MoX5mO5YxK2gT+C62eTsWwa2JMy
dPvBge+T+kyETV4trpDnOZE9VAG3+blVbF/4HJWOyNF5UKnX7C2GJNDU3LLReCuv
eDhbmoQmKLnJb5+9Uxd2+4bUPbSLz5BQUjwnkldMMZ9ic2kd4H4veF8Y4kQ/K3+6
0QQWYDMagyJA6PDG3DAIBgKC2TcUogk0S+Q5+liC9yeWoycGPna9P0nR/9LO/Q3N
2Av6psJWBUYT/EasrHg7oO+e3OEXw2fXp+bPnDKtuNOTP1A0ZNjFKXJZQskzGQi5
xxYSXohtXDYN8U5SES1Nb+0CqbXTeX27uYIo7To4EXEqHU5NZPt4PYfLcUKrQXXQ
IlnuGNQUbrj5Tx8QgNccC0wMdJ1JtL56TIjCsuDrok4ultauLruhOSS89V+Twaa5
QehOpx5z5ZSWBUUl/oAauRAjl7pz5kqXa5+xXNVTqoN7oSbsRqb9CgGHkcvFZYdT
+/xQsiabKYGwp6kI3FPXlBDakCiryVAHG7UAKrBjXaQWvrbOpER6XGyTe63ojazo
LHQeHpS1K6JXkKWRWk5GOgU0xrC/YXuyxFdrcAeF5T5ezIaeNBFiyf2iOyc4BNrl
G1rWcR4csGWoUoK7rM4LKRz5EPCOnRF/X2liBuQpoM2G5bkWgJNkzNSaVx94OCA/
LJPceHONFjG435OjWDwo3jqVRLN/Ax1hHge211y26z6S1HMt6QpvKgH2xLNak5Ir
xLvhT4EaYrLsgxwejvAFurBCe8vvIg0kebc2ZGBW1McHTruR/0tuTXbFBTS5BM5w
Zz60WC92IHGKRhvSAacTlXME0euC5DUbXIC4uHvjmn4n5XswFGXyUTcZ4TE5p4UG
eXnI7jNOM31tiFNsgTeZDuEG90fGLtPDf6EghLr9pb3yHHOHskVSJPYkG5ExIKlV
szs8m3fKQ3iAIa/CPn0FcXeNs3l+Nav/F5XYHBiBWp8xXIURefcBVR+27WL5szYh
UHTS2ZInppEtuvNkfxVKoX+6mOSLTjicxceG1dM7nrYSF4bz9KmvDYBz0wujuChQ
+Rcey447uihB/0vrTZjeD4xwKxeffjcp7rBU+Q7/rZ1yIDSuoGrNrhMpMDGEBAjz
84MqaD/8XDLgV6y5LQ7EWJ+p2Ep5GzrmFpvipj5tYCvO/5bOdD5qZ+Wm+t2eTjHG
6o07hjCz8YfFOtp42LykmMsz3R2Qx08qeYfOQghkJWiq3ZwW0z6k++HQNWrteAYM
7aICwuTBSyGuIDO9tsYfTCWHCqoR171f31e3UvvgWn55otThEt43hIr2StbDlZcq
MCWFo35DE5sD00gBy1Uw8jOrbHfmpoOd+/fk/68Cm3rkhm87hO4xGqd5soQYO+TG
I40Tqurmu2F3/AJAUL3W/MLk33burHZ9CvW04RJnQo2nbu6rS8LuvCnm+pfYYhX1
jKCQzn0TNxo98Ysb/L3ABsxc4bPruXoBzX+T6Lkn5v7nAbHcX/b6k3CaAG0hPwLK
qGGtFU6kM7HVsMaORcrt2G41WD1qbhe566aDJsUf9MOrgaDLKr1iDJ9xKfBkzfpA
E7uCRGfGsk5JWzMLp5XFuQo8Pwx14Jk+b5DihtbSlVtIonhcGRPHMtMuwkTglMk6
pETwdWDHZMIuYHkE7Snnzrd7HopDXtMpess/1fz4lX+S/ZSrcCm4k8qiS6UKzFmO
8DkailOvY35cbN/EjUrtknTLfgjdtqlpPiTJR75QtqKBd6DXfyIuwYVj8+PyuENw
EXbOFCTmgn4qnuFpiSx73C//SdW5tWQzDMoIXPI6EWVuDlnh+XqkYVpzmq2yQETM
QOtP/57kmRvGAjuQz5ZExXqGtqXjnpJI8IDXHvJelO0V9w4rM0KYkqTH5O19h1Gw
x8uYxrAU4Xo14cEjOu1DI9oCtrDU80/Np3DP8Zv3QWBC4DdRNulAmcbt+jwd304T
sqX9fs+t9lBo1PPmoXl3GdTzz3oHTjNCc1M0Gw/s6NQtrtYhM4sVJawRPh7KrEcK
eCYACR7RWTWVa2kzcTq2dCv++NHxil+900tiORybQTMr6+sNBw85FP/1xXBhB5ip
IWa/BHQsLmtuvS/LjRpuEYR48fkBqyKmxRaws24g2M9n+ZDWlT/QE9j02L7Z5hze
c729Gq75wVBkf4gmy56HpFHzqolkV0/RhZGSuvoBdgl0i/iaKz5/8Xp1pzOAF+gK
JMsa+MSEUMegOfzBezgu813BKC4JlRSb5EwsAvtBxS2dlEsct7v9lvm+0zIqb/Jq
2+ajegSGjSvYAqGhiywlDTQUYX+0bJIAB/+4MVHvaaTSdg4qgbpLY56/+WtugoQD
x4TBH906Rlmet7ywr2qadniV18+Mekt5ohaU001WU7fOY18art4HqhIZYApvRlQu
7BPUztdvI90616/M4q9rcGj2BlvFkMGd5i9lhMs38f+DYcx/jVvohDYpm49ss846
5OJBARwEum2+jLBJaHyxM0fQfaL3+rPEI7Og3TX9nxDsEO7S4PqhOY3GECp/4nAW
IQvNCgFhvwQa56nKWwTdUtAHhITIBrvzACLvVSZijWSECtgnvoeTqDPIyaIcZzvB
Tfq3Q6VJyquhk1EdRowAoCldF3f1aGO55qMsMAm3yqlrM0t5qdSk3reMAkdu2nrT
/hI3wTYfusFVn6HXt0Sn877PteEybPAJ47ZZuRE2q1JyHCZu3iCiv4o30qTsyoG8
KS6lEIBa6DwNzpPGV6a9DwPiHOfwltbcVJ05lyITLbLXXUsN3EnduA9wlPy70rFj
Jifwgdw9Wz21QTfSDzMeGl0nOPcIP7Yuy+haWsXMTLD1O573timylrtPr5km8aAZ
oVN6YWPcb+nlx9fLkHFopgjOQtVFijLgNiPL9FmxnTe784RShWlKkfJy2LpcDL5Y
FpyoPVV7RFY87iZROgWm1xY2To+U8eL7dCBNT8Oj1pfC92YM8vwdkfiKcOKBVvdU
MAXrq2qwVtvNiyDnyntJz66VvFN7kw6JNsBX1rt9a1k8O/mAPzm90YDhS5yTBVjb
5BS2rTz2uGaBrsNTT55euP+Zxk8MyUxiS7UN0jNm9yqrUymesQPDESpWfDg+JxpG
32AFKZp33AeMqFD+hRvrCho4/ezvm24W2SN6NvDL/GVzphEz2eISLuIRTeg36+cK
3ty0dvc8ghpIOeVfc1Dox+VNo3qCByO52O8egFOehxRLI82Gfh3pIyyOxyFeU734
s0VK3Dvfq36JS7houoVpEzFpKdyqdh8yEmvg6WZ615G44B9yeKDUgQJyfoKLeWBz
DpgY1NJODofLIbT4VXFdkXlUpvVC/+JQXPmLUGYlLfwGnfA8Z7HxdqTiasn1qaHM
kU3IoQEh9ORh0FK2xgM/JZP4q+pL3K3AD5+VqD3lVVMserfWbo+qxxxNwBbMAQ1L
sPbiIh9VnaZGAoMu+f8busle9defpaleA+yPr6gs+m31LgoOzB4vvfuED+9FVeC6
nUb/V6a1TXdIs78oty3xUkDZaxppSR7STRcV2j3QmMeFyl6cGigyeYCmEwc+DEt+
uyNV/C27DvIYQY6qSvjKHxH5GH2bRwVc4rQv7y1+4hIPQ1pe5Nf2C8irf1RFsKLC
Dcb9qj40eApJlJXNVZse2JMrLjp/XiXT2hFrMzSLN1XsD3qEcI3yD4PrpvNO0uFQ
yISzyu/BLqaiAP11rCny8wV4+BIqnVt1q4rxt1dtZfx55kzJy1VwMXMDBQOQfphr
4zjn3APE0H6n/8Aq/LPkO3ORzeBybWCkMnmT4ifMQ3M4R14Bl/trRC3NeMWmujMe
wm3UCepYJReZIx7wSae2uCzpJjNnUTX1b1bQH3ZI5dwE6mGPVv9TnSa8VJE8PRL2
jlNOl8FJxicQiI5hhSlWyrG5S5s0fNaMVqMMEIaT8pTSfpD/M8S7yW+HiH5On/Zl
yvt0NVORoMHJBx+b0kNtM+rA8h3T2x3yr5AxLMjElEFWP5JqAO11p9fvT3PoaYi1
yIYVgQi/xdzeqS0jPUntrXI6y9rmL6xc3/AmJRYUdKMZUgNnvkV8wrLKPm+6OyWY
VoFAv+YBNdvrpiw8Te9zudvmu1RBDoih/mXj/SN9fTDSPpnhYN1m9UuZD6JwbGLC
d93MpZGz6ZcIF3Na27tCLKxH8pUalCuhyd7FIudM3pcF3SndufIeShUADkcBcAzW
Bxc307c/TRPzjDeGN+BmkAyHLDOXj6dg3nu2p0qeeS5N8s14Mzfz+fa5HmoJ/qya
Tyc+5pfkvL3RHhB/19tF9VuyZ2kk/PXeNmw9Rutxbo1qjIZrzHW+5atJ9g7ZNx1D
yGZTEfNaFDJ0ZgiD6wESEePK/VNpalZbieFtrpivJO7ybo1LRmiFHg59QtDgK9BA
AWKylmrEsRCXsFhiKt1FtqnJUqclFECHpV7vuCfWTZuZ60XsDn22XVGwV8iuFRZG
W2qOxGE4iiQbSiQ8iHOh26Bar2iuZum+u1ies6WjIlh6B1BMEyygEZlRybWdh32/
YBy9hcA/jXJRwDQ2wIbMVntOkmqFXu6cNblmMm7RqoWPKqH6QBmIlA8KASszK72Y
bn768AuShxMPLaHTTfYodTy9gEP9nCc+tvYAzj9aSaTW/4vfGhNsRm7XCk6uMq5j
wgcezCpm5hUmE/4Mgt3fCPzlzKjsl3vo+igc+Uli578408X85V7rXQxR8ZlTzm5Y
cVb4XPzuMMKilDvQTfraKjkMdkPedOQb0iOyO2G1LVGwhkkxFxP2+rtFDQMCtWeA
9xb2htKg5Pmjp1waY9BFlgQFLr/BVM4rh0c+WTgxqyCTzVtD6FwK/M2JPtNelnD6
aHKKh1kfQx1/a2ZLjZp7efeCTckEOeH7uYl2wyVakeVU7IGInHLUWBAEpiJGezGQ
YZbV2TmeHdu79CjQ6lQE3aDxf8cUk4ExqBkBZM+NceYyWKgYYJ36DG0YkseKnztd
Bcas3raN+ejCpw+NeET+z1mPd0tVcCdz73dtS5+kBxFd7a1SAIVDToon42+GjqLD
k9O/YKR6bfLV41KfSXpNgVdPlgB0WTLrrVEuOZwu3Mtc2rPzYpXgggkxKvbNBt54
llTCdg0lrlotBjD8v4TP2E+Ac7bgILc2v5K8WZ+j38gv37HrWzj68r6vbhDEpLsK
NYY9lQuAnPeRvujBbgflMfF2gvI0cOJ9Ar3WNNiEGgRCXbp1UPT5HJxK6iTsTBNH
0EwEkOOiCI95Gn/u9kCCF3lzXIF91BKHlAxFzcvt2KTK9utLxg3XFWQZQb9d1eIH
mb1w+eUQ8DE1zHZklMnZOiWq0M3xs6oH/2tT+4ky1NR+LT4BuFbe8lXpfZjmr8HA
MM1LioXXvtKntjGIZv1vqZkxtPfIWApvEBrb39Bty4CW9aMvxTnD//42149g/GQo
bgj5PHSPyQxJIo2aQ4VLl7X5Ai8rcyHXlExxCI8uJTxUTIWOdnG9Q7Yo5enlzK1e
qnYJitafuBK7pUwEBSrXTEY335La8O4+fKcnj7i7TqEdMBDSNDcPDmSET4a/bmck
sIJ86LEpQhwsqG7Z+6hpfSkIWzylHnHA0fEMA+IT6fNQwI07ggFMI+8N15mSZV1v
VQ9Bdj//uewbS+IjfR0a+jboh9MPUtBAq5mvpngFz1AjXOYAB47ggA/KZNUVXk6w
qCOxZCBu+iXuDMxoCxPeRHPYOKwaRKwwz3Fd0w29YdGuG/a7WcUx1UpzrVkukPog
Q9MMKob1CkZnQjcNy/znc+KGnM2XFbYjvOkl2Hbc6CiIcvBn7Hm6IIsGguDnRSrq
CZ6SClX+QkmrmOhwEOjHuoz1svw/6+EwORRv1TZnpCSMRPf4VVQIfKLlCdXN935P
w3UuJo7XU+18Vct+ECZEklLIDSqrYvx2Pj9EQrbqe4qwwiaqLUp6JXQX/D2QFIfY
XwRXik2JnryWOLrHcngMQRwr9WWyO+lDEBSez/O3WWXO04hg8ryHubNopj1cEh4i
+QuPFAc0HQvX4c/Mw9ThLfpzV+thEzPwEBA/9x0NXqBc1P0zqGTiqZSVzuxSAEDZ
cHOWJw0AifQ+zhZq32PeFf5LNROCwQQoJy1mmba52NmhLkr/kYmWTF6v1Zp9/ZlC
gjxjh9sL1USmRazZC/7wnlsBqnmk3vAc3hlksbGKBvRPDIFQlllesU+F8cwFU9Bv
s1DKcau49TNhM6IMUpGYiybwynnBNlawU6g7y8KnGaVj/mmZZxKT7Y0afn4p2M7J
/6M5+8C/yXlXsW+1uTUJcAJaKa0wU5q4lDyU0JQclfDDr6/Scg3wFBvQUsc+pegb
rcjoBiEYcysU2BrGIWo+ZCmx6Nt1V/qQPNV805BhcwpSgCtfxwq4qmRDc79bXJYy
S2PSJMTr4bP2PTYJ20DOxSVpPbgWG7YJilgs2ZMYpjpy6Yo6OAgIhvL+EbsijxRf
V+bVkdUS22eSIe1Qs1ODp1hTLo3JLUiAt3uNz04dgU0Nl9ozSpM5Hg9QdHw8AtJ/
ySMXdAPs6Hgtabb3ValvxZfJBZEvunkSsag8fT2Ghfwez2hIUKOh5HM1/7utYTHz
NRtwvutpp+Ws57LLc2F/awQ9m9ymYNOv23is6ozVXzyVUvgwPjMs85t+Z6dS++ih
l0rWjhyCDQJKFKTccUewfjNjhHvjUPmR01XI/fX1DcFWVGei1+FJkQEuKdHVV8+2
Hy6ew9Om9iQegNEwYJOlShyWVYOoskdsLHglCvynnENZMBqryoLIP9cEQtQ8Z6jw
UBYB1CFTR67lOe3xC0bLjLiJ1zAfEBUz1A74g4wWAbHX8ex/sGrayu21yn5L4BDl
wCFaD1o2iEe4nJ6joIiXrhAYdilAb2jSS37ZrPT2HZmEDd3Q70QC4JmToKAUmSqn
TvJizaJsaDwJoFmERTr4TjtuSckmVXZN8cCJU2/tjKsWVOqGxmGRil1RnRPxYexi
U1vw9rqU30wANyAMN28UUj6ReBiBYf+hFrHgSSkMRBAunX4MvEwieWWzvPs57PDH
5kCw22WThW7HHXd4QMcmmVRQsiT+/ET75g8GYsX+ZuNRpcSZEUmvu7n06oN4/p2J
OmOSczebrATlXu8OWnN/P4+oIcIU5vw6hcPwR8d6GEvGw79RsLu5z8lOcqN1kqOA
e22Bg7oXYbn2uRbX7GEHAvX75hx4LXAdomsS/6YWf+lySwWnq/lNeqeFhTPpv5wl
4KAYNX0jjhYN5PrSrqJtxiNYXTftmV+3KSKXtZ54t99Auv+IFmOOSZGTugAZ4IEZ
UAVJZONnjUnFP8MEs7ow0YTq3hWT4XsUIi9iIW48ZA+CQo+ia8l9oh8qJ0e2nWGG
I6wPtpIqFbAS2GVmN3gG/0+lQPSqLtykAKSSJEZ3E3m3tqdtmcXofCL/nGdYQGcE
BXWlhjOUC3qDGaqD/I7Yugu9QbxZdxQeJ4SwT65WjeexLKpCp4L38SfpqSc7JAQg
YP4jhRcEoSrCdKyoAHYanPFV7emlcUGCzpvYktd0ZWyLNv3I6DWLx4W8rtzsYfdR
yRbIxUkzecb0slzburZz/IeknzK/x72IRooB0qbcNPtF/WYB50tGCxzVk8taZXLe
H5gNrEkHN85TDi7d2S098bZygCxHw5ZGYxnPFG+Wt0IVs57gbApDydBTe8X5njzY
47w6vviJd/lqh9oWpk+EXzqLa3MJfPLSV1wGNpyOdhRsJk4rNTOcrjtxb1BNq7ta
YUGaoo3WSLU+8C0I3jfsPrOcbZpbpLy68Fs56MZ1dbmDolzvcmX+K0Yoav2+ehSK
m1NFm/2hDEsjs13i45PpGa3XkXhlGPUAphR9RXU1+PZv6NMf5GdOA/h2e+8+WeYa
roDMWRoeGfmdEqHnHtabGGr4A222Vmuf4bQKf2gO84gsfvlj/M2wyifkYn/Wlgb2
Ym7KBnnljiAYfzOJHqb2gLyIaTUwSzliqKGPFhge5A/usgWvMiOahz2lDyMg36n4
/UxyFhb1KXe4dAemWTXRhxOc8nA//H7bfBK0cRJmm13fx3FAiJ3tw0ZI/dY5vbW5
kJI/uvBRTJAK22TWGU1KuK1fdgdcnD7TLr0gJIqobCIRvm2IdHlaiUDa7P/y7mtr
2qXHu/P9mJ+9a76Qgcs4jZ/WSym4KcPk+sC+5D3fbygtMPof0rEmqf23vo5M4h7s
hhPjSQlYaEqB0E+vURM/V0EthU0UMgmtf+KNrQJe/URKP/J049rcrWGtYpw5yjhO
z1/0fmwst5ouwjeJWt/U2WF0yR5Pry6z35YjQ0lHOcbjE8Vx6UCoSbwKVFpZoNWw
Hupj3xWlJKyRGOmZHV7YuOXyM2CCsjhHJMIuvYnQiNZlmHzc4x8fL7KDCksaVAxt
LS3Y8wDDG1PeKAVItmPF5y8jcbNK3qhqAgGJu/nyJnDLioWNzSWFVuTmeXB05I11
JjSXgPM1ZjAvokoZHmhxo9wMOFTBGzHGXu9VkkLhUXt07Ar6oZXRH972ShDyAp94
DRZmdpz9u4u2+yTfH6cfPdM0bJUhs27BmmySRU6GdKreykCnqy2p2kyv0XsOlpKR
R//dcJ2QvzDpLDV93IJO9DG2yzoeDkBUmBQagln00nKuH9QDcnEUUXWmHVUodZsI
DGVhIn83SvqGoV/TTct0FHaSym8nZp9cFAGPPl/GDYwsOM9Nm7aLalInip4oB+QN
bkhkSJXNvjbGijT+wjsVL1p8nVuBJByN5cJGqEL/5mPgYe71FWJK+pOeyR/CYCvF
J2R0zeqsS8uFWz4vFAv7Ig4Ok5YQXxgGU0i2KgvvYinR6SbeD0fZmxnsnVmU0NVy
b+O8X/i+oUQkgKStm3r+2W+aCHukzR/KUKgXytNN7Nmog3HllWe6m/UKVKaZXuO2
I56GlfsA/XQQ5UR1UO3pQUUhbQmvMizm7AddEAdyEB69HeI8FocsWkThP68tXne6
q9uX8AjnYq8VVSJOW4OTSIIxkwlxgZx+lvJj4vQhx2Mx4SOJJlbFsAjtdPNHvmyr
mLAy43f1bV8IpYZS9HbW6fgAaWVhSflMJ+E4eq43hOBoUtSYuqHkg3cBoPEZVj29
ZSXNcE/eFus/b8gBSV9rq3HMrhHvPOdd2n/1Kqzej+aEtIjYWQ4pdo2Zny78huol
pqpa1TsxFA7+VUtkF6d7hOrAmQVwE2FjK2LL/91JEcwzF+jbEMZS/LDNxGdDJyxg
GGDEuGBTUcgvrNUjVkqhMaeBiDiuPF7dA7LXhk/bpbIcp+X68UzKy7XKBZLQrOT9
DDauhIUJPrOI/+pqwz2IbkY5tWY5aihyiqzJItQkZUJXv21Gf5ju8hWxhQOlow/s
LpvvHeAAGKbXbhgHU0AHr80yOmcueuxg3yEbgmQdPlscLD5uryFXoFL54yUwsWot
HTdIb+/W+WktTRUWIDXG4+S4WNO5aTWuGV2+9zQsbdAoyNuiAhdcCRpNxHxyC96t
nJ8rLpUxUZXgd0NUB+6mz9b42paK7LJITGL3Wufvg9h8rZz3UQA1nyE8n4UsOi8v
WewKi24eF9enhdg2MUKQpftIUoKDGEaZLWrdwGwB686F/+1PBy+9IiP4oUewB9mu
QdjInFJ87PpRxAE4BWMjRPHDGvI1hF7e+TijQY8ZpTMsEkP2CM2/I2c6q68UbL7c
PVaIBeAyxQ2Nx6TWW8JBPItKMvdLnKNLMbEXSyPyt7iy52NfA07G5PQU8tWJUYVU
HencfrQpxZk5b/xtniBpdjTWuHyGuizMonD++7+ws3IYGFKIdwZ5+AruD4Z2NZ7u
uBPvwQQzdFjwbmRjMINRAYK7tai8ZttMRXq4GtFWzny66wXUVO/wMKE8FHlsHYFI
sNGEiVXPGwdORmcpis4evoWwmIzJCoZMokWY5bY6WQrp7Zb5y7THqO46nj8LCFye
Uqyc8EuYX9Kb4nS4KfOdSXvRgH6yt5wi7NMxWFzGnD72t530MrK8z1PMt2cGhJ3u
qTFlKjW0AL/xXkNOUWngZSiyCT3IiWiyd/DMXjVE6KbE58qdTqkLTpyckohr+aSG
nzFzprl6WtXq1LbZ8nVbKAvJ6iQ798sJRvX5Yt2GSkzDqhUEGZTWk6eXvijSuhBX
2TMYnDRupxXctG/K+ZDtD4vsL4YRWaL+3Uc9YK+GOumHvvF9anEbd+Ob2stvBqna
+/DTkiH1qmMc79+vV7texhCVIMP97sjLen1tmKIUiYl7lmBkYSzJXErPIrS6kNH5
Tlk/Lz5XzEGT2Hh495mdV7GR8cdBulb8SkTbMBL5Z/c1+21fuskrK2iBZK7I1da+
VHmVqvzc5C5R33lPm4hSWhABPB5qN+HnTJ5Ylu1XqdB2oyFY64LKBq3cMum2djE3
SXHGrBuhHpbOqxsczMkSpJn2fA0XDjeN/7+WYLzbTF4XTrZGh17pUJwFYUmdRvoe
uWK8VP+jvUvrD++dGxRj2GnxU2J/Dz6WX+LjfZv2EbtjAdENPQx5TKk6sB06xVxR
Av9l07daK0hDW2mUnV2LazRevO/mQlk2NBmcXC0INnhwgYCrpYDlBNPSs0tL1A3H
kfD1m7ZIJQYIjt01WWZmrGgSoJ3hypZfajJ3JLP75N5bweQZDgFDo4i6AAX36fMm
5TsA3tN3QjKlF5cHRq/6b/os/j+S7u6f/ewuJQGx1XmSqfyQ1HTiZEcTIRnjrMDl
yL1yAheWiG83Uy82/i85bmthB8BM+a4nR0llVelHBB8kYOmtR9DBYUyGfwgd7aAd
RkFaVGJYIpIXTzxnmyfHcskxbIcuHwfFLKC4Zj6LCpODI1Au3y77hsXwYwxXdANp
U5EGgY8Y9g7M/M95wzPe/VmC98FAHLknm+mjJrhz+Ii/nZV7drpRfVqoFdfVqZZ8
BvJgfEaPHYZUkhk2ZVIDKm/gz6//pxqR51m9na2HPPNVi8A7ZvRovTGGiuM55KVq
WYZYjIwTovlbZfAxwMO8yN6/BTYAEPf5gi8TQaEmphQtqVpgUVLxgtcZ+g73f/T7
a7uFbsnGUcOj8fWpcU5nyHFZKEq3ZJoAgF6KuM8MPgDwwHaSD24AZaEszIf+HMlH
PjrRab6mB4SazIj905GVbJfqUYxJmxVQ8B1yDeAIlJG8WVwdaFUfzFs4U0GaM9zy
4KVl3jUcC6VMtGlkb+aygy5EqSyLzh47u4OK94oCXCjyvCwu3pZUUI8HTqILwFRV
L1OoNcTvkaqm3UGUFlm84oLxguduOFonLEF8dj0+ZvoHXh+Ra2vuiUjFMILBJxwl
qRB0bw+DM3zQkmUTHkPeXTcVBak/iWokGcPXb+HgHgn9ZkjBdD0I8OeB2pbJozB4
eeBfi4rNe7GNhWxLneWvoewEOrIirnEyBDxM5RuyG7sXa8vUpCb+OCvK2x51ZpG/
bnbA0rTquSDsZpURVAjvtQaxZdNDBXhdbizRrmrfAjuLSuKCSPmh5MeDisp/pwYn
nQGpiJCqI4p5bRfpdjkYStj2a6WG/QpFcFSpsWAzF6c06/Nt5ssZetFoZX7bqlUA
ovYMI8h4zX7e/o9xFUIoY1fdGI1L49FroFzFY7rkbhZCCRu8bVGsxuCY+tAFZ3zA
1ZbsRssEAra7ERuj1FLHM7N9XgnBQnDQrA4NXlLq0jVDs2+8La71BAugt5sdWUPf
cUyXiuikF/cuNwv1dQk7KwSBeJBtKmEe7MEH5oak/irWW8PNvqA+o1xhGohhxkYI
oMyurVNE+XE8JztX/EadZAlo1kl/Gvt2w18etfcbSncs7eb1P1e0u1iLzVHRWWXE
BSsyKtuIkzxOU153Mau3TRl4AUDVIk5vV8iKw6/FJ/JU3HuzkAaLTq2XtHb5NV2Z
MHOSQx3HfUf/wCqmH7DIId3S088wKYqfQpEuFHhG+LzFIucsJYDVQl23FRjLaNVE
mFS0pTxySJGhvUMGlqrrBMWrSaP4eR+icrQPNxJ2cHtKFq2LXZ/AQJfrmuYHcQ+e
b8qZOfl2sMeRgONQEgnVARlA8bPOWj/MEYKQkSJVAia02RntLhsfZHgTaj/sUrE8
ITY7m8e1RFtqvgnR6GNdzSBuTEKnPaWN4oQ8cvb0auDjlxVdSGvpWg6BDggjMPgD
ONR+RoMZOeERS5wxOC5itEvJKeLb5onxmsCBkp2Z0qDscJlo099nsMC9s4Lu8Z1x
B9WTGaCu9BcT+vBg3Zmf9RojBKUxDI66BC5P91ZwE5IDgHx6IsbV/RbwTu6t1Yrp
Azh0lowxSWmDt7biMeDVl4DibXGRdqlRG/SLHme+aCllQwlCzxnr7Y0RY98Xw9f1
3jEMy+Ik2VZjgPwr68xsVM0nT/rYfIt3EN1+aJExEk4QU7JUCFaFTelCSLEvVKKI
Moodw9EGZ/iVHmzfVqueVHBsYJu7cyKcdtLDOoQvAuRj8EvbwWg9ZwVB87TEQ8RY
fPKMypSyWqUBx/VpyIsE1k+qWxNaVPkYz9rHrbz0HAF5ZV1XGh0YrOyvpUiUMtdx
nBY/i3GZ1QTfUa3DRuc3dzv4FUkd2dR7iPoa3uQB5SrG0HUeC4fqUI2RUwA+S4Vu
PPvYSEeMpDaAwbwgL4Ov2MJ7USb1zyg/bNOpA7S1b8rGutXtqorSuqzy6F6MH2lS
9ejj+6Dn22vx7TNwRStF1zUGM55F05efna6rHMqGh7LtXDrrYNphqeYNMix6/GTG
YTMJJ+9c73cUBu756n86JntRlkuT/0J/RGLRohOWpDWYUXzxy8HD9PYE6xMP5rMQ
Gagw1vdGeEz0x/twSaYWfYeHtASk089/UZmE3geQGsyep99gYZ+rTJrVZ/o/Nh61
yDzeOozSUzzDyjJot9yRyq2Y06WUA5+ysJFi1VkfIumlMlzPHkMerURLU4VtCzpc
IsG4C4p8HAR13tWC1yODnGP+/mBwpk0cyUR4s+jmQBRF01HpRCPrrAp5hYzTHB1M
ILtA8/SGDQC1flctDKeXaRoXMc3AJ5JDGXzHuDg2aOfDeUmnVcdDAmys93dhC8xZ
iEjIrqFLKn6WEYHU/Y69K1eRJN5H7u9uB6M0sN5n9hYNBTOcH9CDGUZpH1K4ePGV
QrUHbUH2+bjYGOodmZqSM6DeKtpydHFECRLigRyKiGGZ2JOp6ua55+wCnvVOwklv
EYqi+NKcIAkUKNYRZ17QvaIADPYlvwhgrk9/ATLWcdGb2kqiFssdZfJzOssQ2ypb
PD0ipjP+RWFJc7NZHyb+VXooRZo0eP+ENhyx/QrXea+13u23CdResA9D2uGvDc4k
QjRwtJL1sYKd29R95gD+KghCDGupZlXdZO0usSEoLG3YVIT9U7GxlneJNLjwFNzX
WeFl0/9Tc5kOTMc+alL9jd8rhpLFKM0SgV+7MwrHwpn65plVG729MPMajITPS4y6
vqSzHLQoNRwFFJV/n7LEugAf59k9VcqPtD+6Sp7BxVCn2VILXdmS2JmXEHgU0Xtr
Mbmn0BDD2eFiw2NJI7WkdM6NRb4YZ7munV2fHt8VBQBMkD3kHglmoZPCbRRZYgVW
IofHBlMrsjPNUhXoJXdyzEseNLgLk0JdbonNMRM/nrv7A4Ut3ZKVDZ5JEMLF+5Z8
Xu8wGwX/yMCJk6bkjxDYnWfkaeEmQlPZ5nliOFDV8TdJpi8qjkTlX4Sh6+k+s6BD
znH/gRJI5/ZzVRB+EYdU5RM4totntncPjX5qWBTc4L/huiyMQdubtqawUEEcCWS4
chhtlaWN4VKYziWyZ0mXwD9W4XRj2CMD/+ydKW+GDuDx5SYLGp0umhWS2r+A7CLd
uFCBTnQyqE2m+TSlN4NOvxcSqSmJX3xJCqAxyOiIcuPtHhMuuVeoXJ3NCyGEv+g3
984UgRxlIfucXaspuvFgizOyyy+S5alE5xWf6YHwqmslR2Hzcl/+VER2wnoG8QKT
J2eBia+3t3X+/tn0IqGupq3zwmG0fu0PpBnHOXqrBpsoxdX1bvzek5M7ikvfc8qm
N6IFe7cn0GVl2dmOAgWYzm8I23w5SKVXm/guNJCF+H+WDYxgFK+tddGfX2PT/h0x
cpZ+R1xzZN5fI2HS48L3hohdFqvrhrk7avCO8xcniIVllhIGKfia2YM48UHqoVSG
AhX3Zd1iqBt0EWmWtsXMU6D6XIMnIpGCIju4t+3eeagFhXNuO1jE581V7u3dh+iR
1OxzioWGrObuarX/IcuxJy/4jVxLjBVXcG3X57UeldtZpwleFQ3U/4tjgFOjEooc
Xh3IW13Bu2MeZdC36AtDLfQ9vD+kZTPXLYHHdQJQF/tfGkbVDpGioA22DDJNkf56
kV4oBeOWyDBULf6GbJjEjLgTXBLdF7ZctPLT9N69ILAI5Ndwg7pabUnLA6d8FX96
fpfiy7dvomnW2ChTfJ5thP0qQhPT6W3CFX3HA8TdFjNBtmuuJ8vVxmaM1n8tKnj0
sy3DNkkXWsIk8U6jJb49RAHmpKAC26XtHthKMJys4NG4G+I4JcMR2weis3PsYPYJ
QAQX1Giw7RRiGUWsKgBWHhYS1xkSKpaosvQazOOLG+LljJmwJj7f1FokeOfNxSZp
PicFbX+5diuhr0EJU2BZ4QO6VuDmw/eQ9NHlWvBQ224ywdeE2gXZ4p8TCe8+/mj+
ESS0cQtbzCCB8+R6XCP5lk5hSE/auDkABx0v1suijDAe6Gf8OE44vqHpNVrdNQ7g
WTpKxw+gpnfgCEPHiGizBVBGd0QE9D7ogdvNIVTq46Ya+ce69FBDXS48V+jmK/Xn
NSjluXtgmtOpq7s35Af02SZXkdKzkfT9z0hesAA6LTZ1HJWzIOYMbsD4nDAptjo9
MV9HXajkS4p4TKTVKhN8a1COVlsEz1Z4jxqe3OSt7bl7pHeOrNsDHzwQ6jHdfMXg
TTzbOLwiEMqlYaqBobUopzycWYN0BTUlztsu8Ql8y9XE0REpPdnLbkGnk6hCC4rz
L3SXaC8au5PTyur7yzlL54P38SNS5pkiD5jFDLdXfIGI9ox7/EQiz2kJn4I7ho9I
4bQk+yxk5Y+LnJ7GVm+GfF73JRm39NyMGdUVD3vG5SaLOBS+niPPaiDRBOjLe6Q8
g0W7X8gAsE3IdmyhZTtElk4O9rjA466hkBoR4hCjjuKl19/a7QkzjKzE9ZZlXi5R
PRt9YcU2Cn6x4rINiqkU/K1lBaB0ESRrc6WTCDr8vlvrZh+hWGTUdOXDBRliBezj
j0get4jouBQjWGQsh5vURow/retbm5pIowOM8x5pOsu0qmuyMVf1AbDFzjQwyaJN
BUmVzPcakIiUnRaYKvQ23VONmvg9hG1nwiKyvzwqG7JWOG1IUA84UYG6Vh6Ggb0c
5HY8J00vIydwOvlfh7riNKQ8i7MNTDpeyL8dF9QJ+l+bvd17rV/zDEsRGuPH6IlM
Lyv+aPtQZ6ITnpDuGzfFN1V0SFuUl5M/Pb7LdX50AKtKBaS8kiMLYx7g1CcBjT9z
xhZflO7p0vYlRmWMwoS3jz2SpTuTOspoiSQk/eWzWmB2fzAOlN/BxlT+ODUxHjjB
pK/OW5emNXKweXZH/YXKwIt1VxKkX+wU4RC8gXDlrWOEu0hBNaV3RXa4tDr0A2Ry
Qhd01qZ1A9mPI0rmitlP7k8E04UH1hqkqj+mcPPLpNFsb9xqXhFhhI0ImnEii5EM
AbRFXCdxAO8xp+laI5n93n8ojkO7QeXR6JlUqbmxCs0Xa5a41CpA0kdimvnGvjfz
OaeOq9bhXqq7GkKdLkVXyY+QV14oGI9Z23KRLboCK5/nW/2F4IHFj1N+oG8RPSe4
kDyEnWXpWirfVMKgZsAxSZS2WG7dBn6XdBjRNeMP3yeeSvgCAnInNGapTVBAkLn/
6DgyMkoIWEETzOukmLG8URdMX9LvihqTvRzBzHKiN0O6etT2439AWqZrp2UYVKsx
csyIP140Mp+lSx4ODhrUMBRnSsxUMeuBMx4bi+O+/U1JINDYUk9ue0p6eljYvj9q
pxZ73WwFuk4v0J4tGt+WKgk5Is1P7OanihrTyzMi0DBoB3q6c6V8QFMbUZRYnuwI
ANM7JyEtz3eaHq52y8rBk7fG41qT04cFsqBubao9cTt8+j2OJbLroYicc3VNf4YG
fKkgTyjC0bl6fKVBIU4EmVoS6tP8HW8egsThKDPuLSRHt+iJKF/j8joyiWMHb09n
Z0Url9qO7YKsZRW+2Vv/7LzxDI5NwbaHJ85GXtzDr/7QgJhhCCaRqP3gYZTH+kmd
3GTdbybk8PIQikvS06vVA/ajWrNPLU8GKvkYbaXtBg65NcH0aa5UPw6WiOjXhgYd
oRe6gL2kGUtScJJHPocyk3nbDslFhmJPE0DkJ1I8vjqTNhmqEozEi2XShZlWrTVj
sCzhjlpHv33PwTqk8EUw63GuZwmj1rmPRHhIdqnyMxdP5Gcy0RaERVIs9eFD7ZBU
ESZntl7l+GlwFRAKjJuOF7KX/F3Li3ptzXXhr4xpj2GaQk9lA8JzdTHYlSbZd17a
yQI6DaeAGMfvWDaTlKR2YXWb/+nmyLzBdghQ+LgRYztCTTlnqvN/2H4tAFWXQqxh
oo5XjLSDcADwkSoW3hhJjbEP//EBm5zbuIjrSfQXCGk2lq7b/vdNUSWqxDzrJQ7Y
Bsl9asAFtj3wzw8Xsd1S2CP8O8PKxGINHgXnI09dTQea5R7iNWlf6LnJQQZWo1w0
ilBxiKYGAuMpBDGRL0qdQJNfRRVcuAAQBBrhcfZVIZ4yjF5TxLldy6k1H5i6dJ8o
CKALDZDUQi/IsXdGjP59nTxAUasNU9XeOgedRqXHfdNhMWn704HD6geEcod8gVpO
0vYzCpt+WlaSw5hJzX6mftg5CKHqgK4nSGkdB+KR2aNk6RMap223ERsk9avKUI/I
pFkJUglz8KLjcvV0QJjMj5nhecgmW3mRnavtIjkQ5bF/OrDJmepMNDJrzmTHahVF
WmbAUoHTD2PD1GLiF/7M4K5kruQFmysA+md2wiXlsYUOj6TntFdI3YJBGUyFk4se
yRro9ImpGZAKhki9FTQfT5WmIcrfTVwgAWlOkt4TY5grNVmtuOFxk9YXmq1LXYVC
kTw6inZkprNer6vK8N8rO9nDu75Q1gkgpEW0VRE0ct4p3Rcx7smx7OIiHoc03jSu
btabMSSU2RYRY6fnixXHASgb3YrHGZrMgiE7cBRfXqvRtGzV6OiZnDQSYDxyH8LI
QZKqZwO/AwbwkP2vf15W3ioihdAKAd1ZkDN8LCy/wo3ki8IDwHBGnoD47eVWNZKh
3ZmMUTSm8/AQb1Ty9eVfSX6MH3vr+VpBrGKxe9/mGhxZigPocdyHRIwJAtCjMXes
tMcHDRRlXUIcgUZrfdE7662g49pl6/nKV4rKBZbKZPQLANI9HV85GYOoeVLgjk7A
T/ZN1cSGSAUclkgG74DKbIKx19BrRx4iZXHx+L8zzPF5LI8RVquu0IDU80FB2nQ1
KklXYGxQHoeX27j3vHJaBGT9CLcQDTIJAQlYHrMIOGXB4mcSo3AiaeiVYWXo/2wQ
8Ln6pchclAn7tm+mvNrsnIwGS5Dk8tw4S4r+9K9ukp5pQPrIdZU07nUj75uUjRKZ
WGNxOVX6Cf9/E77OEaXxSCmxHNuRBNL9wgIqiGzFpYbkfKXZA9S+NTHCn02AIk11
hSIhfr3pfUVlODXiVTTyAdSreLmHdvBctSgo9RirqYAt8NpgXteQ7k9cNE8xxBz7
Xyf81kStGESK59GdCmdUyCFRAjh9WLnLmqFEVnMA5DQSxwnnOF38gOtnX+1BmH30
F9KX1C9TgbgY+iJX+QsfQPV+/4+KI2qj/mvV80tY5qBqLDmiR9AR8TySo0g4Uah9
1DcNJn8SO0LS/59RXcH4N/7AMEoT1CEAulwMEPQ8cGa3T40uZhS9l6icT153pi5a
wyQeWK6qUp+0fnLCkct+H6ri3tlKQJS99tUSNWYl6c/qNXlcaiyu5Ca3K20w5Ebu
7hngt7M8axqnRSlD28Cyow8Va3aXmcc/9Db/n5gGb59kNMWbGabi8gyGvpjYVRB6
E0DjdvXVFy4nVrF/LgmYhtOLdkSr+VjOGm50aKr0GHDneLR3PkP2cMp10/9fDlv5
+iGFOxNMd/VL0/Nm2KNajEyvSEZwrFtLRZgWSyYEzM3HDxMBtrkqnB98XIDTLAOX
4lRhw7pfd1dx3srjiDSSmRUxvQ0lvLm1lJspFgQ3DpZgAF1fSH17zCtVNqZH/FVM
fK5gew0MEg9ZsN4y3s0OY3wHP+j+T4Q1RFlQ1qBiWNNP+ZWx9E1XLzboSi7/lLbA
bX4n1IOf1RepKPgFMRMRrLve4RFOzcJziH4W+LWyq5xMmnG3Vv/wDG2wcvROtppE
C6SzqeN7ArCgMYkxZlVWcU56tTmSwMkYw1bnbUAgZBaRTmnZiQ0JquaM+F9DW/mg
NKTbEYc+9wFrRw9g3H6d+rEEwm3O5MwUWkVloeJodpO8uPSeTC6Vm4YnsUbX0DYH
GzTHhUCuz0u1nbB+gB8PVLHAp88ISiYw8DWfpCAw2/B8PdzQ69cBoAxlDYmeoqE3
W0tEJ38pJJOSf4yMQeutCuU0zVPAcyBin4cY5XILs59GTk0JMrBGAktY5x7bWNUK
k57avRIPB26htEi1Bnlv6f35MSaKxAyGqZWUtuDWhT/8w546ulVKgYFtt46tXe4B
9qim8zhPUNcI4+Z+tz8vTn+X68Jz9azf5EKYo6WYEu2XOjV4+F9RE803r3te7kPK
WksTa04Z4mT3jLwUDzn0ZY6w8Z8+xWf2rVeYmG7AAK6eJXOYNR+05DPoA0IqAb3p
iI+QluiQZLK0VWOXf/WUAYGuwr4gCR23TOOyQ+MmMgxJLdwEff3Z1rz37FxuRi6f
zpNFLxk9Me3RF4F6Z+e6difunxEuJnRKmD1K6i0iVe2HtbzYzpORLaBr59f/ZGgO
SPivaPopsB3tTp9EH0sbgC1Fk9wWIgDxbMzOtmLUcmHGqBnhhEvzs8n3gPkh+NO4
tiL2ERD3aFsVR3xUZxBvezciYvFPCwTATKsMt3TOmTY9Wi2bAJbq5QAdrG9tTb5W
UxYqAYAJsoloQW2RxC5T/ahlehAoLw+b2j16+gI/zqoUkMXS49VwSNF9tTuTyrsv
JmOZaHkqA55/6Q61O7qECgvZOzOKJ6SGzrXkN0QtqexTu7sU2/ZMXuFWCYVEaKv0
i93rT3bfqw0s0DUbGqA9dNjyO3Z9brMV4TYHyPUygg7iiSpwWd6F/Je+fj0ftGw1
nP7fEmawn43Cs7oQpcCLExlgEFMciyu/0hF2L7NMbQSX6QCSv8jq8exNNoja9/oX
5sdD/hyDtu+LrNCxFLFZdhM5+C4LIUoYSKSZvlUnxB0J5OJfKO9T5yn3NXdCQX8F
T3+BBdmFpXCkjsniDmTz1BuufzK+frU7Wfi+aOsNWCBJYOhZg489tdlLBvU7gm8x
E5nD83htgYlxn1sZzgneW5JTOvSh0Ey04gO9Z5TqYrzgflZnrq+BP0ESh7K4iM7Z
uV2H965pLk9Ob0kILQ+70lttnmx8YsudgP5KFBd2HUnTZV7/yP5g0CCPQb0TcWNA
Je43qGWPcD6Uu9Dofqd5wn+QKAlgU9PCODLxbO2+aSmAoXTTK8c5v1Hde2h/Mxd5
TDSkpT6XwSfRbFfRIYR+jLUXKA2b6Rs2bWjQG2OGgMBIhtuZNqFisw8VqQqNBPhl
W2c2pQ7BmkFmvuCyKCxMsedhj7TG+UFjGSV0XIwsaUb5eykL4D/cSAo984rlLXsB
DSgnF1XryA6yrSvAMgzvVZ/CADibI54ZmnZo2HWRMk+ZufV2m7DWfQlBga1G7KTl
Bf/qaIGS6d7gWIKtDY6tSOpaXILjJ9pXcE3CXrEZ3FB6kdGdq2VKwcel56lNEXI8
1f/mKQg7MvmidBiWGrHEZG9m5SZsHIMDq5TWJnoGMDdsAnjfYaP9sJQvUkBhuJ+G
8DqBXdvQrlNRZJYrR2JD1ZyqtmPRII2XGuLx5bzt3gqZ0/bI62jZyhSKGHaNX2aZ
QkDp+FFk2uBarEQUHJOJ4EIUce5bxiIvNCR6r/5RUJ+Puvh24fEMHh2eX5sK0jnR
FC/82N24cqZLhScL/q3spYtypUd+j9Ng2m3VRMemQnCgcuHtReN61yKwAApY8Sjy
oxWPswi4kPlruXW1wRcOH9iQSV4N/L85Tt/4X4FGF4Cl33Y628mKdsDtIH++P0RZ
3/BlAni3WTj7c2IwxyRm8UfbuoYC8BZsZ9JfoVWeF4kPEaIYpc/VPffggTB2qojC
Kdq29XCfMBmwr/dkKnucpeaafthS4NhX/PVC2j/S/IuqCijhxvliZDxPv7yiGp6B
eqx6nFJJGtVxVxVl6tdcdo+kiy+es1WJj+1/mb1cj7gr+vqA9aRS3i6M2wehBW6I
Hf14fH1qoqnFx5HhrP5kEs9TUJ9FD9A7PEjNSc9HcMh6o46GonwcxQyX0WtoJZX4
imMoEQBkYpHTuhwMrW79wBhlwD4J9qb3ZfjI4mYhUFTFcujsGuv0pbyDUb9Dbl0z
mz2skaKhhg4KS8FszJlkjFxXJdk6mNCfTfEam3QeHiFoZnWSArmP3fikWo9n63dv
EuL/UOgoyrAF/bwQocUr4SmnawzQJOARbOA5Vt0RCjRY6cfMd74Je4ydhxn6zIgE
GxHzSVp8tVmiuXETZuHhoHgMecA5DLOymuqgsYI21Px1a+gYDoU9B3rcww4KcNph
m8EHrtL0WSQi07BTekW/cBcLFOZ8fQ5z0QT/SaBw4hEeb89evVTlrIEWJb4QLbOR
475qbYiJw5z7zApiaGKMBEoN24qvGp1cFLjbQsDqqBSRWryRH8U+xiUb0ZgZy/9N
I4oQWOvQ0TL2ia4U7kDBz2zFNf23o+ZQx2PnLWT0rV0VK5S0d2p36lgWzPO2H40P
jRZcIRKonzbHDU7pJEXfsAy46Y6YDerWjtkfWrQJVMxnpz/7yd/+iyxX99yKtLlf
+x3lb8gIsX9HBnaritDTPwuHZQIm00fqZE2Yn3zgF2fPlvVdGNCe9SsCMmEBvEjL
n7FuDZ4a3ntzBBY8qfYfT/d2e9y1ai3fNCrryEMaDHkTCICJpk4P7P2hQORnQtsF
sRIGRf7k5UuirJ0CuTiRSCnFuATbF9zubNMjl/9YS/HJcPFl5nxA/m/y2Kmv8+9c
W5H3nxdgcJsWmOZiyyXfP1kKOSDxW//m+SEcipw25xpDu2OmIDC7MqwDyZYLBWBj
mfDtWT0NQ7FsxYo0ALnnrSZSqFGzqNgQrPhR5N5HUtv5WzumbX+Q148nX6Evt6T/
S6/0rs/1mo4WNqAwNSrsFQvmiZx+/WZ4qZ51Js4kfEzG9j/N7k4CtOdoHG9dgTIv
XdaQiIsw/Vz99ODL1gqUwt7KITf6KpkPJd4f321rVCXEMVVX8nWBezsgh0kGQ4O0
+z8bxFy9k7XQBlcK2SYa1gXG4sS6rAi3f3jnriCksT5UWZgytDdAxnGDuS3FJxnF
IP52NjlcUmqBUI/B/1RygGXQRt/WzvIVLxNFxHw6psd+uH0FmQEvE3ZLR30mW4VV
0NrPBOfYrxHxnY/hNCHrztagMgGNQhwxf0X9jMHaoTJyuakem9ivQ6Ohy7WzX5BA
//QpukYobpj+qTxMXCFzUvougTc9RxCvan5TQ7Vo+6Upn8lrtMLRpgw4B6W8PHo7
r8gyv5kkqp8/hAv02b3gUvKXGM1fwJWHE0D/CbujK46UV94WPpdHK8dDdr+qA2p/
S50x97hEwZh412kA/QHomthE7oO6OKyL0Oq77uyAS6IKSPqlhHXa9njotLmBVsDx
12wN1nVwKxIy5gqnXaITOabv++VemYmwa5pW7qXIBNSlBpjnMebJCuS/2lIvAJaK
YilB+/J0whTFsmJOX7pRIqe4V2jK0a9QxIviXkHAu7t/7seEXUoZWIGDcOZMETiA
d4XDTCsK5CePFU0t/83iX33m0ucjvV2W25I5ROVivoZ8ZUXTNVxOXWkGR2TYuXCZ
Y6t6ZVANR+pW51NPjzpv0YlAZF7G6lyCX84z1T3x90qJrZTTvJCBSHoy3CCXbmX7
8HF0TOl/ECeRj/yX0OjorncBriVCGwlMZrurGSqc1QZXn/PYzYFl9LqXgxkHKK/C
bJzjPHek4a879HEb8+jI9PFzk1gCaQ+/fx7h0PgbD1Rs2fNX8YFjkL4gaqD3X6og
FggzUxFKB4FsRDeCrG8XE73OJeuAhjsQh6/rbByztLXeDKdbrjnOHYIaRtkHn5Cd
n9PB8uHlOLy6MillNK4OMLMzu+epe11FQ3z122Ppj1jMBt0kOlfsmmvJzST9pxD0
v0IOImPSMPYOOs6Bee0uuzYCosUUXjY3WqV7TnlzI9wh2XLtigY3/5ooVZd35PhP
PH27MbnhfknuLtHzihflb8yqFMPW4qVgMhs1HAaRTZopboqyY+xK4Npnx7jKJc9z
ID3evLa2beRg8bsvBkX6xXu7EtfoR/M6Cm4Ah8jMamk5qCuzgf7GRTc8CVAfqwpL
8RVRyh4QTn77ntXuUnxfatxEajjGqQphqmkqVluEoldEpdbDV542tuCkAy7caxof
tX8bphM1b3HaKCgvLekno/lb+f5DpGugOqCxMfZ1DPFuZk6u5CIdhUbD9FFG9CqQ
dfbZH9i6/cjlJ4b6r/4Sq10atsjNOCkzCj+AB0Uy8o6qoLHKjoIfmaBI/A0AgQGW
zWuC8jQpS/PmNbAy2ZtrxXO2f197WkEsOiU/KRJFpR/EOrOTVcMZDDrfVN4QKNXm
eAn8r2KOUVPJflQ2FI+d3bpgb/qPUksEA4XnThZLfEtEtvGIFPQYWSg5hO20Acrv
d5QJrLy/YcZPBTPjfh3ZLvn3M4sJaGkaXZ1kEYljJ58Pr6Ck6Q7DbUtgRR+WWcZa
T8B6QOU254ZR3LbdXDW/DA0tVi7CxCUfoaaVs00iOk7Es75QBByNYQFNTU5hTTg2
PQau8z6HWguPOJ4iQ3IxsANV5sdbPYI+h6gGEk+DqoqGMc+pMiAsWQpXfUczrsBF
HIS6c2pd0DZORP8j8+GV0Px93TeUrnaKPryydQFyCbmjx6ZwT6S7+iitJTCbXq4s
J1CPh2debglyQx+lUh+orwL0/2+b0n0bXT24mML08Sp7pClkgxQq2C/mkZhONbco
1fLsxuC1cKHh9hsf49UtKqi89wTnzWSFZOXX2yyWQ6NZQfuT4KCfXOuRLb4A4Plm
8htcHY1oCreQIyrkAp/yDGFCTTnvfkK/jrZUjlblq+HUZ58BbJk6W7LX8D2juJqM
GjN+ixskvzqEtGq41k34q4O7tZOtwJxqsTlb+2DD1smHa5pAsP3S5JrazEGx1eHw
csCWZQaCUYct+sVLaPKA8qkJdC8RlUWS0EtTmuJrAUviCSeYQ7FA0a9+hz79F596
IPYyApAHchE88RE3GJxlENXc/mQILN6S/0g6jli8RWNMfeRvOwkdbvbiWPOSTEY/
StdqdL5nDEcD9oazlzCuAI5mA60BqErAbXFlQ8T63/IAr8V3B1ijfLVEjSiVIjST
bhJrB7cWXWVmgMARdPl5vMshsw7hQy4jwL6O3h5u4YnpicXxwNHvFsY4GmMvBBiZ
HFlUEx05i465t7DHew/fuAZ5D6a0+y9a0r9h7nTdfgHAaYOlVwNI+UVG5AwRfzh4
bgFRkTbulmOHu+Uv3MjtiI9HbSfrbfqVMftpoIc0cPhFHZ/ZdqIqKxOsgceWAmo6
uGbE/Un1THe+NuouL61tAhuqy7nDi0zsQS2jo0un8YEUGpA8pO813DKg8cYWFUAL
ToEEwuufkLf1IJemhJmBbtO4i3lW8lOG+Aq+2DIPogvAc/MeojFnDH7yLv7igBtJ
Kc1YygA763WE61tmoopc+QfibTDDtA7fgzHxIOKXA/5+k8mPV1Dhr9BL+7ZsVc3O
Y0Z2W9gC/2q5ZhmAm0lDVUP8dViTbi7ZCpNNPKHfsVCoWDTtEpiuTjFYnjE/hXRb
BVrT38gH7sahIVu6IWNmqbRs4ujxjYXY6QiezOl5nfuyf4n/czy5clyaWovo5n9D
nlVsRQdAjK9sFxMEzhmXf+q3/ybHnTZV31EpUUXS8iFHdT8C+gNFsabdkI3arJza
LTncIFJUhGBjdvlE0zyX3FgXb7mxEZScdbOuFMpRC3jnYvxoTXCKTRfL9Oclxcg5
0Or0QO/A6P/kvlGiwwlvdSqi8NfXjjpWZxTNyBtFMtcyWjnfOQW32OR3YRHQR5Y9
e8hi7lsVOk4vr//Hb4PJ9UcgQ17ZcxlA/X+sSYck63VRG9Ivtzgn0MFuMhrejSLT
ZVD1gmiraBrU1Bfndn+IIYKjOqdSjuzfSkJQdXSjnCqgOxKyl7Bpu38jVdVOJR1P
JKPbdXQPKoprg1D2t1cVDeJiXq5+inCQpn5is9JhFpp2vRShKUjM8YQFwiTOD/bs
MpY98sxSq0XobnvleJMl38ILMs9LJq01d5jzqYuVSUJaa0cwwNXvghAbTHKpQxe4
zQu9R5eENZQVwsLVh52cFBHknN2DXiI9w58shy3xvyvqJLpR27sgIhmmkfNiuGUR
644IHr+NExAn6N8pFdwekv3lW0lvR9bqDpVLnMeSmKQoybLYowzY21bj+Q6uONCG
Ic4Qad5t+pzfF5sEL5P/DSyeMMpjJTnun7HCM32cE1Dmpm+gGF4PiAa6pCOLAl/v
9cFLwsdJ27+bBbUILiN8gRUEduovlunjs5zeDrdO44FTTbivsE5sVBvoS+kVGbA+
/ShvMAI9J2FkUmwxlYAAx7dvFfHMq+0GcRJB+xFGCQ1dACtd7SWPcY6uVGV//CHn
CM4l81iLkJC1GfM+GLqZ3Q7bzYhPKGCW9xP3nqkQHuuDa6PUIt3PEkU5hQEKnD8s
pV7/eq3hDp0yAQZVSiSBVqv9eB8PDnOXTNd3G9ZK2sXWBzTlB8x53zXcDC1NUwyN
9+HXWzbXQNA0Cgiparg0g4ws1iSh/OMvTCL0SAg05DURwrkcALXDFUtVKfqRSZQJ
rrXsFGi7IYGzpAWIYZA1ILEoOKjW9dw8+7IVUFq7U1oxEaqm0t9MRS4aGccdOl3x
b52rX4mtmnlEreE+bFVVFpuIRxOlkvd49vB4zekRUVbbPTpW5dJbi3nq888cAy/n
hpB2NuMc6ycDvEBLLs0MaPnzqO6AVQ+vI+527ltnzJfYmMerWU4lWTNmyGRp9D+T
Z7JFO2f6bPkue3UtSzEvQJuhkrm+kOcXxJ/hgIc/Jy9WL1o+SuNj2PYlrqz8+y3D
iViRiQAYiEzTL7T3338kAxgvBASrTplp5CMZnSUiA8RacP0PnFpsYIfnI+lFDFTF
kBRiC43xHZJDPCdVknw/QZ7Eu6vAPKoI6yUjJgh82JnWeXXUov3wRafvJL2L89k+
CUVLGmrOPyaAiPRjtwdSW1WKPJxrNNykhzjlQsVX/004RQ1jI5aB1ELE8xejCMeL
AyeBTg7Fq6PAC4HlBFo1kXrlOMSpCP9CFWdsS05hLM2dMI2+zeO+uTsiGprDUrkV
XJCbW8C4UDXuJ/JlsUoouothiofYkbW191qdhJQW+INrPKKAL2MC38iPLl/qCfQ0
tphw9tDinlJ8q0H1b9fhzLST/SEKv9D6yS9/8EF79p+5WR0W1mQIPiR9qmct/Z/X
g2MgqZKCYtq89Ws4M5FgWfbnOiQOl43HUaOGdTJ+8+q5skNrQmPhYe661PzRomNP
RPWwDXMKTTeJcd7B2HVh/AT1o9laB5FL02JyvUZziHST63UcMQ3+XoFIpZcB+dln
R466cSoi2MkUkIUFADaOWGTzKQ17QfWg3iYrz4aliO/somiEbk5jzJhWwREcka90
5VYjCEXt7cGQa5svlIjx9JV3JXMpvEPC1+Rc6i8xBR5sx6chl4DBffPY7GDVKO9+
NpWUF1WNkjZ4SBzantEjklHc9j4JMblIhrbPf+h49vRvSzcppJ0ifLAEXZhT+JNU
YrZ3U/apGxzouSBjUr02b/rrLxYLNvlpLgnDK6X/p1GnMXqL3LE/5pZnRzLCeo+E
pApnuz1LZGJTqNaN969VaA3j8TKCo+JmlhJUgaqyfqCkSJ5Roi712K8OAYIOClkI
/Ysm2MB3vajBjpGIpsnH4kdoLLItvkAuPvZd5f3czYLs+PNAYPxVyGg3G9HxVjx/
rkr4XvK/49++dRElkJO+4BhfkeadypAba+WgVm70gersu6BbtfUmufJFmWeqKQfS
mLGX73qgtGw8SgG44sILJzpfEALAqeyU5AF8lDGVzoSaf5yoswBBEHAlvtyZrBfa
UY6ZCXn848BKu5rtuItgh0uemi1+kUzpeAueJ0mEuszyIbMMBSwKdCmRdZKEhc0j
+/aXMZCoYtsK3/3dy8W+MmsAUw9xQVEsJe/dGxhcOJ6iGYWPnHQR/4lQ8rVzImNg
sC84vwBufQJMTcDJped0rs2pQKZd6oNc//QlpyCPOWlUF1nMV+lFYPO5ATezphxI
/BC3MvDUsxmMDDocqaZDIykLCg1eBUQ7hX2WV/JzEZSMOTocx1Of+VaRcgatq7EU
Z3zXTQ/JYnLC1EdLoPE+SPhsBV0GPWPFZlyJFSFB10S9G2rK8ythbCJvGcnjjScA
ij3Cfqb1pIl6dOIegbOeDqIDXpEu6B2R5uV61NlXgmDDIU9QnRbdpMEzF1N4jbM2
yGvUWRvfhO/faCj+NA4HbsK9J3y+odyIu+1ZBZrllfwsKxg6ZQ+W8Ia88frK+Css
FAvwqh6KGD7IUmCuL9be1x7nAMK3WlUSNDsRIJjx7hlE4ewXE8QqV7mQKm1Q68g7
V0tfcxu7Qe5Nsku7eVYug7+EmqyOc5IsIUH4tUiz4AKjKTyO2L8jvig2mw9gjb/j
Vi7ZKk6x84xBJnM4zvdUIm3KqGMRLr10IPVsyC3VNlsCKFOuEscDgNIXPx6+9JiX
S3yHor9Qhu8HveMIyUdcMiOfXIq1/VhrX+8mq4QAUmOGxW59Eq144ks/K3xOalqs
3uhZQ/mIdDHuNe+fo4DxU9W7sCxYusy1t5dfb45Ztq65ocLFu8ylSy5xKjELTwLC
v3NbQtGvyNiZgfq/NkK3uhqsRcB4UM7iY+2mB7EuTz/6BTOGdRDw8HnjUI9N7FER
ky5MfncPb8U3oTKVgpSM4tZRmGshwLtBYo7Nq+FtjlvjS9nWduwSJ5Z8TadYcKuc
C3JhTo3O6vyUST6GVmd/oBBn0C6t7/ZVAkYMSQ8SBL5WGhJ3jjNeMzL2MCm2bWU9
0u0G87P2jYOda+2z+lFR10s3IGUXqFTNwu0bw/sqtvGUfzSaBxHzckvIY5zXVEpO
0aXaR9B9R4da81vxF3fbOCDjpOHDwQTUYMhpI1xbwbVraFpJ9eyw0qJf2K1hwHXJ
8n7I0A/EuqOKQAzEarhiMTy7CW0qKRl2E9X3UDm2U4wgm9n8b4oETJX5Kx/wGsGq
aqJGKBXa8P78b3xy8eZcy4xNTEOe1uObOtA293QbRIvFkK4CUfJkOy3j0Ww5+TBv
T6bMklAAbLcELdj4kNZZRAW4R9msjHpaHxkkZbxFxgP7XTyl4TaZFOgI//7Y2HGa
ihHAkKLChv/OjhWEI4ngywl7LtAd1Fu5sR79GXhHUFSCR6VhDJohHtAizZM5FV2Y
YkmzxiNThuTYbLG2yMsfl+/m4maQc/hyoLsD/m8Hex7QpDcWVRdbkjHskeYw1nn6
bhubXEaPiD8wgC+u2fQSxYapI7Oiku2sA5PYjRMdYjEa1Uq2wNT3cKn4L/vm6tMA
QdbZpuKxRZKxFuB/GXCiuX6yEobYRIvSXh2/84QvWGKJlMfnDNCBPoV1/SyMdEn7
mmzPCT4rsckCLnAoQWVLlHRUxQX7vIQ08LxGMumUqG8YLGvOUlLH3+0lsvlrT17H
gcJy/R1reb2PQVGOardBJB0Rjz8FXWNm8GxFdAPgxqw9GM9xfvNTnIF20roHSJOT
W+zo+7EXPD9jZv16YaQg9uCUEH4smZaLze+ZvncjWf+ajmusIxPEA3+TG02983Yz
fzUUdGBvYYQvPJIn+AI3ddOKZJ5EZzPxP8Oz8bmjkS4r7+M5TKjrjeUUAlgsRGcy
a1fVVE93WCHVDETK5ToXpMJnz3xwOSkzEn5Cin32BS2g03jMqkMSo5zfYyZyzDn+
LT8OESo39nTANG274JcS6riBS8QuDv63C7Lmv/jhbD3J1NK38c4gt7ZJLaRlDIeW
adnjTZaEi1Ll9yPT9FcKR6NzC3bU3JdBRKaKUQbvoY747mDOmHLbVLVUsk+ciTjP
OwXYBZZ2uKxcyKc9l+KAxbgseIoipExxLrc0phjy0EHh5Nj+uVBzzKqNDb7Sw7sE
LEOUzbhVIh0oh6EK7H94GNFih2bpnpPplRjqwty8f5wauDjHXogVlNAkUyRZQf1d
Xm8fuO3qh/hE0WKQONGO7qnqUKvMhvabHjLXCwXaZWDSw0+E8xHGS+JulUXRMTix
e2KAZ+u8yT6rxok7QKFlnFF4jaehNqblQh6fGHbdnT66IURxmSRENaExbi3uPg+d
NRO/TO5ZV/Q+BltpkQdI1kuZKaDatPQow8Lb5F2sgRezp5SVVmHv8NCQVKPEyXi0
ntwZngsXSTuIsGrccslx+8cJhBDN3fKMUOuNWfJD9mSqaycHjlKfe8mLRQNCLZMA
OO50MBTZbd/FG0cCxuDDw4DyDZZU+waX+lTaO2wk+9qdw+BOmu2sK+SG1/iGTI/6
sAvQGeSg14bZuPGTQ3Du7ScNpy7R59FsZR/qrYuUln5635CB7Cr5TaF1Mk6kIlbf
Ua/eDw9IuaxpHiS4mA2sFcXnmkktTp/vnPJasKNeI/4nvkvJRKKAOO2l1PL7tSVR
fVsNjCdFCmKIA1kPt1CO8ZOswdJ+ZRjFaefCRKz7HRlWxqF95EK9Lpt0S4cLPCep
rnDMTmK8C7akgH6MggTRJTkomFA9np/FdeMIAWjx/3XjkTaaDWcNU0fhKO65wyV9
NDhEKyDTEDBqFiWPBa1ent8JJViiFgunI2WgBdqOI/YbmfbCnu2AhzDX01gZwMWX
Imwa3bOD74kE9OkxNQZ0HetxfLSkYqoLliRPFE4/tY5RQghHJNQGPqh94U+OLhL+
G23sKbz83P6u6/o/M+uoOalv+GQgL0hhc0sEcB7KoF+Ayx7UQQH36JYyi+yD0Nq4
VzBkM9iuhCUg08vG2SVVlcO+ryrArmBVq9yw9fmFkWT8YDhVUYaUhzcGoDixl1Rj
woq90Rpes7BfyuakOwa7vsrJrm6fWQZyYcu80CcbQ1qabPmIZoABqrY+9i8fk5Y1
wi+F0LhgyS21QSzM84O47YJLbEYUr6FLbyyLFqP9umj7J71NYYuQPX3fW4j5KREu
TjM95RR8+aJftsta8Py0Uj6BUgGYlxzRt0zmqDIgzchV9e1iFDYLihD+m/mQf4bt
9LSPsVVQ3gC73V3QaNei7bptj3KAUrP3XbEew95PisrmO0p+iLDi4bX+WlftKLlO
aSrVgGmtG1Zhu7l0NN4jrOH56jlkj0zbSPDjYZSpVBSs+Y8vEzmph8UeJ3i4TFgi
3WWgHTs9iAW37qFNeVLf9LZx2nn2W9HXBd4fmImrSmGiqGwzV0FDbBGJScWFB0ua
fOmd8Mkpc5H5vp9VfDU61zEHBxU8+EwfJKQW9XMj35f33lUKSmOlpx1Pe9p9qBLw
C/25ed2pe/WhVgaI27wWEu2cDCzIVfK2bZsgZfhORa4sB5aBRBe3+jVJdjyz8rej
HDeBwFWHm7jwBmVEWQFda/Y/kvvyRM9Zpd17x3CvCjSb3a8NoL3U6LbvTHlFCoY3
WTn7tQ66fAZndp/zJMxvmBn9WNxuLP3CwPP6Tno9KNEYUaxwococNKHBUg/sxKzw
e8t03A1DckVw3RI3zCpuZ+SOjisHAmyTUv01HCQrlLDRJbY75OxUFQeUETyekCs4
jsVsZzYqweM/tSYFkScsCkm4Bfg7XfGBbDyU1X9UqiicVmJjcv7pDGIrPxt38LHJ
2mo/tcq7ijPJ3KsB+VwVyX0OW/T8vqVMurk5cQpzKQ8A8lmZCysb0Hp46YYVIkVV
J80YF4frJ8dYDdIeOopHlsx0+uvQEq+2q9Du5MXXlHWMtYZ3E4JJoBwtBeTjuxvd
swlEbmQ2PRZsXq7+4qANlMrT4ioPp9Rt4V0jGawbYOMLnk0Xq2WOs5xhItvNNr05
ajQAXSTXsbHrpMUNpt7fbxJcoBj/KpGRkHBH0zFIioiUm3kp2JJn86tc1Tqwpswe
Okg6/x/J8Ot4e9CJE8f7NuXcJU034N1oejU3lBHEtSO9rKZCBhjNzTRgjPT3g07T
C5iiikx7nLfHF87V32+kl/x6NQu9dSJBfscTrOvhciBy9fPb5hVdpvQso3jZiIxo
bCJajKttfMiLuDP+J3k3lL6ONlSH5vFCYlGa9VYlGDkxVw0hLtMsmJknTR8r2dXp
vHrLDn1+ryIIbIepGgeN+JNq/ZgYEETFX5892uCt5Z8xDmdMxGC7jtgj93X6UAcV
ZTI4Y+AcxWrYOYzYxThGxIgeNrddOiUikHRwJhsAnoWG5jfLPRtd9CLtpGeNOk33
FVydEoZbCkoLcKmTnX/5LaW/x9qispFy7NLDdC1iXyuvtmBe1LUK1zyaYJL4ars3
Pcvj8dzuj4bhA7D3hzb9h6tPq+D12jJBzc7HGPzjjpMbQTHYDQ+pWIyh9bPyI/lW
j0dfoielcMNamUjf6OSNMy7uEOAzEEVl6wcb8DAsngOU5lhQJvysAV982Kb0qeDi
rOWA+PYAXePKhG5U25TUZicHKTQu69C7oegjtvSlVfC1A4k4OgYXQYm2s4RtGifT
9tvqID/0DpJmiuN2QEn4pTnhYCrFm6/g29eZ6ydcf7DjkJKMBKknqw37YjpAWF3O
e5wARlfRxOIj5QxSlsov3oB3zTLNjC4BQk8MvaC+kdgwB5w+D2iYYoFrE7wAHhfY
B7x7L8l2pFNHU+KG52UIJ1YoeD/ivJLRz5KsJmIYznIb0YNvqV/MgljgUT90Cn/W
1sE3O58NbmCdaxAoSx1lTFtJdOe7d3oXqp5KG0O1lZA8qeLAYpMJ3CZRXaXcqG0Y
XjRjIb3jDWyIg26Fa4/8WhSpacE6gE38NmHnFS7cH3tEBpcIfr7xTYYFSk6vcVjb
NqZCBMka1X+xdOrgrCzkNlSrS3ZCKK4QVz8QldiQT4MRQcJBSPaq0ish2G0tG06f
PMC93QYqlmaIjwKEyiJwm5ehsWQzM7+GvcmJi3umPWBhaP8pGPkRElxFECejEttU
GTwbqXulrCObZov2xgREeJkc304ZgsHkXabRMn3vTtKTs8Nnm+vnPTgKQu5jBSRA
MtAA/KcljYu3rUKBOXl9kt0cKeSsfLC5awJozuOfipuiQelGh0SwbUrghVvQT+ut
mlxrKOBWIApMgU7MY571opj4/3tEQu4Bo7dT571eAHZ6ChT2T7qN5vXbeT10HOCK
8gXvXNmSErPCyNI4BUBpG0grPpQo8DUiRU3PebxrdfD3j8oYfnoDxcpx7aelrJNx
JLc5JD1ARgt/rvFTq3LPk5QWpBs4xMqaBDBfeSJVzbVJ0BBKzMeKXupdxbnXxq+k
tx1at61ad5VPGHSt9zXeRzjaIqNm2UH/B0XEm1MpiTWA5bSfJymMk120LvrUPSbx
i9H7lFAuQ/aE690MTSBkNJ2zT34KgS98f9VgseLn4bzXERkPk5q8BJpbnxn3Lq5u
8jZeryrAkIFhvOUq40gSUL58l+mpNzXOjUXiyK3fFKb1ExN4amd+PM3yDnIjzdWD
ZGjMCjSQEPvGk/t4Kg3MA5NrgYlsRMkybwqLPnAKdgXjNJNZ+ZbK9OU/QhoEkf96
zPkGxPFrNhLwnenGjGdGT/f3/aNUnkkbX5VuVLv8ma+SuVvTbEWCjhyV5Af8U/AS
BvmazFYH+n3RUiPq8cKiPIW/R6sfnBTiL56oekiJoJKTgV4SGWsI1TBaDavLKlAg
VGr3ev9k55XT6bQRBmTy6Srl3PYElijaskJfhcAfxRn5c4ObXjN+9yye2krJ/5mC
AjQG8PmzmA42b5PaKXl+X5M9jHkQK58FHHGQcN/0Vl+asFd3WI0aS3sBhGKR1qR6
gFOkaZc+qSkfG+qB1KJCbBiTYEfjllEH6C7WUmPloi2Rua/lfPkw9cXWQzea7sXV
OgZ1yz5IA7YMJehhUTXphkeNfe4MZJjDLgFFYbT8HPVhlCURM6Sbbj+89DtYfJ1B
64rc8ZZFQhxBUMfjrfAVEnfVyA6OL0e9kh127RdVaRjlaWqhyZYcOwAoDYCrtL8T
t6Dx6e5Fei8E5mOEnNHDPG0R8JAB3wuo+BNMsgZJJ3ElUwIUTWZg5Ayu0jyB+iLK
tsgrRBL1h/djHIPH/1v0cuqGQeyIuW62cMWp9v97/CRLNNpnQL8PUjs8lTov64OW
V89ZidWN8oystLd/lW3dEOR9DYJn8GA5SoBbVp92zeAhzqAsuItV2SCsyffd3BCE
b2r6+7iHIaY8D8Q15Dpv/cheYRbOuJWVEipRKvp2UK0PCvWP3BKaGyFZvyiTXYYo
SlcFvp291E0mllaZPjNES+ZJdbmaUrMZ1lPGg63zOpdgXs0XOFLtfxfAXFPBHfvd
2aMsegfYgn1Yxwj8hPt3vcnizCnpDQ6GspgAXUPr1RNZSlSxT+fhMoiHQmWzCrdE
vBLvVXeRkAQCN54BAXn07Cr1DzDK9jizDZUWk22TW7XVVKfdv+JcyqEgOeXFds8T
jgK9hiEhGtF9pst66FgC0x0g3hS+rB7zOYBW3ueblm7S3QVuT/L4PFMaLHvVJFB1
YdxEDVUQa4GunYcUpLo0JJWHICnlGIVvrglcm8lDqbYCWRGqbwGU3BbH46/mDdsG
zA1QLHXGb47kZdSG1PfZcs5Y+9BPZzAId131EF2vyabwyn1qyU63f8AO/8/SZFfb
kNkEmcX/9pe5gvjKXZnd9rvAB7rNGWeH6fqWFvSjWvPZoLhyyT5uRqhHRFaEFX6j
oJBeGXJyLSpv4+Y2S3WFxCTdeyzNeAJDW6hKoxILTmI6wCkdacQz6p7dRkNaYobN
L1bZex6g+axgB+3UJova1ikN9TO6Y9fLsI2GNzRpHt1E6oxw7Y36affmzckxjIAO
/YwbPgRxqSU+0FGiP1gy+TI6b8y91Q3X1wUcR/2ZL86K+WHf52imOJMm2ZXJ80cO
kcaI5To2vvXE0r+oFVo+HRf91hfciHPlIjjYuQG2gswGqf9HhuawWekql4AKK8KM
8HHv4oPQOLm25Qi8j1FFl/qeDa3YAeYFGlOvNHjUBo0xqcVhywzwXvbzKae1RS7+
vINSPRvzZGBRhZJk6UC7JUfY9Rc3141aMhqil/IDWZjtnRt1XL7sFsb3yqgy3re3
NGh6TsVdjfUehkZb8iwIoKoWKOdgCL4+h0oBtRkWUUv34+IAa2ovdyNEahTGAcEw
LhtBv9fBB4uF/7jNGA595WNRp65YUDLYVs8tV0BzKv39568eH+/A0DU1nSpAhPeD
aKXx+sjXCKp3Yn535x8+0KmCqFlgL8RGvFGVCIXL4VpISf0LunxZcFjx9igxlyhh
AgdeWfCoJUXufS+GQUUV23xjqnrnLDNfy5lfSogTkD7uaGBulA1I6jAGVVfdtxGV
fRmEOdq9GUslKoNRzp1epRd6Ot0cZvE0d0gsE/IMjxz37y73QbvgL44K+aTFnywa
kvpRzHDNHId4DQJTLnNicYOT5d3W/9cyZDAARPTwoc2YkEbB3ekrA94wwa7kMP0C
O9RruOhNPwoUXSzeQffjJzxrRbwJ6c3zBEDAekdMJZiC7VlWUEegwoEgGSaMri6p
EKBrdayjFioY5USKjHMnb+g0v1Xij2gFpMSLpnib16CHQQxM3nufG4cSdnnbRG5w
+CnvvV/hGOnE9eUD6hJ91ArBYvne61n8ZtFniz0jfXxs4U02SY7Dy3fAkhKxXsAk
uq7GI0Ge8BkyAFxgG94l72NNOOHPMA1kiNc1/GD5+M0Fit8BsOJX2YPDNDcnG0Qf
/pwz5IfpohtJk9KeqZLlt+Oirsc8dB1TqBJXkeZRHMYst3pkPmXRDA3EAR4lhCZw
k31o+kbZ5s8Cku0w8mRWyfhzWUcmo2zUag3S+eLwhpED+J3iRe+ywyWmsK0Ukq/i
V+WBkyhao/0ccqiqUErE3tcb/qw1cf/RM4BsSOAHSDm6gtfIPRPz8rYBqud3znhe
3XFfv/rKpNJHMl7NFt27d4dp9d8Uklpt+oYXBDwqeNsEQXhUGN/hgC6p2qma0iWQ
AQK249HlVRVDi4Dvz+UQ/+yEQpXGTTFfocLNaQQX9T9HBRcs0fvufqgrYZR1KSuQ
e4E76TQ2vkk9LtEmjZURBnYz0iI+EN/LuhrWlNTe6vpN+Siq5iURiY+2EbpIdLIB
/Zz33fTsWzR5rtErObGQeHkV4ZPc5nRXuD4InjicfpLLBHBQAEYG4SrvjPbt2+Am
or81hEApQnLTAdMEQjE20XYSQasgLovOnrDWGehNivTcRrJNQAJQlxMkyog4GRUJ
PaEdf2l3pNG6fwVWnuJ1Bmrkx1+/M/bETS9VcRzPIYo1EFOLGetrVVCRnRKORtnb
vO9lXly8/e/0Mzf6y/TK7AAFzVLfP05xm5FeKhIkLCH5EvHM8q186uAdmXvxWX8+
wiHvK0Fh2UxEqXPifNCLOyG+SO8XJdVGHpJPYfsOv/MXUbqxVPGlO7so2c75D0y2
4DbpqLqS/Sd4iFbtLdr7h8cR+yN/4ULjMgZjtBodh1O6ImxH5elmEdMek1OeekVS
KybV//gihUHMlWz4Bce7mQS9OD1uMPSzZ6xlch22IvSFYWchEm/Pcj3AV7jFbFLJ
s6i3LCHRLahBWlrzrPNv/w==
`pragma protect end_protected
