// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WQgjchKpxU6AOVskJI7uoHxJW3qSCFjy01/btKPg2UdqKKdCxNpeKLG6p5yqefHG
0CVFNzrj5yDasmyNIHOlSxxpp5YICcMqIvzrCUgXnuBvCyvJmRKNljCBmN8eYujx
e4skyOpxGgRifGxRjx7Y/xRAc67+pyTl1xMuc8S/oB8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 183296)
5RLDqqO3Ra+iymDNMgJwwdVvTigoU5cqZChd31pDt3jXi/nQ1rt3tcNhoALZd35q
GudGZSA+JhM8MXlEsgdXHpmPjAR0vurcMIYh9Txp/E6YDpNux8KlR6nm5NW1GjCy
1WA2eEHZ068Z54jRrdYdToyRIX3o/7NaKVomvwDZGS5VBRA5NcIDauOeWCZK1lXI
AyVR9MAKj2ib5/73/mbu56HJn5VFArvqf0nTcy6Soh+U9BV5PVSZdI8yXOezDy2R
EH/LVxvkxKD7FxCXEHJrkQI3xbsid3m65g65YHA/N3G71EvqnPmgNFFnBWJHJiBU
AECwgmVGsn2mvSTBjzFtpj6vAL66y4iYqWPoj1sAe+e6MEmiQSRSg2HlHMBJDbVm
8AJP9TzO9y+nPFg2ibX9u+J/2/TGWABkC0Iljp9sfF5ZIaNMnoJRiVvVg4QM6ABb
1XBfQgL04EZyxZPv9WIDx3Ry5aZMlWMHG32VoaiG8jG532n1pUfMZMW7trLBqjQF
eCWd3YcZq1YJ6gmtuQIkB4Q+ssK2rk/HnKVnznydiyV7ivSjZiUZTYqAK9yH5UKR
50+qvsljbi50BhbFzXa/u1/SoiPIF6ELckYE5uCqY0YuNDMkpqw/5kuDNXdJPf+t
xb6rBkoFmDDS4600awrWDUJPXjvJLU9f0vIqRX9S4kw+tP/CxRuYUTrGGBG6wzky
p7EJh4DW8qBxFLlRFTHE/RfzY5W5GTw8BzZFjLal9nWeUZS/uEZ8NcJRlgy7ADed
IyB7haPo9tn87SELRozkJ7sYLERH06Mknf8fzJ9Vstz3tQVMkDSdpav8B7qsLEt4
DLMvf81wVtd98MBovnuKKQ7ptnerCxVWfUy6nSVQ9XRvTS8KHmoHswFBjOvKpg+R
gfVgFCHcJxMDawwv+5mFcEV/Yy/2S4wFUoqg4ea9TRyIO2n8iH6xrwnIuULmMk4O
ZD9EAG3WTv49bOvwN6gLGjgJWTtWngdqfj4YS+0iDBwWhIjWpUvd0gybYF/65O73
xCtINEiGUwN6BsWw7s4TutHgYE1/SQ9A/5HG3sgJdsU5kZyjanzkyxlU9LGrafMQ
Q4zTUi2hjIqfU9tQt9k59A8o+3C3ecAeDVbVI8QTChA3dKLiYHE9JHJkNg745FZY
87LT3c0heRYl0XyHj/QbPXgp0sI7THOPgF3zuSzY+XNbyfSmTaPiRZVYiHBAs1xB
uKJVVbdm4IicXbEvB9BuapxY+fY1ayfmw1Uzt23Dzyx4Bzrvfn+asSVo29H60V0c
lmqNLNo9KT7xgzcHuVkwAx9VewDDxu0FLdsgW4qWJKTM+s1XKYJ127l8D3/CCb6+
VuPDKUnOfpufMSpGpvngEb7OBnXfclZNRZeGTH+Uqmq2j3uzBL4xc1GamhZKfIc0
PP2TDjKwbmyxu49YnPHhz7mDqV7bB++bdlknFBlguGMzOU5/lgpsFsblOBJlXbzF
VwpHTVnJTSpOshAQgEom5u21SOXpDxwFubWpgfqotSXLgUP2vAtSNrfZrURlxGJt
EtAgmjFzGKRiRVl75LClTMCt+3S2ecsyX8v6Aj1PKUSpNbsJSmFrcbzO3reoLJQt
NY+l4+Jm2xW71IULHkwO5HE9N4WMFO7mlwEjTxG6pKn2ociUT+IJXbkdrytK39qX
d5K/qxRl/l/62OZ4yESPE0EkYVqpYbmNE9Sley1+NkKbxTwJoPxxRvHuoeP8mNFy
fiwN0LXvk5Bw5hM1ldLIE2157ivCP0FXjTLqkbUt03DH+3h0N2pb8GDcA/kZL+oA
+Ngb3dHaQaPRhM0zlxMxg+W5p/oxXyF0iKzlu3xNB/BIK07sYQ4X0eyQspZfrekA
xSJPuh7ELZ4dvag4gKINQPpY/fL431pP/uyxIYpJt3rd1qED3jgheo56+7KoYMNH
U4CtP6Xfhu+mHNdqR9oAPW5T73/p3RXEYZHuJrHxESPZUfajWOLaTpTZzid067EX
MCKdJ2Q3y+wvFUwXlF0yo1zjBft/vuv+REMtyWJd8wyg6Ua9Vwiu8HcPGrsBTubO
kvlKbDwVrJbJPYUYAR8vMtoypaWzMic3Qa+Euo6RAGw8g+9CZ8Fdj84k2BN0Ojp4
ZaG142D3+nLlLWu07Q/7F3TRVxS7ewl6MwjM+8Tuhm5ItyyG/cTP1a8TUsdM4Yvw
NoNmqX38hs8paoUU4deLG2QOBN9EvnKpjb+HG/odDCu6ifqVtJiQHgKds5pLJkgE
3dP2o0a0fs0vNGWgnNk4bGnn5EOI19at9ZL0Rx/tQQyUEnV9QFqCvndmiTIrmhhf
mOh5fH1zzshOviUuIIMuLICBW7wbgg1ifRq72/n5iJ6ULrdvHtZFRaA50Fa17vL2
Utu1EeyAoo0ZJcy0yDNjDet+pVp4MCrAusEXuc5IcyrgYelv1e8PrPJ2AmpIKoVN
FnvFbQH7Np9ys878vuDBX00qKmqJwyTQG9EdpdnrzHQuIwV35ZIjZzbz7EuyPDwD
Qi3ogaphUPTVLUx0D6NoD3WnplAZAQgUmRkUVNIVn37EAfJYfTSluJJHxJhwqWrZ
yqTJ5LYSIdbcvoR97aEl5u60H8KMwmZORG8+JLDRbkaHhr8ggqg2sSAjWMtyNb3L
ac7pTYBCM9ZBWNptp2z1ZwE5bYBv1sZtMsEsfHGxsUOa2kK/ffQiBsdDuSiwYTS3
w1dIUimCwTzu989WRyUI3vYNLG3gU5jAcWl/akl/6BYlvOOjFRjkGIBAXtuc+UoL
dJj3DvmhvAjFTzJU4Ld04sPgrV2JvqRBpZ9o5bgMXetOinP0TMqJLkHkJ++2DsoI
Zk/lZWtZWX1A8RkONdvZOg5DyZiKmS9nOz/RVFijqTfzYK6nvnkGv9aHqF26eZKC
TYmFCelFC6RA1oOSpBi+0MiJnCZ/WYWKCLRU0eLUL9g7ptSOGvtEWAnA++OKnHTV
L2Snxror93oCXz/U2nW2uWPpZuTiTv24bf+3Eru4VfrycMmXsc7EY9bDKV0CwbRt
to2SRLO+gXz7Ix6gGtBwkKp1A3SjAmpDDzDhKy/CF3Bo4rj/UuOjPcou3rEW6APC
TTiWDtyzWQWzSrznO1GQGLGXcUnQs5kgd7Vx5Xwv7I2km6DO+hrAF07LqK6Z25Af
1gDQFDoxDfByntXQrRvHvo4t2oFD4nZtrSuVYlnD3KdR/1+gbfr9N47qrOLGDw5E
OGAJIRrWyHUbqzdr6g2RavuE6mA+nGChifd8UNy9+rxxZCeTCs1asBCFo5KiMCo0
uW7ITbwIDxKEGxLfC6wSfpmFMIZ2ekyewbXXsW+gLY1xXoDD08FTT/PyMAMMQrbB
To6L0FgafVbvkYwNCLagcJrAiFBuk1cvbKi58xN2vVErzsZkX/EoCYej8KsChNRr
2LcV9xzk8+vAURe8xSsjlr4ocGGjxQAFAV7lwQRDfVMufMfB1WtrFQHMg/w0PAmS
7xqUSGHmalOcTVnZk73InfCnhmU5EP0MQhGZZFXzVAR2ITJrQexqNCYkgNsf/A+f
Df2Xhwb3x3H6KdIaglILqN+TjT1f4xEINhnhXwGjJZrvyfifdl4tgy/UMMI2BkTa
ae1yOORcPX4sNvdhO+phfmyQd/DlxKHrIioWVLMvBd+rXY+88eUYgegvP2ihc87+
+klYZbBbvHlINYWlXTlpf3UIw1Y4uZHtdNw6f3fVAFEfIBpX+qOWxkYrLZqJD1/S
tYsroAoao7p0SWKpQM7A3em3zAPWZFi+lvwtE3dAuII/OmlUl4aGrFp3lTZl4Z15
eK71MYsH7pqVDNfiTGYSNv/RaWxFll59tRwJ8uZxYMyTeKXM32EUxeXOh0kfBF3e
SxLuJWO/j+1sbexjWFmU//2T+o5t0yG6S8LeCUoXI6Zr6GyQWWieOWJNWbmGiVl9
qw0zxsiB2rP+kcd6rZdTXG7W654aeJebJL5h3jVmI9Qq02U+GXyeJRhV7BCqvsB7
k2T7z9aNPJDLCtoWMzwkayr2xCeiQ72BRWQS0OW4c6JXdRlGK0949udq0gD0DLQL
nxY2BUnC5EWny9H805czFTideC4v/RhDLg+j2Wzru/EqJlxK8ogM5PU/YSWU4YAC
jxR3h4k+RvPKi6nngcc7p9Y4CO2gqDCwsXqNA5NWvAMH1qcED4UzDSRr5exFs1eI
YTwwj7QZFXixQqZEok09nQognGIVt2imCPG4IDRpwYfVdlFQtYte31vOOtHA8T9b
Yfy/mHNZUxinBfeXw5GDCrsu3V0QPL0V1+IC+ptyosigBveuB4m5PCsk6pfBKseO
ajEGW+mqStO9RCihMDTUAIQxzvxhO5qq5LvTQ5utRhX9X1nvhVmkyNP8k/Bfo3/R
pZIsR5JzmDz7nXQmTe1Ajtov+HAhqVBT3qAMtUS3ZGBisetfRBfmUOSCWa9cQLvr
Bp/9tJ0hYiNWFKA5kMLpfV6kLBmrBO1I7fvDSCCyTb3Vv5nu0+e8zC8+WmEkvozI
4x1uXvwOMTZnfK4NxMxKGITAc3pgDztqnpanilMgxH7z68asWb17+MILcUC2BSRR
21xPrNYM8CZdoJclNs75LN4BjUm+Y+bc8/4w5H4l0CRmQHO/o+WANeJKzR4XS/VV
98NDdnUlIliAPkhaAug63EWRyZuvl7/XDX9hRzCzuS1BnA95aXRDtRZ5W0a0okte
WDS5QWVlji2AFsAev7N0sAorJUcpvl4kXq6D0xzVMpYrEQvyeUh8bYaNCzCRFhF8
ftLXPdddYgOBjtNLYE4DBs41a5vYIK2UWNoimyrs/wogObI/iq2H/ejYOi30yJk1
B3z2tws5kh2TJbU6lW24Di1xSZS1xKah2Dw44KqZlalLNTaAIG8d6wFoJMqoZyAG
E9HSr0xnbgpG8K7OGrnmBssfcFuFp0tlD5fg7RIkh672h2+AVSqPI+65NxzixzMi
kVnKJaBeFnNOPhbO20gNhxyfIf1kjwKMc0YlDZr2CpBNkqMe7dNqlxKr9jYBs7gD
kjgUTkNG4Nt9AI7L+U5pLkxVfrVVPr/FMPyqJ0a2yZUAg31/MYoXxXV6h+V9W06G
SIiSiKnHmYNn7TXdTgOXRmWeOpY1fxoxI+7OlFCl+iH15Zyj/bdBtfLSbY7rbY+l
KYQXohkCvQw8swiDRJtS5Zgg+/OQCNF8bquKTN93mzy0lljia0FN1Ay/e0DOhFQ2
yYNu6IPVvdUKhE/RRyqqYVNBMWxfv4foOeJxJy7DBS2XYTvm6PxPBx/PVURStn3n
t4joK/d1zrxko/5vMNWw9aSBf7gLsXqAgSoRChIEcBIPkcvH7Y7bEzDNbruMCxn3
chXUX1XK1Xwlqu+RDfVjdS23qJCgLfWy8Ag3ibaO1dIPix3Heuo8a/tZm66uAvFb
jHKcGhVkJrd8GJvYxsyh0sRrkDNvUaNiez1ZQEMfPfYkeFc+srqB9uxTmQ+1vJsO
rHYnk3e/ivssWS52YXiq7hrlv5JeAwtgEXRqhSeRtFX2al0HR6j+heInYDp88aEf
PpfEWPPr9CwrSSThu3eUa7WekUbUgDeMLPAjPcDOS8MHdIobhhuVvkwtIfNdeXcO
nFDlPik1GOSurdvFBE8MuKzPo55keo2oNxbxOvVE+uQZNUIBqwSP5fDMH4lNxA4z
3uBQAE16SrVJTZgmOBr8wEFRm9H8vVSPfSQYQQ4ooGZRqe1bZibpu0BVx6U4OD28
7z2stzFEgcjPlo+nAZ5Tx1DJt61Cp5WblxJPoAiiz0Mo+6cISY6C/oWcIoUuirmE
0dUz4zKeFGYuDa0nVCh6KXdmUZhN6fAI+deisg5rkqKoIQTtzW6hPnbBjbRbcD3U
Jd67Nc6k38V6+cidI3ZjNDVrueslIEuSflyWPbtOM15jBLmQWOdP7HeTqBYP1dUX
8vPpUgos+sNSMN+KcAIh99QHt+b3C8BjGqfiontdNqnDfGTALShvGnSWxV/EJ6Ag
CFrc5GLN/Y9w4zjSGi4AU8s34X5giAjmoGXHkhStR7LmvGNMShA6M1OSyJuCYj5H
9ujjkAbXMSQdmf/k8FEtGHHtFFTM78N/r46r5Kpyo8g3ElDUORXS7mdPbjaRL0gx
uh2aPcJTbgElHrROrJ20uSVLMLtTS8xpxSUSvz6bUXu7dxLKDYv0VmilM+/LvXK5
j8ZPltPsz43JlvxmLELxX1+ZFup4pL81EHTp1EkaCvfg6NiTIZkwLL5TUhugZxCW
EeymzgD9umhPVbHlrDbIc4Lkh6YGOsBfjD8IL9Q5K3dLNxW7FVVpXl8Cs1z5D0Hr
INP05ZRPqj6ogvmybmQlhNPYhU5g84/dOYzRFFxE7ERYviQFRfxFC6COW29GsZ8a
ChdiwB21/JfSsA86yuguegk9bwH2M4OpGUpZl8QzQn2Lj+lavq0d/loamuVDOWvx
uCBcYKrlMLm07GMozHc5IpRihcgj1xFi5zA8VZI1Trhd7MoQdXohADBl2QVSmeia
9Pg7RsE8guWpjy1RpBDcB9IN+U7/3HuXz86vfpcPTZs0B7J9Dlvbrs2B5KVQ2QLh
aJbr0S/2TYM+7840Fwkkv3c2l76I/rdo4zv3ZhAKc3B9YARbChmIoj+W7+cpx1U3
1Sq9GNX0/7X16FkBZF9yR07sXZd0x+hbR6Y5xGiJIDtbuQFjGvlQ9/ARRhAFQFZG
FlNUxu+WUvoRXyR42aG2xjCJzAYs5G7maURS3nKx+PpAy1FoI4FA0RAA1KbGW0qk
UsN3VREy4eoXab1gO5EjPhvxMERKCBp3MIjkf/pdskL2mTIytczZugaJD3KD25pi
WpA6qWgAF4PsZt4sL76G08+KZlsNAR/e84Nhq/hd3+Jfxz7tPGWThnkxVwNyejlv
pagiT68EC55N+kitAQPNM4yEFCzLVLPp8xtc2sDED+JsSe6eyBEUkKl+cdb1B4DO
KlSjjMDXdEa1lgXUqzZGzT8dbRu2dEXoWli0vWN7P50Vpn3P67Yla0t+Z+3mTUoi
dYEM7ifUgbfkNoi9D5pNzEMAIqn8QNpWOLpqDUApy2bPG3owt/zhM9tG75EwFhII
eZLq8lA3uHK6bwLJZwzC/rAeFBSjSLaQqEgU28jxykb8PZNkO88SHmIwAIzzPOl4
HWUPwPSPELSw87vnv2fsqVp10fO02aUV3qIGEvC3jv5QLYh3QHnYG77yjf5Y2MxB
PA/PERfw6L6iYZ9RjyTvEaum9GwRo4t+fvvWAMTGDJpNPs6mqnGwptTAsaer2ZX3
nx1gKFww4aXrB2Y3qwuMIpOmeBdLWyW0BtIN2Fwz18LA2oYcUa7Yhq84TsB6NvGe
M3/ZslNPGxyN7X5a7HvCYEOQqyqg0HVsr8T/87Pn2hLwKiW99S5p448nKCUzgxYe
PuoSCn9oiR1MdXF0DsVu7HndamOxR7wG/AvuXFQegfujovfVGSKzoXH1sOpcgoW6
da79psX3umBDH0VLakELA9xy+yJDDwcQuWVvuB8eIURJrVeUbfaNb8G+O+OCXBRf
iBtU3V2EoYNAPS9sQckOtGmusA2oN5T/EHVR1KzdpEJyQOiT14sdsCISM+qK/v5C
vMV/zD7lvPiJstTY5VquWQCfxGqYzxVcN0GHShHsX8GraVh5mSxJQyDERL7MEtwz
wENcbrHX8vyEpsYmj2OmUDasudA8cB92QbBBbLdgzGlBhJ/JZxWYN8ZToAT0ZGC4
KXt8ZXVEKkxF+Yxy3YVQHzxYjACxVzo/N3mx3KdMJnArA/JiaszCIC2yWRUG1rLD
SJsdn+cKBe7saM/Jj7LEPkNLT87hXZ49Xws56BhC/cRYbaD0l9ZjOLnNh+4pidnZ
s/s0MYQXZOm5JkkheQfH58GlPvU9rnkh1hQq/c9H2UyLmUJhjpq8Nsa3vWrt9zEX
lzLriOvUA1XwUUF08LMozq9tJ8kJbf7Ln/FivdBXPJM7HXO0QHUeVjbNY71o/An7
XBAqTKnjfmxk0LO6mBeXh9xLnkDRkNN1LKr9g1IaGmBBVxi4RX/I+6mePp2rBviT
kfi/EMYdnd5WMBjRTw35kDQBP4y0gBXu/MUQfzc85RQSfIPGUsvRJoPNIQMWF20X
Hw1ps/1ro8bWHf9cOMA30X1hvh462INOrTN+cxgOMm5i7GKN6PKjE4Xk53tgGvYo
6sglVG4IpDibZQtriWJcPdryJuU8y2a57sSgDFBeYcmRBkE//PNfJhYBrlBE3bwu
TRAsmPfFEwfpiqVrmDcto18N1BK17BPcF0e8SAEQmhoLO+eUVZXnk7F+/frIZ1qT
lql0e0TDIaDj3+GqaZ9oPjaCzLax9HTNwM4GPaKr7g+S7zYw6UjnCqT95fUwfNNd
6yojyjIXH1ekIJeudnVjWOs++oXnet4UYvsPbAUe+Q+geOwdKPcKhKCHrgXl4/a9
5b+hEvUEyPouIzxbZgajHv5WwfvN4m3K/XvSQtXZxl7EkKNkCLs/sLUCslEYsDNY
nQmF1L5ng3DvS/XWFZk9Qw3GUf/WtLPSzVRV4bLmnaGHxiauSSea+Q/9WL3EbOO+
WRAq/plV/rJANyppH1Q0OSjNicYA0d4VHSqu2os56cQ//sgoY1JU0Gv1ZefJ+xrC
NPeaxG0H16EfQSnNeo8hxhP2/IX9cIBBbqyQYdF2pWaLKyStB/Klb5QmUXaNL5OP
VdmxrsJeb0tDMGYFCRu2kJR9rGHxWMfxkqvdlD32MRL5U8TJVclI1qfYTTkfOJ0M
uWcrDcd8YpNsplRM63c7NBd8eM2wT2ZRRpzjndmGHUaBGvmDITtPBmb5lFsyOqz+
QRXYHrBb022IRBov4IMb05OvsEJgMtm7yYo7zWLU90OWGC9TED1AH4AtquQvylMN
bob6bkR4cy+pUXMVvSXSa9fwTG9oRpOJy2ORetnnCzwk2V7ahVwVPoWztnzHYJAC
84JjBlR74yPBkMSnnbvfBJMP+5vnJy9rNZpVq/OSMXXYKkbr7aGV9IW6rc2OVYw3
uyORfdoBtAheu7Xfvg7JTZkiOvpBl9iWDcSCsrrt+0Hh7AitHUW+dTtODsr5h9XZ
F56rScjMdsMkkYBwdzHpXHzl9wVsz/DUN+1EFUtGfsng7NfOdvdiZ0HvzyuuO8VD
Wg5RHrDOI3Hl9M6uOlbrx4f2dWSWT2+rOOKWzuGiA2fZNpFF9cnJkzwPfkcPzaGg
IxG9fIXBmmVvOVFYN7R1gEKn0aSdCfhKu5OkQXdtSS6P0QD2xQ+AQ2srJ9Ko8EiA
ApmPXAuGrx1CkyzYxmT0uUbKPiwons23f4dJ34r+8rGxx1VpSlfkuddF84j/PQ3Z
M4G+1TYXivXPLQ3hwG1MhuEnese9/qruCPAqC98tNAuDB0BHc2wkuw1TIIUX7Bpc
ucMGSqmFNXl4gCsDvz76v+A/2PdHmel8HMg+8mc1+7r/qVOW7b/ew9ePl0XTzMOm
+//jjTiDbUEaWGhl1pPIqme1JP9u01MzyUPNDgdqOiRI4sIiOSEQ9eHc3fYcdgiO
3PnJvhbct1E7SJduHB4f1hbhPgbUf+wIp9djp8MFm+guGqjfkNcoSabCXZWKGob0
sfdxCAuqpx4YR6AC+dMZPGvCfuD9QtwTBnVBC/zMavtPI7XVMTJboQRXTka1Nez9
v25oCtrOdO2cwZ6uzQffStAZTGRn0V8pr+2NRNvCvSZeNXlVUUlwsvivdT9D5rlq
kyx0B+t5KLdcoq37BH7ERbQaMMwAZYWBqixSGLmjAlNTnwsXaJeyIlwONb1HIHxa
wjsANvjuoSnK6cJ0ELgCMABpd9nsWjPPX73NzmwgNkyc9uFlVz5nAOMJUd+UUf9g
i3HPYOSEB8fPEYgmB66GSjFhcyuyOvpZt4YpNX60Ti+8eKRcJb3AgCahhIe5mhmr
2Rk4Qw4VLF11kK3ycFgKn+ijK3YLoryzdmKs0nKr9SUasry3mHDEzUHVRo/fXAb4
4Rb67GALiWKuOw2DDX+v8g4bPzOp7Xma0KPTSS7kGcU9cIBmJWW75jPMm38vtJK9
OSoPpSwqWaC6C47daIyf9JgwtpFWA7XWKIhpekuGPTq9InwduJSF1JDsiEbxNz2V
zMfwkfehoAfnSHrzTTFUW4C8DE6PWVZDRZ/56JKMnSJNy2zJvVHo4MSxhJdP7YBC
22ucgAXdGoPjxdlJIHjKv2gNzhvXXbyTDmzwzvZM4ZYykVJIJGO7a8lIobOgdOho
3El6LCBReS8x4YJRtaDJ744XMqE/ttShlRdlf8lcIisUMtPvZkwn2zP6AS2hmz6k
DbxMMBvCelKBB44+tpsjSEK4J6Jmfstbp2El5VjYYNE+ut6eYdRpO5kb5L69xOer
a0uus6qsherSjL5b47YiR0Olq8J70iKroy7KVNwVhothkolcfgsxYxRTyMMmTkei
rla+3sc4HQNfRj/fIntUhHnfRmi5pxxHZHkJubO13Ou2IlMsJDQQv7aylGTzyE2o
p+GcLUjNJo+e2YI/50gA319mHtHqd/U4C0/s474wbq6jkWfJfF4lJZXUZou47pz6
nTejC6/WVPFVPkf0fsF2xu++/4ox4k09y24vp3CMB3zRpOUqdDKH7chwfqFyLTYk
vdF2VvxPXcFVukYe/kHdTohhzpFYSe32Z4nLsML3wV0NlY0ryLIj2M5XQLoxJVl/
X3Taf5yVtQ4OL/Bd5E8kCM7z8A+PnDCgDW8dp431mbo33GZswVSe0iCwuqvex2Tv
VFjuMycqjdsONTXWVgV2geyGiv1t5ML8ZSv4wBg3fhb6YgThZKKC1bfsMPCmL1ec
vLmW4kVHma6mj5OhVoAkI5DtOBFmY0JEQSb5tENq/RHjZK/kHfJjvnVR4cIx8qf4
j9BVy58QrtyxniB4ouQWzNHFNwlqRfsd+56EZ06EHgUt8jFhDwtZb5O+ZpHI+2az
hWIGiUidZYE/IQmAcY3CFiEi+OZUkDF80fb9UyFgme0929Z1bIrLuuQ0lUvuHBZO
hwsJbkaUQ9BYOi49GYhRv+NvJVJKxq7xD92WwKf2MesSZT+nctU5RoehIi0GBNEA
CaGaTQm41b+WUjsfhl+kTornKnOc3i0M+l9DX7sACwZrvmAoHXj5yOcMBiknAanI
MJuSt5pblmsUr/Lftn2yyC4AUYWe6iTMaMXY7CokSm0CouuPnz6ECUS2eUiGne/2
PeK3QRF4Fv2Agqm1/Tp9m44ztYTcX8Zc8moYUYH50Ty5C6vtnoH4MdYKOC7NxI5g
nrbGZ2LT0nivQGTzy/P3vPtlvesXMi4M49381pbf+XAqMR/SPmAqSY05giSJRyz8
vWrOOkAyknd7xkgeUTJtHg5ZvPyLgZIgBA4rl1/SpsFtjHXbSTFF0DwiVpKZsiGL
PAyNXh/isq4vmIKM9UEuY2j9z4/veyMb4K0UsV0WEHhi8hXAFgYayno441h2qZa4
vNp02ZlPDfakIToQKm1QCZ/i+Wv2b03CYjjHzUyWcN04QGnWWbaUhPF2ZXZyaWWU
xAvMrw+wCil6MU5E/55e689G5t92i6IUF5WtzC+mz9n4OANM0MvQrfbF6FZr1QBn
LJizDbT4xy463WoFbSdwlup9SSNySP4IY34hQIk/ZeLeftR1aicyvdDNFfHmc99z
DZKnL4es5L5NJicrgtTY+RpTpdKw8LFZfd1a59z5Z5qbWVBFxR2VZfXM/+ZK1MmG
1mjicDlBL+PG9K8UT9uNQXimsnybIJa2kvSi2Xcbt1hO6OGVkMr9KtumfZe5VPD7
iAudkZ+aV7axlM1oSzAjW/JWnaEVJB1XXXYsJvUBetQHrOHK+D08gfeEs1RiTHuM
SbCGgA/fs/l8PPFqaowrTHxlq6A1W+edOrjvk/DhRST/E4Se9ctqJcFcLpZE90Az
mTyAuvnfiE4g7IGL4MexRujUeZodtoRiPiF8g4L3PQKsZlMHdLK7siZLXqit7mXX
6fSz8JlcfgQMDK2EeLDYcEfMUHVqi7H4hmuNUgHpIoVMULvMhRLmoPl/wE1Dczlk
ey9WRT0nX6uOuqAtneBHM+QzG3N/C5+v5gjXC1f8/LD8vfUILH8oaIKkv7Xjo8BP
EsrbP1c266e4mxaX29K1sbxGgdQjXL7MKUA1TZKQ/Nc20frCpMxfqGIXcW0KMLRW
davTR2kIJhQl+80ewV/0Hb+3xE4M7BxTg2oHLE3dTnIEXMq+/whCdATyfjQ+MyTF
f61AzILZKY5NXN+yh+5npCvaYDU+Kvii3O8POG4wGjzhjJtWE234d8MKfOQ/CRqe
vbbVeydkzjOAvy5SvJyPg9j5sHteeMmcAY/N7XBBRJUKUuMc06eXHnoNRJEIG3sh
E8FpI5bU+TOofSs/0c6hv4uaZQlVk6ZsnQ8XMTlW+71EIxyuMfLR+sthFJsmON4P
DMU6pCWoox8AKzczPWIuqczTrxMsdMEPTRGRgF4nHhle3gXbeYUCCxrHe3x5VKoX
S/h980TWTcs3YimEx0u7m6LxE+6yn7ctL/yHw8rCbcLBKBEIyGH4LmeTlX5GHVci
yyAKyO4/UieOqfh8ggZ2KKONCEQXMjB6EsaqyXuGuQTkQMD0Pox7jaSkaKAlAwao
CNFEKgTK5UlVzDp803xS8h4kIVfscmAYBBhpc7xU2NQ2mGJEXaxGSpWqIAg3SpoW
fe/ufEjB+mM/mOQ0UEfWwt7/7YKDMZiqxWpJvkjFsEfGQjJ8p+a+IdiBjxDHCeMS
amT0HGHdxwm9HJYQAfpCuwUF4B0V99HMKXgRDpLG3hHc1Rg7JsvQWrO/6SEIp00a
oSITK/rf4gk/FpN3d6hAw9FGmHx3KV9UZCmbYp07KyphrX95U65AVZ9xYNYXzz5w
Y07ipeJ3bpL6DUjUPyfDFbMxEa1hFKzY5Z1boOIzC83XTuEHgOdcdOS9X8xaoCGJ
bsw/beghRJwBNU2jm/7aI7uI417lvw/wX0dEZ8xygG2rM2TsuLf00wEXVAgj4Ic4
CM6Rfb/21znMH7penJ2uLickS2oZhvOf2KpRvNtRmZ9/p6fqZrM+1FEHaoD9tTY+
s9AB5+UNRcBzGxd0jxdZRAR2P5g04jRNmnPh4qzAqFp3z8ZmHNRn2+LYjwBxJIvw
DyhS0TB+JnDvoKf/KC0Nv9vhhfOs64a87j2hSefHCQko9g+K7T4oz7WRHkYrtAvp
KUgHW6YSa+4IZbLs9ZgljYPc0fT8wVH7y0DjJOmYlcBbskiY7FjtNtRaqdI5riSY
xzZUZbz16FCTdgytfh104reR1J8T+BQ/u3tPGNe0HqNjJ/d94tjv8CQv+oHWiGDV
wQ/qvGhxy82dsZfUKouANjWzd0TTFSPfmYq8Obz9L4eg2wH6Nxax6VGVS0ljvbB2
s7yf3OBT8dBIvp1G8PPS967kVGygLXCFhX495odhxROj6eo9GHO59T7C+W3wecn3
cSh9qRlBtdfGbnC3HmXbpf8mXJ5WNkxrKMpvmPtOHoMe39JXIEyqBE32u/V45Ikd
UBOatC+++47VpTVBr2JwHMNuoWtSMs0oUoNdOS9vYNEvWPe6IabfWkDsKlfnYwBJ
J4DB7jCZR3IfRnxUsW040LxYJKaxfPpd+TzM29CpF9z4iYILNRZ/MuXkBAsN0P3t
J+TTxOek0iy4icgj3wHa3KoiZD0FdSGPozj4G7KR1e/wGQEeb+iMV4jD3/X4JeBu
Xjmg2anU1uFGWMnU93CFeFPsOeSY/YpJjs7HA060ydEhV5qd4b3VEOhMdzDzpO4r
jgA+BLu4ikpDbDt1MVRNU4w6+mdH+QBgqnjNoeFGm623Og7WZCtyicP6HrcG48UB
sEXaj/rzgYYrofUwfIPVen+1u9YjrLS4Q2Oe2HtYUlDXOa1JvbWZZ+q+W2Ex2SOR
2hISPmJpB7Wqx9bf4x5mLzB2CFuAAC0pgY0S7Mxn0Wi0lyrmE3JbxfSfT/Mg/NAv
Op0Mk615l2CSaawM5olufrj95JQlD+08H0eE5a9FW+XvnRl2T37nfmhdG54XMnPp
12GWQf8lNVVg2ZMV+hknu6alvEeJBXcDUKYQe6nWUhunJ229aATXIOKR/qe+Osgt
aKD3AzBVNX26N+9qGWSHNQL7By+UHWLRMXvKlUAm8OirZWOHS9gYt7WUTVahFLF0
daxcNHyM2YbqoO1OMiLT6tM+nPj1QoezsbJ6KQfjKMz4m8wKegDpfH5d/8qyT0QN
l+p04iPTvlon7feglb66hdUQrCJxwVjPi+OPszb9UgMexCGfhFE6jd6ykEkKHSq5
h1KpwRJNZNifdLeB+qMma9AOSrIV+ApiQK2w7YOnz06wen7n1A4jv/LntOdB5wLZ
D8gH7XRzWNgeRLuw87Nk8YedPTngNWFUL5RJRDcqRYM7nVXv+2/78akzvEunMiNw
u5auWjBvji8vbe0vt+Le+fflBQ9vysGfkY5tenuadp8mLcxJA4Q4TXNgquPuf1Fp
CL6Kk5Pq8NcB1JxbxWB+vqFyumEhizeNA8sUod5NEi1WdfAK636GGS0gYCXJAP2o
13ab3FocE05GLyjkp9MKl3yYvThkpDR2sm5N3TUCzjsignk+i/s6yDTOEDuFV1Vw
KwXsQJ0jG0w637RlOjOJD7GxgJo2RzCfGMhTeOQSAihs4Zz1v4xD1G4rN0pWQ45s
WHsGK4Fv+Vnfwu7gsOHc8Pcah0i2yAnUhkdXat9NGr5lGhF8b4NYrAqLuu55Y1yv
RT3nA37GeIJcyXwReGFUyQWBffBiSlW+cVhLwI9vyYo/jmJ38zwKy9avkgxx3LDV
jmvpQTEnaHic1qq4XGCGInPS86tkL71dy1aTqvxaBQB3PY3Mym0Bup76R74FT/Uz
kVdcd7OxqFpk3CaK6ZOiYjXEXgwWl7ToP9887Y8snCksBoPqCvpfLB+7N4xoWBob
ikqbeL/1hhkzyywp7qjYkbizfn6eufPFDpV4xP6flW4RWJf9alm6kiFSTZWrJtID
5FTI0JAikO6N4NIA7/SBek5E44r+QI+aDVsT8K96fwva3obSK7dU8I960+iUGsQH
Xq9Gg/vz3pqS2IhBLPta5vGxoLBEdlXmkP4u+bfnJIW4GqdFTKFf5UBoEP8BBe/1
frxT0e2K1GfUn5STS9txiGCue5+xVYNjg8WLtDTcR64f/aTm1XWWpGgZRpe9W8Z6
mGeE22E9Lb4S71dPNmPvITnRpUNhf2KC/5byuuknYRRoh2P2m2qu2dv+6UXd6X4o
sRLUKTd/+aNblvM7uUpayfGrEcHXdfdf+Arb4r/jKGhjBKyBJHla5SoPJNR+BX9X
7o302ZtysLO1GiVtBWq1c69O/w/1gBANo3+bQcYK1dWS26cYNouQK99OQYRLZtUJ
9/Y6kzDAQWMZUnsbhBnyzPERR8g4YYXfFlBoXvObBqLyl+8wHeBYYAA61Ye7XryL
IEPlf3d0y4YPpDdOlb5UOxb07aK1jGIoNEliwRUGOiRSjyQtoX9rh+W8xrcEi5te
0FLdQuG9LNTx27Hn1FMtzHV+4ZhmktBEw6RxRnNCl6tJ0gT0Lh4qW4LCdf+xtAS4
p0cVns4AX3UavHO/oX8IBw/MsqyM/ZhblMN8mx+IHKMKR0eWo9DWNCaa2KoQRmwD
E+/EBGS0gCVSvZXxLBkHJqraOU/RBAwP7BI5MGxYZ+h4i7r1B7z0dFmIBPbkDChL
No8ib+8Lt5nRRN0L7PUqNEfpssg9TFNequfh3/YHD9ZPjScClH4mj+Spo9wKQ1dz
VQPPntzu3DYYK+cgJoJGd83VqgP2mV643pMtO84kOeiyXmxJ512a7SN+k0rlUYaa
r5hYh26EHkmIcAwNDX/+sxaqhLbDBakKeVzUi9LUQtCG/J7zofGgagncCmppv1u0
G0t9BR8ANcPkQUdElQDoH3X5BAVGw2ouTWmbC0hLhubP3tX8X1IC9HBKCWHULBqB
3YZHkrIvZV4yTaMMjJ4J5BbAulBB4QHvjdj+Q5J3DSz1O+vCX6eLgkcVrvPBYMjW
QWP8YmnOkpWTM83nFtPeAu6DbW6Dgz55Sp5lvAbHDZy+nVK9fzl4T7GWitQReMJZ
zkEq8V9CGzIn42QFoVthPSsRqop4Xq4RDgEENhuNVu9g/8UH3xQsYmcNC9CV6eKT
cOtPYqlTj1UXNGt8StcPxhGXTQyTH9p3bqW+o7Q7/yyIN+APaqQI6Hz+gFFnrvRK
xFZuttUVaR2z4AdGL6/pN5E6IsKPFWxZ2v8DblHvb5EyO+dL2U2ILCuenNE09DE4
d8BSVV0KJ40vBRyNEViwmdI6M+hKtjRf4+aV0n2z2sg0UlYCqy8O8g+WVV85skx2
ZN+Z0px/xDc4GVMuKX9rghsvtFSUwBUCFjUqtnVppfTJth+aPeUmJcLWetpYNQLb
XFQu6eM/C/umc6LhgobTbukEe366rKf99bs6C5mFINi7PUql/XWtr9GEiJgYaOPh
/x7111rzllSq8jiRvqeukVbwDkWUht4yDMLCOjC9ICxL/zrkcoBcBZug0wU31sig
D4fTuxyKL0lAgsi6OJL4zClyOG9sxMGJdm6Q3htXkhm5MbbpH+ffa4WrsZ2CS8fj
4HpIS9zOR+26hTmUWhy3lqkNGYt4x2q00enJyaP40c7m0GnugZ096IZ3nk/Xqqm3
ldyXkpt8HwgK4hoZQh1VZp2FVHNiUe7znwgQfwlpJJ0qtzBtpvArSvZwk4gcZYcV
ix2YoyBVwoV5ZL8qAdIJ2e6DDoRH8/81kFzMIK1mpUKcsGQPO9TRldt8xMj0b71a
NflhwHPzqFf2IyQBwzt3p5nXnmNiBgr0TglDsyKhD1WY1g52p4GgOsuWMgUZKhWZ
l7oSxP0Gfn77FxxdN7cYfcNEJllPHdSTPEGsVGua43BEq796yebqvgJF0Jg1OaJs
00uH2pCXPO7ultJLMDrSVk6+Rvn8pOnhFxg87dBqe/bGiP5yS8ano47wHzdyMXi9
7xU4cOpr8mHCp4dL6Kvj/zj8cyW740JoTUyyCfX1E+1RVDqd1+Zn/sfXyjuo0ait
wJLWpxzrcjY3ECPpyRHM/UDRRGepGTm/MJB/npHqXEeO7FP0yNdRtjgkMnsCr5Hp
jtqdKHB1nAiIui7+fwbhj8qT8xxG+qfmXQvc1BL24P18GXzbU5z7+3EpaqX/wqCo
i7YERdccwHEYTGjsUhomWANC4sZ8DluGaDijD6Y0jT7mrbPWM9wx5DGsTXjOsebN
UM5Y9xsphIqdHzBuH8QzI6y5c793CJ16308WifpZLabCeAuK++yYwLVj+jpU7xew
n6+0F91vur4ziqeRGsbot779Fl8xHStUVTdUdYyY3AHPCIcQvVggqebNYBeee2zP
Lt96B9SZIurKaTiftF8jR70wGiRW+xGyaqBzpg7oNKdY8WxObKNsXnJXZ/Aa4SfK
H+RksBvTkX8gD6gBDhGJ67Drg7WI9Z6LxdZESNdKVS1mVEc0Tbz0NwH5C0Oyrpcj
ETgbHK0EGpXlBBFzIupsuaWZF1Qj5f5H/alKyYFh7U75hWQIUWgDQl9CSta1F75A
IgRxFQ/gmx/CipAYcm72vCOU80vgmCaGMwyP0qaR0azIEdTe9L7lGiJ/0/DVNlJm
p07RBz+8xnL/iG+KHKqqtB/VFZh6Lv4Ua/1FT+qtotMDTevMh/A3NLRl44QwApDG
Zsd1xeFu+LsJ0B2o1Us2bcYOFEKIQ6DyDEBDmJahjx7svWk6O6tYL1CvyhGWuSOC
yGEmPXDPg8NAJHid9LMyyszUyCuhoTxqPwT3H/KtTScpfBeqBLo06DlfgZQIzEqA
Il7BBshHpoGKGyEDI4g19ZDs0UY2loRHgFFKP+vONhAmyWrockqp9kwsphnExMUK
bVIrXdmFt0QBvbcIoqjgQQpIdObI/lns2GgbxuAZfwH+9Dtagh9Yn4j8C6Xn7m5G
IXdMfR2BFz+K4EgyPWe6n0lonVoJv3NpyQXiMYovP36ZFdZB6AOQWYlBNhQPnT7+
lDKNYYm6BslQS2uWlTiTv++ToUzcwtqmSj/ET5QTLlOBrnAidwzkSrQTbQ2x0H8Q
ZCUDDJFuHBVmoo4dhFfv87zM741EbyT8t/Ef2+i/1W26S9Vuo9yxyO4toJ0uvgaB
3q1FHzApHb9I0b6op7DNauMFTA9Kx6enpNtOHIYVL3zAvCqhIauvjBy4sUmcfP1f
+U2IRqNB2+MVvn+we2xJZpLi6pi5kWmkwo8ygY069v+mF72uQ26ZkDEaFW8Vs8Df
1th2xMXCm7zZ9eDH1PxT7xVvwK+JNBkTp0LIrYqXlvU3cTUwuuJR4hRRqDHXXayE
1MXUwNXBMt1ralW7aj03VtENvGArbpHOMhwA97ABaJxOKGiiJikZXfkonOuUbyfh
1PAnQ8mwvW1bknLMgyCKyHS3GN2I3aD9NAbTOQt2s3wzTbYmzil19egJBJZjJf5A
jgC0Ge8i1CPDfqYbwQ6bJ4vPyY86fgf85cVsMiVu3kO3GAKJEFyXNtlLtxnJpRuF
GqysxLaX8Y1X6yBMAz20qBuYVNZ1rvCHkJFIoWFatTwS1iSVvR11jeoiDBZVQvfo
yItypiCkev/8xDuXdaO3L5aNdx7GdBr/Y7KVWgw1rxMZdZmErl0dQUNPJazA6hEJ
fwAtrDnzljpj1XXuRMrz0QsZfi+SRzUOxgTA5Ba1/2KBSz+S04HJ2X7H0i7t7H1Q
2dpZ3g03xX0aQqO7pfxZIwpsfOF87AIZtuLM4stuN+iwQrtfWA940Ou16WwZcTRF
FDPeqNYLF9k4TcMtG7nlEZGq63y2yD3zof/HuZAw+IMW6Jc8tB1xUMaKqFElMnru
pQ+jLrgSi/INTliC7YSOn34mPF46PSkriNaL+VSRKY9J+zicUJRo9/nRdIbu0rDZ
YYhfnCOpTgswY3CYtNfrsRHhdjMlnymDxM6SmEr0xZ0mbhR3jzELc9Z5/+CU3pf+
52DyqDYnDLlTyugE3t6xhSxay0YKElct9PM1j0kYcQBoWSkGjD04NhH2NIawdJlF
Xng3dLy6i1188dmyCuuyg0ga0xJQQaiVwYMlRavlrfRophMj3YERPvi8DTDVguL8
Cy1JzC4CTjA9hVhD9L/4zwh6rfDxcYUlPRLfD3NE0/9Z7KfQgc/pu5pWYfFvNBCK
vg6prEgNTo8B5s+zoLAsbB347SmP17Gpu6dtbYDne0MyXDrExIq9MeezhQ6bkZyo
GdzTsPxHFixcbAC/16m4obVxhQZHzjkxhgn3nBO7vx6rhDDd7SXO0mkkjTwo4XOH
Xw35qSDe0ZU1LA6W7fTOQZudVtQl9I9RFXS0gW8OyEw2Zt5/zOxBypnmE8BBGweD
yGjri3SILmedJiIHKmhNy3ijZts+OyMKXSh5JTeGbQnu47nXb+xI0PZT/X/TgvBu
FPM5qQV8juwbSY1r0IhKgHZ64AMAydrSnL+dEbGJBxr4HDEQm5Sj6/DJKMNRLIrn
wkmqUDNRTDlyIOp9SezQvSPWj4IzNCvUmWMvGAG/h/9g+019y/XKB3NVXP//+Yp1
hEOLCCdCC55DIIF7dZ3tsq6P9fkAyDlR4RL8T9W/vLmr62cQAteh671AbnLCBfnC
F/x+qdUKv/nDc0qJi9jIDnlDXm9hfj1bvrH0VyStXCBqL1cMAHvk7RtD17/iXE/O
9D1ApYD/o8yVes44XpgGXq+cWPBtR732hU6uYiH5K5X5t5x3EGK/+pg/9ba5ZCXT
fjYDtRD0NGDLS6AYMExRV2g8DlZ2CJhU8UfXYdZ3Ruarc2AHBPC483Nu4x0BVqI9
A/VgW5wAX22PTMGgT+n1gGq+yNXNCoXcQXZanKrkoeF9Gzf8rq6W1IzsrEX6VEe5
JVasKAg0sAa/7vZ7sA0NseegiOmaXYXUq6V2Tu06b3GF6wgfdS77VCqra3jg/3Cf
Arvx5Js4XmqAyPKQ8n4yfed4Y5y6wQcCuDJ1xM9T6KIQoK1OmTqdBBf8vHwdY4ud
vKwO7oeE0Y7XSJfP27YLDBO3u/l9rYWjRX0IP094FegtznQuYIMghsBNmrmwDWr8
nXv+GbqxplGVF5puNjtacucSnSQDtIdUB0ha0tePD1c3Cw4Bhr2jnwELu9pmW835
wjsrhd3WxOz8FSn4V+oWkeN1Uh/Qs64sb/4qL67dFnhA7KCEu7RvmqZvN81kYzKK
sxqBwDYZCiiWXJpY2rjN+XXOvv0PIUS7NbYVNT5svYaRg1pesmqSzs3wj0OoiAqM
7plZgb7AiUDSRVWlgPjMDvu43OAvY/9FkiuWdRv2sgJTep4ChuCRFFIgUckRh2dR
EDsjSb822OxByTDg3wiaVryYItmMMpSOHz5M1+O/p1psO0VECBBxXbxo62SDFUU6
sqLCgMHwMHNPYh9JrXWvFPz3pruXTMZ5LrsqeCade6upT0GdyUtaq6b7QTLNOu0L
418Y/NVSyXPhL8ULdOaC7cTawFffZqq5p/tvjoLL+qlU8ZplJB0awCysmlnHGD9Z
bUbL8oBFRKpjmISnKhEGvLqApNDDFkFhbamlZPeiktPJfLJwBChnNPaaGuO2+QYj
c12h51vu1+i+g2alXwzAKhraBPKmwCkcbLhRCbDkCy2yNZBrJdX8QiNBCr6jbepg
qanlTwsubm/+A+034s98NApZZ3s0KsbYhfnEaYCDYBAQebdD4z8vAmkXiG8naHPv
gCWB0MsWg8asBwqC9gUxxRIo9YMe01e8avd+nfQxUN+gOhWEYYSsLqJ5amk0wXz3
uKfg8KSSAy8x+2C6V+y3Cyfdw78fvSoU3tTlBLuIXNNrcwtMLCkUqLfFIOS4zWEp
xCBNjoZyJBMaJhkWADYnTBMTER4ga9wLNM2GbRRCTqzYmsQbQHMsJVI7YC5rlXAd
ynOSnTczU2CPgypxCpw52O1LbDWfChtpuPOFVQfnUD2CYFOKSvEX+4nLfi4VUl6j
eLVvwrS4jm1uwqJeRQizKGqrP6Q86X976IOH17YmZQzZI9Tvx9l5vFpUf03baiY5
c6KFm48A4Rf/C0nQWYlm5IVBMB2iwZeTP//ugJP6+s2ZiwZD7YV1l349HQdqKDgF
RwIfdPFripRtEj4QlHaFvkqCpK2Ux93iIi2CtXRfbLGiFo61SYGBpcTB6tyDCpNV
UIo0Lxpu0qZ8VdgYC+vBNaPbArxNZgDSYZccGfMxsFGmmL9LSGxsac5G6NN8rf3t
9lGVVmx0wQiwtphEO+cqpGSIrf/04tfDcjtToJjLLAWYcl9k3izQBWm/2lPUvJOr
xGc1U780rz2dp5dyfa8ramgPQjXK2Fq7J3UqxdCJ38zd0pBVlLMmO+L1ZDD0fRXs
BHJkRtMwc5o0lM0CRSF+bi8SJP6BM8Lsq13+SBZkSyJedBzy9Dfj6QrOknfNDD1w
cedXAQ3Heaug4VBQ5Pi8Wi2IvVoRcMdyTdWR0k0BrdN5cwnF/gfCYjeuOQdb+IBo
K4qLDQ4rGGjbKsQ8ROsK7uk6sJU2MbGenznN/q6F2wNoF0v040FwPXgKMSJ7Q+PL
4Tce0wDOIwlcdiPfrk44yJj8cLWx9gOlJqQ4HuD0xninKsqaZb5Z3T8nb5p5j4Yo
HN1nRX9kjZa3Rff5Nh2YeCR1MCmxnPtvvVoonn79adQpdks+kb9wW+BB9t/cGyS9
GeWUwWkJBjM+kVzAnWckj7Es7AtUg2FRxMig1EmB2a6a2jK98/GTkIpYxaNvF+M+
PaGEFj2hkQjStszCJFngiP3SB+tsM5r8na3xrj9gyWw2uHuqaJhUvT7yREwRhlBL
TYpMyojbAGl26Cg2uwHFSMyy6beUPSjXmQDK9YM5Rm4LPt4VrJKZs0CWr4HsMxjO
LQdWJ//VjghvnI8E0WNMLQUiTUBS5N3Ge3p+LnQ6xofdZ/5dbr/mVhbJPrnphVHd
JUOIpiKj4xLqOIons3mlTmgvUWC/5UIg/pzwbqZ7eN+APzv+WC56EmjwaSwbx1rD
RtOy7YNWcRPLV2WVXKVUBXagkGgM8Sp6a0Lhc7WIMdeGQObpBw/V4WXPAP4Do4Ay
fNsEUK+Yb9Nn8McEWzLbcUn/N4pEyYqj8QCjx5sveZTNpBRmncE5/9eAbZ2x3xSp
bmS+Bur3A7tMOt1VgWFsCDrVPWJjaqCRuLhUT1X+LnqwPo8n0UveIhdfAPtqpP50
Isz5ZbJGUdfVol9qJ5appUZH1ORa6nq0wm1hJjhQDRRdZ0Z7uRGFkz9e5Hbh5yXa
MertKEkKHRYyTnVe1nzNYtFMv9o6d5fuoOuEAVJ+NGli/Y8Ywq8I05hVbye1J5u2
NTw6CyUyP8LXy2+426F1DaD5/TMIbeEz4j2pPD8hFuRNRRUkIWYtqdqiZ+WQVfzM
zUewvu0PBxRIEdL3fqteiU9TVuQOf0ZXzLHubSEwGb4N/JbEggBPb5+lsCzYYPob
bJ/aOVyETgH8UeHTMqR8o8gD2aqx4am4R4+kOrN1xK3z/Sr4m7aQUglF4JROejWc
00Sjz6mEznDmyZwmbMwba3x6XbDVf5lK7gn0prBMRk6GiKs9gQDMQR2hzynfYoC4
vorT5zb4cAtReRwNjEC7xin9tZ1ZAPKuoS7NI3P09kwHvbUBecWjNQ8wPKRhPiNn
pWwZfXaj5uhty3pFlbK4V1jfOSCnmItPEkQh1tfYEib6E+XAEvvnzw5Oh63KudAv
wqx8XgQ0G3QGxxOAOYSkVLVECByYGp7rYQ6EhtwAUv+RNAPeH2fp/3JLmoom/F1s
7DRAxTGT5KhJFfZPxuSh4JqiqzVsXhyNpKXCNGUCXqaHriZM+e8K5/rKVUs7B2UE
0aZlRyHYv5AVK+ujGe3msoKgZIBf0yZBYvTTNDeXp1fukw7q4Tftfp9Vc7xmKX7m
KHDESCHpi/PxsosNprze4Obqfb9LVDB9zW61evHKRippy+VYp3cQDmms9WxrCnJ9
aJqjcRhvZOxyeksaPAkl/8QdF6ZRbR6EXtdhb8GMf2M662ovnF9GmE4GOUjVJlpp
HCjr5b88Qh17dyX2F7Gybs6aNRc9CPV7xbnIdbMpREioYgsGn8nQujxfp4fT3+x6
1JLQUqfUwJO20vG5RvqYREQ10dYCjP2HyEAbebG6kVI3CU4HzeKX5qqM/f/iDTl6
xq7aT8Y+k+mKVOCMyjwfNLbeR4RWXIevZb7zzb1BKR18FthzzyqCrYVVTkFhRSJg
2jWSqnejXzQqU3XF/wYleStfuCBvQrBCifMqywEWFX62XXOVOxqyWInK1Q0Phu3L
jjXj1RiD8+aVyJT1MZc5VjSYa/vAuEOQvdqcD/BFCBP0ZFqQ4TvMBYy2L1s5PjNl
n9+neBOEHlVoQ3sxn6pCRGLInML6hezNrJctLBhsSnTv8gpQ5BmlAQjHfOdj1mv/
aVp807fcb6jCPMlllwJhYaZr9bXyHHMmFUjra8UEQrp+AMEP7jzVcocosyGYayVE
SZg6MNxAWsi0MmYa76ycWqFunFQnQtVxPZCnxE4jaFs1ku2EbOIPCDh+6JgwSVBs
3czlgzzXOsYotXMgfhxm9dhCWwG9seq7CTLQ1g5a8GoA1N8VfOeTkZi7uhATkaQe
qFyWZ8rBg5CFU6VjsmXGrtidW3beObFlRON7h9cKh3xJGVnaox8l4UanpnCq05gm
jv628aVGnyALjC6EXVVdPRmdI24imEWlaRMA0WAMSC0nkGjrWnjAIgBC1GiJNvxm
UGSm+6pCIesrElZh5JsIz0t6Y19L8Bi3l/u4DKBMUVx4SelV0zRYFIvNXVu9F7Bk
bq7Fa327GwglfNG+DcI7PDf376D+BvCDQ2AFnIujdLOu9KkmyTzfe+54JeXimxSB
h0vpPKGpK2L/6DZeB1ERZEek3T6YbYZbYi6OIvs+350QmD/chynEeAJUnxNFfdbv
wMknb5ZIDGK0j8KYd0+ApdVSfKPaNLSnEGvlDv9v6oZF9Ox+da+PnnwFRi10eCmP
HIRcKwT09/vo+wGQF9Q9Yd+5hz1HyEtHDj9dvcKYguVY72SKn8mzqX+f3QDaG3M6
BJP6QsQxGp48zoVCIVBBbrfpGfZv3j2NEJ1Fqvxlzk+aoZKasQl1hRcNsazUHzBb
jobPARS+JAkOzQUZeqPT/bGN50W/XEJYODDYyz9H8od0YN+n6SWztoEsAXME8fth
NjvETs+IIa13vVr9GKTRZgOKNYXoB98S5MnTCxbrXkf0rjzI7Lrg/4nzqRxAAXKr
/DAdYX0V/ze2S637o1bzKxH8Wb3AVqhy5+m0t1KWz6KG9BsF8UcXaCfLLmmoDTWe
Usovizj+d1QHMii6Cuk1I7tv1Ta1J3VG1akWysYciHeNLrxB6/0Jhgi5NTRZwn+F
PY7oHYuMq5anoUdNItbyeunQ8EBZ1XidanJZPZl/mXW39elMjw1mHSThA+YomEWX
UHaPld4hbjoEY5NyadVWxDceoa3DkgGCP1j51OC/mPKoj6LE/aFLvTyczLq2uM/q
dgqxRxBf66baHUDowhqPw8lHOrx9I68L4lodEV41t/bMzIByk5pmY3NRrWLBxSB/
4yzE0PBZBjERs3kXuoq/dwelKVXhuyTRyu5ATrGuGmN3jdnXsgWdPtZCuzYxw/If
Po3jfJRO4Tvt7eBJNrFH/N2ht+GX7MWGgIElsfBzB+oSzl84bk3qE1FpEZpPeFpx
NskagPqR0jNtlf1Ste1zcfiF/tNeqJ0JDgW1164wvRY0ZnfnOP0NHBmHA9OUjHfe
0Bl+cH3qM+ezGE2i/uKS/7jSXeipuE6728I/hixNyCOK1Akd347AbZ8vPI8BE8vj
OWYfYMazhJX6Ey/JQacMCgaevQsYoiF6BJnHjfNW2U/Dzzl5om7WMY21OcGhlXlw
zoodXSFjLrDvjwi6pKkCcwEUcoG3SLugHXkSxcYsCHw+l6EiNzPOXCYd34ZF6oy4
eYUr88NUmkIYknuLfvrHrcdcJn/pGaI9n3RY+3Rds84yjPI9fDrncCxAW/JvFx7n
2lsDnt1+B5f6Jkkh0r9W48bihUSVqOB/8fkSlnBCJiqBrUrjU1riFCtuIVIpX/Az
USTDb18yo+bZYjnhhAQJ8WVuw2OTVe7Nk2s0LOHfi2BQ5Id1hbOs3V35W0/Dahap
zZ+x/16RSADlya/8WCv247wvviYReU7QRRZai7C9VmCZhUuS7rOflBxfTkTG81Vk
adq4/lRzCxKvgdib02M4aLLTneQQ1ikISwpPkIZpVWOVFlVnfXOr1lXSn1ND/Hna
6iuJbnEyK/zBj73o6hbNd7GDHUv2fAJ+MtSqDMvCyoFXlIFZQrbhwftjbXQZaxyW
Im/E5c8I+QxxlVash1vH0yr0mEXigItMxVWMfAvCUhr+gbjEZ7p8f3+1wPUcyUIu
819AD05ec1Ezl7w0pkAR30XSItNvuanPTcKDw6x05oZAqSClx9QIA1Xlx78wGpmE
ZrzebfJlodaoCduNWvrEmvH9iT6+YjlIchjqs94fjeBuSCaEGZvRv18FhwHeuriS
2OwApQ9kX2Lyvnfp0aL4Ou6UUlF1pW+UE+T3IYHgrnEDPCGvE0nhG8i7Ax9/XbZr
iKC2+g3OK8/hFTX7AXM9lM4hjgsVANmAqlb0wDfvUxk68a0MlzlOUsBFnsIK52bH
zO2Pb3hkxIXVorsGWFDqF0aPfh0QNW29qtv4nq7MJhLq5p2DEreqXvyxnJmBqPTB
scPyQ/cWQQNZQAUeYCUBI8FpkCB/PxxcPhDd5yvGZ4FP911yP3WtC5bI9LdVi2Xt
Bdc2QwWtZ0kizFrRE5WDVWQn8ueh/g+fZgM1uSBnb9m3WVRbmV3Jq9ejFUuJlT1z
dONHMdW6hGAHWKd0ujyAAez78h4br7MPZBTU5E3Hvp1DBfUHKNaVtpS1VzUbHqFS
OkTGtPELVYsuPsqxPxqc8sX1fH3rsMrgbab+Mq/1MKJ/2uYWyUExsD2/6SptIWwq
8dBN9wZ6i2tC5Isz/hecdCkFL1KJPanpOpC7a2T+PZGX5r686rlcztOBHNUn31WN
96TnKaNrZ+ZiXkVjL6an+BYQuEd7Jvhb7Oi8dVmeek7ONVTPHZvvrizWqrzZILrz
viBi7sIBv/58yGVCptpplurejE1TWslGpynq4lGYioIB0NAI2CV/e/SXH8WDJB0E
6AiaY4h0Roj8gm7yFu7PUJOvqoCMPu+tMdp/oUwhgmIpK9AbhhBX4KqYLfHHMaF1
FP6dj1sajp1NPCnBXfPZur6ArlO6yenJW780j20AMrY8D0rrSGe1+w1PTY6HZCQv
+mUoPigEA/c17d4S+zUtSBMPFFk+w7hkdHZl4VF23c2ObZt3a4811U6UhzCpGFYD
IKW3jnq0cdNddZ+PinpS9FLvR4QpfLfuO3kdkJqVwysNEPhxB+JITOCDcLLJzSGd
fBJYcVaGu0430soAoy0H9fhGrqU7WZz8ZlsNenqDsnXrFqbN4SwHmI+aJUq8s2ng
9gfGyMy4dHMkp0JXXqCYvX/0W6DjzyB8Ojd3Y5+pUn34Mj+6PkGIbcDg6g6TLEu8
tFVO7DK1PZVJDjMROERKGo9UyZ7M8pufJBsOpfNNhNp2Dare/xh9g+oPtEuRpoJC
hScoUd7DLmfc861M9xVj20otLgjjBRjkSoRKKuvrtsD//PfVxgJV/tlI5MY1aS/o
+hLFNLp3uJYXeD7ZvMhkrbP+l7zDBjr/fYHhH7AOBa1Fk3R6gSzEQEe1nOuZGV2Q
XhqiX+BFSQ+Oy1AqHSLPeTder0nuu9EvBx5Yt61o8XxvbYdAeBzQh5Fj+ZrWmUbC
qaorl06nFr4ZunRQ7whiA3qb7X76d9IR4FBOIcHERX/69F7xAe1z10MizTVvLM9q
sa7aj5mpYt11xEupx+FGtk5wmqVljHnCzMIQ8A8OgOqlbUFSptSGP8xJsbvi7PQu
MmuOijI0q023uZFonFirONU/yGn7RlKkdKrZVlZxbkdXhJChnfBkw38FwmWAMh+q
IyaSkzh6i6EJ/Tr1EIUXc7WFrvFSdXjC9aDtQPzlI730r7cxc5emEM21jmZpUw1Q
Siey2BvLH1LCT/k14RYdRIajd0sfppjx4HYWv5+Y/+yZnh6S5/BrcFwK6phgP1QT
ULOWeKcAlh2Gtdprgpedy/KUNZOGdwsZK4MgtuufL9JDD4JaPxOyXD89p9BYWVUM
KUQFlav7IR9Kx4m7rOWJOzO+gF3gFX2NGR2p4lMqFpcjfoaEFxMtqFevVxnrHhXs
+UX5JjV1XxCG+aWoRyNMZV3RtzCn3zepKkxKAF9kwJPvJIswsKUafr97PYW3zqch
IOO1hyOfq3sFzofDAqlrEkcV+sBl1sPML4sa9TbwLYrrxi4obtz1ZZSqdnSuPYsj
Gi5knlNh9Pi+TK+D9XpKTfr/O7KpGo+ber5dX2bMipANMCEVFubiGaj9mDu+X6Ko
3wYs6+0YZ12U1etGp8H5LCPCMtP1aUoRI6cRlD95G0Us0u+ToKyd4NBvirX+ts+B
E02CMu9Fvazve5hBbJ/4XnjxXyNYwHeahjojPpDUOegpIVQDvxs94r87b0HBOJpo
FtU7w72YApm0Yutbd3xPSE9Nft9kCWwa9Qp/8iLBdJNiDXshdATumaX238VKtU7q
vDZKdeC31EhdyyxvH4Dd7dH/r614GWhcLVyFM3zJFjvG/G3v15peASYUIsaBbnbc
Xu30Gla0OraQt+Eb22fmhfCTgX+wqJNmQnsdbTGirswrj+uPg1zhmlHfoAWltJPQ
cmP+o3azCyiCULtf3zP3TaItBwX/mtkmVuMvMEKLqMo4VdLnqCpXruAIRML/90Se
l2KQ5LfKlpj15E+DPj3IHHPY0qB1rIvHDhohHD1oWt8+wExVRdgLJ45YVlJbJKKP
afRf2/ek+re5n6nl8xk1r71KV5Cf6igo3JXg6Jq59xy6KrEdF+qCq+DavDK3olsf
HS9lWdC50W5ohBr+drmi9o2AdA3boydETeW6PK9gfUgHHItCLRXf0YDTt0CZrQrj
sLK8HmCW7wK7d8hAe4kQjZZtGQZGbFXyvV5Oe99mGUuJ98Cmi2nNQpf0PAZNiG3q
jlh/uvj+ApMbmAXbhWy9Wdy6Ojbpvr0rMBWSbngfgmWFLjW3kC3Ocb2OfDxQ4I3t
kMLB/8bD6ks0N2ObSW5SYJ6uE+4c+Tytm8aB+XA/864cHOTW/FB99Rgpu2VPte9V
UP4sje5ofJ8/ZzAFsZwUlQKS0oSEKbxp0A5+6+jTr3/dGwtnbSxs7y7/Bt0Rsqh+
/K4+q6cDp0vAHzH415AKMs0gY/W9X6mpJIfrrJjtwVFlpcBjeG+jhjhMFO63a3oG
NQFfWI2iCwkikovrreSblMvJgegeXAkierpSytPmJ6macKi6XoRi8Yw7VS+9KQhT
c4uGqziSOnHlWFAghA3FM/LBHHMfMoPdw3YAWB5aYubdNba2mxmsqv52cWcosCu6
sWeOEjOLUSVTERSOYsX1K8dsTTQcUCdQfM3Q3aNMuZ5dk15o5mJkEG7BvFAVL4UP
aq2T3K6cEVYJYBJ8aUy3D1DFamQUsM+ARrootiLrw11wpmU4ZPgSjMeSoIFoxoiQ
emBnNJsPWRLR1akpc7q7O3vNh9ivsVutZ/LlEFKkFX3qLl5NUv5iHJNJGogqu1yT
Qd3Sts94siWgbWPcvgjd+hpSmHD1L3i7S1RRA581d6ysLsfQObieby2E6okDGahX
I41rBN7m/IqShwNE6EmZnZh86nAiE7R48OLqi5AFFMvf9yHDDU7YsSQ+7rrD6YDU
nAOwORuODMbOJfbWYV1mNnmQFpdurs+Co8iZeuLhWGTA2iqU/8t7Nugzx8KXmSoP
GB2RdEOwbICzL/tznZgMAtr4+f54R4O51MN37xN0DPtnHwdH+JSKzkZtOUNEA0tO
iGjB5F+xN00IGeVLi1DCWg4MC91CUOz1t4y270FkaNCxEWRhvos2AGwSyI9fSgSN
oebmQNBi116WO65rFGow0oI2b5DvJbsipXbgysaQhBufAjLhyvksQcBFU/1VVgKw
L11j3/CsjKqgVx94LEkdsrupC4bGP5oqJAEmqJ6c6krzSHo4H8R2WU7tr/msi66q
EHnUoSAMhKr7vAnAd/xC8KNDGqHPOAfpfFX/PY7QVwkpI73xHndCfatDs8At+vI/
zDRwx4xs7zQ0hlitZQ8dmG/afzEwxK6k1HWREOxzlEJxeJtBruOZsmLnPp01YgoX
UzWqnzR7Yiie8moRJNM+3d7BJCYsJbLFl15CIlBZD2B4luEWtxnzKCsMlqSrrFu7
cU6x2UYY3HkGxEJ2C3ZqNKkpOQmlNd4H+oCY8tOk+ADTJ1MWXmHP0A2RsM6IcfqJ
bRwZqxOWOgisP5QbAzR+QfRDJkuQT/ZJF1BUxaCeb/AhVuADGKkTuC4c1r+hURMz
qb3aPcNt892JX79ljiAdkK7rWewrfVsweeFaGYMSyTa4kDlGKy0sH1ORjq/E5sUP
cuYaQDn25pbChvi2NV4Lp3DWsejuOYHfZpCpvRYD1eqMsU5BTb++XKQJ/ziHC5Vo
IHOcLZDQyTek28YJcoCoUz98vT4+CWu8re+lMsoPmtoZYxr7g8e5WOah6NKwCiey
iO6HzQzGSEi6bqhD6RJ+zwZDqgrlT0tDzZXFGOsEZshEk39cAqa8x69sJFrCV99h
y5q9zKBtQD8hbmZxVnRCu+kQCwXswRlb0HiuJLTmjtal4scjd9lSUGWYpo5sQ84N
dGt1Xhg4zWDpfKehpRf6icGxZf7cJgKPUdF36nqYcJc3nWPiW8X5hMaEUd3IrgB9
iIfhW8YCveSCQ9yi4hKFSBQCI2M/5WWzdbEBvOdkonTSdTZbFSNGQROUaffaZT/1
poIevwbY5ARy8u4xy3vlILHhJ9kZJa5W+qYlIVuhbkdZV+7oe6D76nUY6375180B
LJiRuAxaISuRxdWlO9Jd6V9JrbIo99JANXiA6Z/ltFar+v8+eUEoyhDyawUYBVwf
OMKJXWcvrKiwYCLoM9gr/0cDa4dcEk0AIqBbHv6/ucEl91ax8XjyTuFOuXR/HOlN
Gr8yCNfsCu42KUwEqJE6LdrZtZEah75RvSwZs0VHotCPhPK02+o0rGvJxwmYhuki
8IPe1kuib5ej/20J6WaXTc5Ip7ZBEzGMIRnstzU2e6tUzdMZCi6Ge6qZpnC/D5y9
D0n+yFH8DNgfgcnujkFn0vp1I26956HcU9DmVA0bqLxuSBQdBlJf+mGWFVrqwYhb
/rTvOOJiP92kgL8NzKELPVTuSFnKuIDR367bifa/0l9JRtyRDdumbO96o8nrb/Ad
eVWwg4ZbauEe5d8qcGO4534/UGV5sbIFKz13rRokIfPr+4RQmne5nreRUy22BZkf
JPYv2rNQRVYjf5TfKT3sX9ojWxNJid54yPRMUOo+oAHBjuXDtJkuiItF/elwVOiJ
WfvloyncU8gptswR5wz7IqCbcOc+4bnbu1nCshyQ679TtDLm/s5VTk2oZ9rNDP6Y
FzaPU9xE4Yqw/sBtYNDTmCZKelx7kPs5YECbHQRX0aQBQX5+SgcYrfYJPg5Lrs74
Ss0wEkCy5aTeAKI5kVkpV+Lmq17xfkeqS/CgO1m0PjnDG36YxJWryEldIKqnt0FR
kw7W4ItXUisNL0vQIJklUIdIRAV9aTONnWgglTrXXsTBziCxbIuByV9GzAURNbKS
ZXvcEUWIn0F5CML784WqXlLqxkQDnpi0Lrjw47cSLggzK3vhew7K+I94w4ngGs0z
Ed76t+ajvmujjFW1VoxRcXFB7nL+ER02OGgRU9yzl31vKpW5/mbdyZEpmuIMzX3Y
SA0Gfi5BRVS3kNh3f0LbwNE67AX7PKdLkRoS1ruMljKo7JylHZB/yKf3a9VV7Edr
shGbH/moy33EqzRVmu1nzLTnPa6saK3PVUuSCmvehIWUGLKMRjSmrGr/arRSHJKQ
0bqkcQR8cW3DIoibbAzk73HV0Jju8HVRGQPoc/NhCADUWsBi1ZnPLewbv9gqOK/l
M3a5TUsoBnvd21tLmZVqh4jk8FPMd+BQsSfEezZHENLXf9BZYMa7P8ZcA2nLO4Nd
LTaXr0VS/aus6+FQou9Z3U8Owe+SfqS0P03BDCrjpYoVPARw1QhXItwO4E4APj5l
uvirhwntYOae4tuxEVoqr2pG/jMt0PjFcWMZ3zWH60jukuhF8zsog/X9w+yV7Gz6
9gr9xWL7KFD3oLeWWOvAr4o1l1KKuNcj4JjC2tq8+iQilm6Jr9Hlj4hL6tpAb/cw
PAdb6r9lHuMpOo5JctygGerQusNidRjcp1oYQYBWHLl6p+jMp5qqFvFfwZoREFRR
u/U0wGxtQOQEcAhs62D2vJnAj3lKHy0QDGxDqvv4vEyGjmk2X/W1A5cq96dLTWaC
wA8rYpEGwO/PZnB+TZ376idScp3zFudbEI5hR7cNml8kTitUny/IovU6cf9x41j/
KgNIJsx0wvHbe/zDlt9/Kz7q/2HwvCNzX07lC65tVOf0G7W5JLeNzEWCne1vSLAK
wcKBYcFE6soaGESRAF5Ue9Z0MFuuIQl8DxiQVf/r+fVU+xp/qFYZRQrRieF76XCU
972MB0AenQ9OTDk468BzE6U2Acpr/URedXsGw8mGOJZ37Jmwgc1puFfkfUlmvHn5
EO9wntcQsyWO0nD6vdSubBQSDacSbkX23BRJbnnHJdFSjN43Vnx2U+tgDrIGW+ef
iAdoSMzaZhg70fnxjC3WEb3Sw3oD+7A5mkYzL61y2NFkTzX2RwMRABGzP6a4g65F
tp3sZ2FHJh581GwI9T0t0JQ+y4FZYwEi5V0hymkOE5n7rV4KjIdIf6qk51NdaZu+
MQDBe15j62n/zJNV0Fnwilj9dM3PwbpG6X/TC4vaWagSjUgXRqyKm3fDDe6bZ5BR
xO4CAUw73saelZZIcaQLhY4bN0zIbA2lhNvdcJXioYTIQf7+GJjLskLQGNHvbhhJ
04qpnZgmR8y43kCAg1SMjQjZgNb/ybR7l0UJ5EBSCUmkfd4Z/Vj3Vl2wgorDo54e
bUFZS7xYHumBAsrGWwtAvSsauYoxgDk/3J5EfSJVvCAcewJFxw/aeiSHgvXjCpVd
OZW3TLCYNI1HvO+ErKwLHEiAYkXexwaum+UuN0PzRGTk71d5esjsDpnSuR32k0jn
tHbmSbs+9GYfRfmynBpBLBAQiXXhJX0wPQmLtcTTuwYCk9+dTpz4YCd3z1sjgd6a
OphgTqyQJlIUPiPXT+PznNaFjFoXDRKaCXkZFlPttUoiaZsA9MEJ/2pqB2HktyAL
7XcRwCN1f5olKs6QGjC7avRZJ61wls1seQmYYeb4ZAtt3zWNEOW36gF1O84QI9o0
ymcACVE6bWFmVruJLlqBdC6jVO0spr60ukNS9R5n7XbcqnJPwI+Uf6EuJZqhgLEb
KyGCJphGknyBf5fUPXSRq1BuOXM/fw6yiCd29XMCv7gcaxS81BiZqiW2K6lav7mx
Qy/CGa13oLjqbC1QM/rc94VTIV0kpwS3hTsFHW/YxpJZlT8IRcoMKzaIK4sHHm7o
JRlZr3DgKg4z+3+g96DH7rAC1tg9cfO9PxUROZgqt+dik3T+zeeAhlueyTgiQZG0
CzjxoO4hO2rIKp3XznQdUYQZ2EV9AYt5l03men/UtkInZywbUwQi5DbyiMNQ2/4m
wUVDdFZLXwrx8TLGfCttQ8DjaV3+INDhng/CZzY6KIopBOc540SbbT/8GxTZ02E9
O+WbCDEE+Dpjj6mt2pS5NkAnnxQPJi0qlbvAwdRCeRnENoLkfMK6dLIY066qKFCH
3SxP2DGSSfuXtvkaHDSeWUhEZdVXTv7xMq8E0i8z14JCuaoyZ70TpeFjpafESNZ3
VwTwtCp9ja9I2XaPp+emuZb3kMtMSIalxCzm7PdUN/WZXC61uIzxVBhMcAEcVAGz
DkKcPRcDz+QmE6Ph+h4FGzvO/tTLzYQ6W2X78itzXyTC3UOEH1DaV+u5mbS36Gmc
cHvU50pPvAh6VhW7kaZc7zMy4R2oY8sLcKQHBVqDWsUahwrMlVDAb1B0ywR7J3PZ
fgg8jKnyG9iy50Oo/c6kXoL0HOZ15FHrUwBOvyMDOCkKV1vUNceYTWAjKFUhLowF
P7tlNJ76UNwVJiVD3HTgQuejibIj4hkBrhh8rwhzC1omdIAT4jYzdR0zfXsvm0Iz
2ySsM+Oop3Zww4HWNwH2y52HPrWvYrPay8/7EISwmh9LM9b4/pJpbO0mGtuEj9d7
LA4WT7ZhIShMq/5vqsteArVmYdFRcwjgrRhkzgeMM1h+ZVvQNhjr+fxWL3vaJGw8
s8HQAJOumamNqGOuKKhBajxzSPUR9F4Fi5xLh4gau7pqs4b7+vMZYUvGB9iJjbdZ
ht0pNxELmPxGKDnBJPCIibCOnlfLF3iIeGk/t3u7EvM0mzJDC8okTYeweE3aeZoD
bzK+o3/Q5JZuqDkFVQr9keMYj2RBGp7/nYv3v8iq8YxP4LO+ol68ui/NrjwGybeS
14L91vPfW2YD9RBcjBiX4j5ucAQS2AovYg9UEoevnEoLPwae0pFk9TiqLmVfQwr7
Qpm+bTCiI/SNa9J9ovGzJSxKjBxlW/j0F/4VvbPXkWxhlpuABmZGyHFJ6ewPxlRm
z/bcNIPpyM/W52ISTk9F5njCNy1HTFZJI7ZwFHC615ZuqojZql0ywiPsj0/lWPY0
6ZcCrfhekCEbseQL9Qs1YM9OQ7lgIQfJGgMYER2lYjKprveSMwV8kfkIRw6D7o5L
s3TqcjBOf4eg/oh5/KzxUNvds5YRZJQ2Ey5D7uNiATH/HW/sKHA90SmwJ6C3MdXb
ZtWLHe3bQ4eHvD1qI3Rq/MclXpT3HvQaH7ngbQCxIdWMNn21XLc5UqQNV4R+eZ+A
wPJoHWOVGXNtX4eQn2vV31iG2rWUOA1TWAk5/ctBM7verGrt1wZzxG5LA8tIBiVq
U+/b5fa2nMS5xBUqOPB0Clt24Pubcj8E6XMbtTSPu+w0399QqQfI2BPckwNDYFYs
ojiQCAUbhbskJqmpx+SqNW+Iee9lrITfQ+vcqSjZchHiV8+69ef+FXH9tcuwrq1C
jeBONO8q1RcD9qwx0uWKeTb17pkj/mBYf/VecN73DOtHmGZf8d5CH4kFc11DW6Q/
5ArfBdjRWl+RrykblrqvXYDgrKwg6jpTg+Fa1oWu87Qu9TmCk01b/Rn74yCrzYZl
LXE0y8jWKi/Zm/D5zd7fqpp2zM+VYTi0eesagnXqsZ8PBdTIO9eIZLYGpG/CzPcE
fLvMt5zbi8oRHiW/tzjrbLskl6xqtmCsZDwGBe0Msa6wW0R53JyxCHEoV7PhRoSl
P0H28oG9AEF2yyReJa8ZKdi9WX1Bb2emkuCEMma0Alp5j8c8c4mItZ9ikXgJoFO0
cAwOlaUWNd4BylOpcQFG6xtWy82xsrrJVTkYZqefE0dn8r4qLcrAgpbYbF/aYKNU
+qBLOQZz0P6Qc9Lqp5Hlbt7VT7AM8vbL8IN7CyjuSS1Y7abR/u+7khW65FW4aDBh
ZM1r3PNyI39MzqmAmjglCbHNwIU/1wlw7IubZ42Eurz+nehZN4REOPHPqKLd2VND
js51MrfBUYRs2GTKqPocZGkzynp+QkRKSyflh+PaKAlB6loa3Ij6NeBilWXeecFZ
WDLz8Iy3WI3qux05kgRGd8yAL08rvNQdNxA6J5LpgU8pKKaL4x9ZYCrQspsV6meW
68/tKdfl3HqOf90sgBt6XEjtqAojS6vlvxIuG61QEop3Qk0P5Ll8+X/4gpa/sAfF
hXh0gDu3Hjbn2ndI3d0zVY4FjChw2jZmmo6OWz1u2wKVwwRtru6+gu8DO1nwd9pa
aO92Qw9HrGHlWrwB0lnt2BfAldbM2NbAvaokm+7aH9VSOW0EyeJajjU+0DHckUIh
oXKeulYDzqXwjyMkjBT7HtEw8d9XwygT6rvLkxEZ3UkzyoATqsFFOSJ+teKCY+Ch
Ua6eaksQ7bSGWahhkSLQie5U55VziWsFa0XJHWXwvvXcj66m8daKmqYe4LI+if4q
PMLFYeOhBxkn7WMHCqkdr5PRGMjxF0qb866Sm96zZpI75PXNAMNt6w5OvAeqbvxn
IyNccBSuxgu9L4vQ08BuCDGyQU73loY7+kvqZDay7wmGevLq64kOG5ZBLZMSWj2r
DkaewXvc9/IfwwfhTcOxMonBXhHYS+hAWE1aRe7EshS7UYjrjRPfhcdZgCDu58g8
JkF75/aartxMe1juipWvr02DGBlkoXoaUc9Ro60sv6QOjwfj8NpeQwFVu0lv4UDB
6cfQ+3dCL83XDunFnKj0ASb04nrk7Y25IwY7njmBmo7aMDE4a2Ujq2OtsztnT5D8
OArLcrDskN7EG6OihSY4K7GpIsuH+KgoGKk3xpihwrEOgdgnxDeFGv5W+ZWkftnn
NH+GFz07XyPFOTPOZ5zX3YmHT2BOzpylzFEUSwbUJavO91T03zs+GG6yDifXqyY8
VojsInCXng7nzj50K/D8OR8fal37FHTgLjKUkw0+Vqz2XwMRTHewAZXyp8qw0uPJ
ge66gZolma1baIgMe1v1j5hkQuLNRm153xaz6PTbsSobYEJYZp6AhiYaeyfHD7BE
2TiURyXQPa8OYxPeiMr/dU9hvmfD+6bg6+vxu+5iDOinRas8OuAPTRh+e0H47lzw
du8mlqBNmeiW/3Xewmr+pN7Jscz7EgmaRbCVe/8AR/b1dkjCCBatuqp1fGLfuobv
bywucQzgiCHmfsOSjdkOLfCGms7op74sJ9AdahX87tzC5dbvZLS2cQnW2mIKGrqF
GOEKTq86LgpeiU+WZRuVI2J4ChNYumI8ZK+i6Q7UL/YpG5LkhbJG4Pr9uB70uQ9W
m19SIL+JG5ni6e2yO8it1BXthwelQvkATUsxzZKiIWPiPsQ6iCw4cTUabBWK9g17
4ACfiiMEwGNsr34qx1Edlh4JG+QnAfAJMdkNyjIo/1RdU8eXaH6uP8DOQiqpn+re
vQbtMnk8kqhy1kvcMFpE6e6uLvu6p0+AxySAjt4+wKdXAD5NIWQAjZDbRl9QjSaW
0MZfzkQvyrX0bhiRb/wMMPN6EQ7qpNt9YGh+hwXfAPgMMS1D6M4ZGRBMzWvjHttP
o7jNKvLCO4XtXEI9Wj7b37DwpO6I7+Z6dSiHHo1HExYAf4Tzl06YCeWszuSjiZ3q
7Ey0ZCYsa2ODISlE4E4/WZTEuUnd+yapdtBJHeXL9jiP45xT0fGYteZgOieJd2gA
chRKOhyCGA3ZBdig5DlFxJPyO2QcLMdFUmwbtY924W0fSzVLqPvI7IXNWed7Wfoo
pI+71J5/1a6ZKS8DKVhyXNrVcFg4bRHyw1WNVwwJgArP9MDZt8OSurlm2ap0+0xc
Cj0fAvui1vdKPMLZhM3CsKtIAvKGHNarxj36UpLV8by3iKFCoxyi4kFjIlrDf5XA
HUMBUDpffLi/pboYSky2VgKTXjdAjHi07crzt44vDD0V2O8JchhzIComj2kCnnFm
qiDTrY74dBfHz0MSFupsm9AZRR/VPnGmUo+drmexU/97rd+tOwY8gkdISbEkLlWL
UW1eRUu3+ECWQhLJYxhN19o7wvCKRIAyX0+wxYNLO4JGmTXQAa+cUPwHCVJAWl6s
njQ/ZapoVYWuFILl+A7/3mTtIONxRubf16nDYgS9pE9JqzHnY97nMqtsKFHTBeGo
RiWQ5Jh0OKRb5S7Z9qItKF11cNV01mB0wWW+15Uz4hWfkdRSFr8egALLykBv2hqS
zIyUAnHAOFPFM/yBhTg9rBE3AEXs8j13Ex97Ir3OpGWFxw2fA8jKWQcedLpbotTU
NKIEAcvSKRWRxVgF0ggMP8gRm1lQmGNzofl8wKzTOAFfvVXMmnnJ4MIqwi3L/9Af
qjSJJrZljXZnHzoaDdFaaYhSElxOyp8lXI4I/XkW30tvhQBfyh0afbRE6Lx1LMwF
sXm5I45qS25Qzgiis+Rxku//L0tepSjZuajtSb5lUOi03cxEag3JJ6PyK02VTsd2
VAtgZtoUFBekl4JCc9qeFs5E9tcEnvAS5d/YC9da5PFfux6gUJ3aeFcK9dKZewdR
7YKenrlqdfqGRgbBsnzhAj+hhYZ3TZrGtkP3ljJ3b+d6mWSggELHY2Ko0zpCbxm7
2ifv4yBCAHEIrjUALtxrDPzLuX74t2xACb4phvO32/jX/uMTYs63IgCFwxkDje8J
t9IZMkFdzWhrs+AssAm64gtC2ZMkRoU2goLFC+J8Scqh7QbzywjLiTgZ3lxyR7Rb
46j65D184OnnA3L35qsICs13JVKNsbUsLewoVDoKPK/jo9yLosJkXSPnXutT/G7v
wJRk4UydlNcLjghoxb71G3U+pFrlekb5/oe+vw561QnIYqK0odOsjV6FZJmujAl7
/PowzUDzTIvcXAxiODEFRCIHyu5uES7qlEAdGqGYcGmI2uZcfuqM7P+6oK2uxLng
2ory751WDB3n56RBRJOnP4wxJKONt98ZIjamz0i2+yzT9bXdSECXbYYFsFGFCFLS
WobU2/ucrMfr/zN2rX7oscF9g/o91mQTsC9F06WMDDgO48e3waIx0OXUxlGw2oUh
gxyqi2dKr1yfjzVK2C9CeC/GrmSQZy1ye6GCTrw50D1VZrp1Vg8RdmTh953aR1Wx
EXKYbd5/nG6OnDkA8O/gfz45BS5hd1gPWFMWThcUFCO64bBVt0siLtj13B5vhJpm
6y58cTzD2ZglUJd7XKe1IEP15ldnudJovsultUwPtAbZ9FBVcQZFtuDj1Sy0SXXG
JaFI8I+xfhpMMSVGNchvIa77gtgG9nf6sc/FwYkAmHxnJbiaAnVywg47uZ38jHYv
4F9ADnYPPYtPdwYDN2GkPEvHHJSZmX3/IqPpoazdU/phpCBJIPMEOUEnI81RzMa2
4K4TlOZF1Lnny20VuIcleQZem2qBBB36ThViI8yHiU7AbdO8DX7JQkoOfttVCd7O
LkuEGwE+2Mm8Y+hgVWiM8CYaHq2pUCZAZbVz0/WDHcGtyBmFDwnJUAp/JBGWTsJE
pk6LbFHrhN0yZbDKVTRwguLDzUtlkX/LDgjHmw7FKA/HIcfdH08V5iRRYCJBuAog
g9QQeepZnGaafPNCgF+CDILjsXks9oJFp/39/7rwLrVn3ae2VKWDwapCN/LoPI4V
A3n2AMg85fPCr8bAYHollNEJmxLxIMWzCqNrKTiYsORE8vDT0KmCK4uG87AFsojN
ifbGG7jSdsAK5Dqikj5PqgrTudHjINPdVQJazzyCiya0U3gz/DNLyCF3pFN9AZTl
amwSwSsdqGxDjGDZt1/AoQeVKER8H+2m9MwaLkk+FxlNqq2K47/EoDaJKaDLyDN2
x4eMnF273RT07PAcaFymnwbLDViQeF7rmWTvtYgcrcTiKBkG+SXzmP/e2uMGghSp
qWSh85GPMKVoMM4CGONRWZ4xJV5tEQsewnha+paFoIzRU6gEmRfVlmYB0+3DW1l/
gxyShMn5HjWCl47w4ZHCvD16bVnWegYQtjtP/ja8f96WJG4Wuusjijh/+XZe38SD
4BIHqzDi7v1p/HKRiIOaLGetz127hwDdpZXZyYHkr1Nhh8et9WY6G+5U+cpehU5k
LjAIMOviISh9mQW/pu351mU5OJXlSTGr5AefsPn+my51APF4CIoHn27pnwMqYMkM
AF9lbACNYMpatEETbTe2IThtITXBbP2ATmaTBxk8MfT6tem6UYxPyq3mJJP+nsue
XWFBxG8vUjvGgJE/rUsgOW1eY6lxvCmVLAp+g5k+q4NLA1wnCDRo+lPA2yN7Ut09
bSRvlckp00Vt4ogxgK6cuSk5HcqpzFtvyvN7zDwiZ4AViHZf+c09Y+elOW00Xk1n
Nt3KW+IX9U1TljUwbKTMMj5+rRHbIVq8o9iEF0j3k7sJBdRbfphoH8nZwpnzjMWu
blaf7VgYEWkLrNWLgsApFSZeHvTjmPXWxR9hTaCFCGf8YBncYrvxA+7UUdrykxCn
IdwU/zbX7EU0YtBo9d3B3AmR3okc1GhDG1Em07UM+HYr35UZwgfoXmArYOTjb0ke
Au0mc0K53fwkpXqEDA82locH1LOBf97NchOUC5exuNAXXWJmXTimrrlUvomH5crd
3S1y31TcvlwhAFMQZ7UGB/CM+TofddGybjXy29mIq3x+kXiP/aesKm5H+bYDXbKI
qCurpZmBuz7dU2fKn1ERxMgcRpwSMZC6rFsaUbglU2YZo+ZkzH2L+QqmAJNrXKi1
Ce8lIbqnT687iFOiIaj9prYTEb8Rt9o0wf8JPkeQRPgOxYlGqKonvnSwYVWtJb0k
49g1Tik/D1J3bjTNJ9GLY/qGjF3sVaaGyDDdpWFWEc01WrP41Mlm90jtXkYMCPzp
GSagsf4DmaWjUhYs/+Gg/NsxEBsqwhJwWl/x5KvGz729RIKs5FPvyfA0A4/XWP1v
FElKQMtS2Y9OZh0+ETCShrwgADyGOtu//GT5G93OELmPGgLMBw/flSxLKm2O8nfE
VihOYE/efZAyhZjquyPSckgvrYxUSL1Dme8lcuPS6FXwF9Ntbxc4AHv+Qn77Ywir
5YLkHsfaxKlL26uD/sb9aobSyJ/6NH8Vh5YrLSEHUeOKN6u0nhAdGr4LSp/8kmfx
BU4FKwc0WZ7/5DEQ69sqNDbW64dwFnIV2/ohT7bpMHTeoccfCmlO7TNkocIe7eMw
fpuNvbYKKU5HxFtyzThEKFevr/cwdM/wwzmx2ybCsXwGWQ7ff0lEb3O96Q0R7QlQ
JwzdopsW5nuVIQAxflav9VN6qeO6jsKK02SqEYxfgm56t3skYgd4iDp2Sxz0Rcg9
nzyV1q/fWjx1dDzHasgcwthXvBZ7Kk3gFkTFTyA3RHek+BSlbNgkYvcRFDTQa11R
yxIcV8xS1aXmHoctjGLDE2ZGpwhIagTFVsTamS5Lrb9RqZALZmTy/e96gOD84i2c
Z75Z0ET96EcXid8p2di/fbzyvFWpsy2npmFp9IimlPoYm3+oNg6ZDGnNw/Jm4F8I
+hdJqBm7mXeoPUibhCXKI2TSUF4/me3EXqska5HXrYcnvGCto8qfKmjvpf+maXxe
QAaT0EleIEOBvx2B6fjX0CcW7pGuZGyt7++5bbkElKGH3MpC+UhBk+nRoHnp1UlQ
tHZ685bqPxuTJt6Kjx9+eu55RMFXvPDu7mp0zyudrfqE13264qywfqsmlIdw6iBL
NIl/KyYoFoZL8RcVfbK5rLIxNHih2LqtASDeN6tA0mju65/hynBPl7+YoSYc7773
bnjYaXg67zFenXa3NnSOqv9IdUJe87409Tb6W+ZXv5FupifWn7HEaK9SAlek6p7j
jIZYPkMXUzJ5MtD95Ue9JI9TfvYilKBfZcCJ9d98qc5MIh2lOLlO6u/HzUlpmDYz
FTqoR7oQkbIZ54WHzYFqKzvsos3PQg+w9STAo5oCT5aVsJVF+CA0Pr/EooQu3bMz
NCM6t17TsbroVvDcEoivgrTQcTGuDqLQDY13n1MoCuiaLtCxjvLNtNYc+VeBhR6x
FqUmw6Mb9EfRQxXGZ8IuAJ2342AkLz05TS5EgfjpzdgAYTbaFXUrEQPQ5INiFR56
EXw7j8VdPXsnzDqCcRX59f3U6tzGAIJqQ8aPAMcGwG1/x/MvYPgmiHdl4F4snQxF
s0V1HT32QIEaZJUWi4uPO9fikUj9pIjpePKMVl2yuo9O08Z4MnRvzx46lNbp9omG
rgWYbIQqCZfko+nrU4i1cIvVjpekHexxLG1inyc5fR8K7nubVmQuT7kDg/tvtGrE
sMRDhuzUkvrYT3O93P4Bc8Dmeo4z3GP1zuA1Dsv7LKEQVMFVM+7EeuXHzSzwCRw/
bEoJikKgkbVoCIIyMwVoc52AOwJ7ElyUAlksbj1pqnWWk3CI6AvJX9wXVi4JDfXE
bH7cZwUM6gpSrcsXIAeSoN6lLeCZAevlSxGGQGSxdvel1vzMhF3cMPWgJiDndDUM
UjIDstJ7fPCHOOeEakt3o17RWd61ypgb0/yLS/IG6HisBBRiIGMHnaB+lfbNFkW8
DuklhtCQ03Ljn2JaEreSqpN2sNJU+gljFbFz001gyXC/NLjLjxNgm1rGlbSMxoJT
xZGYLqZvYv3DO+/hXltLD0FVllQbKces9ao/lKVYM4W1kjl541GorMaHfejspCVQ
uDuFiORR6DQCTAWmziSiEvSVAdDofwWV5o0+c5cAfFIHa77233/kNPHYTCz8fXvA
4mvuoo3q94RIbUYD1JQuQlZnBoruDP8DIrh6WlBLFq0fdo3WZ830rBRQ+jLnR9wi
1vQzpu1vSAYq+tM6OuqCd7qzRHU75EzIJU1dUJ12hKkxqNW7K9CCxA6m1dM8vMod
KwHn91QXqyweg1oqD9C28ybCGPBclk730wdbITU2vUAKzirn49SBCWJa6lVnKTBK
Ob2yIwl24C+ZPutmlWePWU3Bf/pOcT/4IOWP/MrKs5PYZ3ElMpcvYeYHElG9RkP9
YzpOI1qrKodcsM+FS3vcVIJYP9ZzKyte+h0/Fg2foIrwiomKDxUie5D8ZUbckzid
H1l+jriSKRfxIWERC3fOu9FdrlYPBf4ZDrUfL6ryw7lZaCQwmK1m5zwd6gzhSuFx
Vn4p6odtRZOrJPKWX43VLIrspiY7xSXbxE36veUaxGJsHzlAqH6gAGguRzP7ao9t
5oeg/WfePO5f3Z5VEBQ75N3JEmhyK0OiaVr7fV5tP3F7YiiYIq6SpeNRxjxyLwvZ
20zTV4/5r+zyuu/VnySMzRq76QIjTGIAAgGOUoUDymtzU5rgoqITQCZAhQLgtNfL
QY9kTuXZ7Y2E+HNKTeKQuN4Wd/ZRVHhMlR0E6snuyN6hoWUotpWkrQveeOPde3bp
q8zee/LhGnp3RJX3/9L0sezO8Eo4lihxoZe5D8y3k3QFSAb1aAIkQIz/64nSR8//
XOnpcnFrxq8FeD7HbxBOnF5BQaQ7S4vq3Uq/nTEa8QfuERIVLKVIWASUlcAr7/Ke
n2+IR52RWlJCTIPiAfXnC/IeZiC/kNm32I/mip3XzLs1kfm4wBix9gI21OwW7ABo
ycPUs/mPBTttozTpwV5lpAzZgBuuCNAGR4NN3xdocwI7mxl7Xg3ouDJvGSpWr8uR
wgGFIotV8i0qsofUOg7oYVBa8wrzUPVPNNfSfHvqTkL8OOvFMrwD2HJ9HQicwGHs
5MdFZJlwGJnN7dNnlCio6mhcv/QX90SZw4eGmqf1AzWMAmIMn8UgpyLBefJimjS+
kVjBCWU3Vg31xFmNmzPJ15NLZ/Gm44AtLou1al65BMfVeiWVnWM1SXRA4Xk9BNd5
xc9kkMnbsrztQFvQFLcQlwqHZrzN1qfEs0UH2zh55CGr+jYCFLv3r+CG/BAI80w6
iL4RhLbN0O9+UqvjaOkg2SZt7YEoHEsBm73WIgUebGQ13JPWtBHlGBiSu+7QuO1t
N9LMWrtxI/dea0P/UHCQ+SOknfXgrfxWZ5xv93lqP/uZNFo0tKmak1jQ911xrdll
ARoBQpu98ldNcDtZ+1byYsYl6wmVL8h3uk0NSLf72a0RFiYJWELKpRXW2b9actCH
KxvnozIu5SkhRZvv+JQCyIJ1WrWDiCqyDb8LPFmJpMuyGhLTcIrL0cXlYC57HmlR
2oJvm2FKJoTXu9wT4bEHpeCuWp0YI91GMRG6P7dKQTSZR0aFjI0onSvjhotMFKzz
mTklDVQnWb9b67XrrasOpgph3llUNdChVe+hTMQEeQRi8ZyOSkkwSUoCM5i3CD/1
i6UO0tYF1+N2yNFXWK28FJBMdTCsoZWcqYX5Ygnr7PejX7ONPIb95boTp4lJTJlf
kp6mHZFe5NoXwXvkJw3T9WViSkyGqSPcwadcJ87iq99MPohzPQegS/lqX/RW4Cb3
oOOyswrVzlsK9r9MWhye9kPTAKchpIXg5WOT3CYykmgBSg3CgZEOU6hnpLpcvDm3
wyEv2uAnN9ft+czm/gwsyL/nOLjCgLiQygct3XYpgIGtHBviImTBqgopaJKI7OOl
ulEhwoEPYGR/GG9ONKnflwJgLOjzD9oaksHBOdhbnZPZ5E5i4HsmSdqTvAnpz83B
hHA2Jei1SgSs09rdrQDYrNhewKG1pU4rskEuyyDtU5Sn1GjTu3a35mSMQAlewxBX
z9emC4IFohUJKFSL2ZWb4SV3I0aDgRQr7O0/QGRgQN+SVAXjVfbARdk3uShdEk6+
Yo04mTejMjQdqlzmdTv4O3IhnXradz/YcSGKZQGozbU863jCTAIQoSET5A9IDYCH
BHQoQAWUYKFmdmfYafgcyhirWAU28Ys+oQuL0LrAGV4yUExaOy9Yf8jByP7a/Hs8
/kfABSb6df2BWFHuNSdCkhDma9OvLIeYRrTDhw58cwZM2AozNFZ29NwxcNbUzxiL
CS3bEsr0ut3Lg8COUF8az1VdkeO6yZnrNNKP8Ydp0mwrExhrTPAn+xbLqgjbWXgQ
+w9Sm6EMBToUDmRMDXt5ORGMK5v6KLHyjLLOTkFwQ6QxHEySCvdBHxQClgARwl3i
cHTwtFTDimdeTI+4WUUrifiamZW06+CCT8mXax3oQkvKCW+/NIrU/Coh7JUqxEZg
KgPfSoZeylhCq36r7HjLhpMUWPzbLK5xOhK+YnQgBvGypXXd8cE5PU07pxOK0y9j
7j6Rj/VbaL+530i4mZLEuV6cExK/hh+kKX2bK/GtWjBkDDxSGt4RkQ8Lr38XxiQS
jo6WE7cMwex4/GIjcoOprfX8ZAfMxSHKS125oTShZGFzk/h/seo7/c1d4YGn4d+7
YdAUj8V2f0sKh1Y4dvQnMp0w3CfHZlCbtDTL/iIhR6RgKVTLfWzMVdw/v+PNZVQQ
a4hc3EiPJ2MYAPug/2ao5pGWRemJ2vCsPtxzCWezuToudYoq1nHDWVIUL3ig3/9O
H2CGdsLn5AHMuw+empWHNpI5ZfnzOIEci09uw6q00/zLXDY84wkmW/E2xDYfFGBl
Two1+zz7yaGEbOWaNyVuTHHhRx/mV5WwfdJh5Px773lMcNTfgRSIDxesxv7TDVrO
Q/hdA84MzA70jZ7Uki2bAKce64EbLWgXj/qXSboMiO3mFsFngjhHSDcOhCCLhtra
k4RiSWeNibpPUCMYEr4O+iz7wMRolI6J18/AixQurBZZJAV6B1nd2rv6JRgJeEVi
CHGta+zutWqqJl8T+ZsUF5Ojnucqa73j+v0C5t3i5ltqW7jZE2xQZ69QBR02p5zI
G/tDka0KglP8HXHbPrtxLgoBZLBGfPuwavtZQ6mE51aLq/+YEIA9X8zWlUfB08ZT
/dPY44Ha0q3d9q6/0UMFSm9xI4Alil8OaIzUcuoF5bkTq7U/94doYWG9IWEVTUt+
0BMizJKIut8XLnt+jISxC4HSPA7giCz8W0S5sq5Wi3nNFJqzKuBRbJWjQamqMH6I
0mmoR8GxoFlX96VT3EVIaEe0OVxYmopuNLIqBasxFgx4q9W0A5pFKYpsFcDgRHbP
W18PuKSU/a9TzFgqaOFH7+YLPPmFEUQzRHrK/W8Ye1ELCcI1hc+912CMut1ySVTi
H/9+JpT0Oe6Kx6+f9HcDH3F6wioWlVwUTpWUEiie/A6KnQ0us1CnpiE3RA5fGCBF
cTv/f+ipX/REZBzVF2UNJe4ZTxmg1n//WFUlLQMTSutLrtnNHMyw1mlsodjHjtbn
F2h5mBxym7Lj/21l6Ib/mSlKkYQwX2OvWLu5z5XISlphSJmj+VSDcpCW0tYZMzql
tevbO1FH97fbOneAN6qo9ZFOvgD0xcGDEKau0Fie5Wzy9bb+w34RwdZ42advFMBa
qaXEWtfQtbK/AUWiEJuUBjC1t0zBlCvsJfHlBHCIkc6lNEhdZxQha/3s8Fq5KR84
2s7H39JtKGKrc34MbkhCsp01MoLouif1hz0HhTCGJBsoGGC4VmNIMwD2g2grUjBf
Tk/aKNp9WHymq4n8BC7JWiqlK3g1dEWtc/LdMjEKzDEfq0fB7eHMkvW+0LBq2uEN
NhJ6uX+/DOj+ZZUn+UFR23QrczEBFtg1bAqirOc7hy9sTx+CzSzaRl7eUP1DGS9p
Zrq8zzXj0Cd0gqS5AUtvGQET7YIK6nUtbEn23HKiUYcy7jOaNdw8xCQQJ6/TDNOV
GP5VHe516pabCE/1/tPXac9BQ5mQe9HJIKVgglrRkJjDspVJPKDkJ6N0qbt5e5hC
pkTcj8GOWu/6axMbFaaBby33t/uBhfuN+LAH4sBo3+d3IGBrk2jOVuB40Ya2Hi8x
Mt1uiXYR8WkQbzCitjDLPoS8ffw1qCPBkiDzZKBN4YQHlOXoWHsmwk348I1BzOR2
zBYzQd6qUGldJsZhIwLG/5bya4Rl2WlNKIUObr2Yjr+pkpEO/oro6QBB3D0nHqAm
2caeZUWWwYsHDj6CsIblbOBHCgq86KVu8Ms8K/YaWki+LtNK0wIfAN/tlggPKv5s
lULUHSOv9vmBteRBCWCLNMFW0Rd1CKFWRo7it+DzTbkc+HUvut6BzNKDa7M88zHF
Y2Pax9gJfGpDl+YyhZMwtazgu58/hxitY6Q74EOuMQY3rsJNorGguzOD5ll9hJdn
7ILYZACMhAPrRKfGY67oL+t5BrP23cu3DoTGKlG5B/fPxW20oqS2QTswSiW5Mrus
mu7MhGtvAXwW4Rl1edQUzOROlud8Q5idKVnrP1sr82fWChCne0fn049a8XnnHmVI
wRJpXSJ3LQFKCtYNLsNEz5e4LTCrv6QUbIc+xs4IFQ4STcTPETmQBJn/jlw1ewp9
ZSig3UenUQ2h3ZtoMCa9vN4Bn2FGs/0ifgyFZ8zEggFrIU/pTEcHhb3Gvpb7xGHb
M3UNT3aAD93FCN8U9iaI79iIDkPaZ8w/hOWvTTE5vZAlKzgLD3eHM0rYgnQA106N
QbLMQSLIeM3xEqZsxVSBc5Z/MPHHzTVtQ9m98PorO0dtNYtMykyl62IuD5coa0J9
epMB6ZUiF8YqIxto/tKa0jaibBz1r9QE40mK4ahBEp2ddr7k6tlRQHsve0DVM/uZ
k6sGQjhTCxD8EkineK+sobxPHxa0VyFsR4F5LakfluvSHiPs49sJd4u2lqJ476bf
NIRMZbK+2l9AtQtTIa6c3s2u/WCFv0DUDq9pUbNdKYNIvLVBw9GEeb7kYxkCq84V
VBfEHMehEhM3p2t3Nd0mOg5u2pQUQZ3OowQdEn0wQxXZFgGAnx1x+DQK3uBj7gfn
bD/0lR5cbbmG9HnRNhqTp3HziiD8HVQz4NfDCvqKWqNjAe73oa49/Ylg6ZDHKq7W
9AQIDadphEhXr2KQq19KS4vb9pCaGmdmYghT/bu6YufjJUXUmXkhWlyr25zSyN7j
2KgHPZsZWllU3Ya59spzk4vr8UPVTq0Jb6dzLTeccqhULNTzIzoCEXbRWFdssCqD
dqSdZxv0b0aDtCljbPrBAq9561YQLFB1qGkpY+Npu+SzBPsBpi4rsn4ZNMPNvvp0
SEBsvaZmmm4ld8rQzZASBF9nZ7LqyXVsOaGtaUVo2MhbRuUDDVQYYlDcNrx5Zzhr
BMMFNpSR9joab/wtkkahc/g4jzY0t5jHoGTrfXltAIJdKmK2YpxZt9h8PMH3DlBB
MA8We6udez8hAd3bLeP5GFuUoexQUdwL5OdHxhOD99V+fAbcHg3sXNyYOP5RGOAy
ZkktfnifdOFzW1IaroeuWbDCWB59O/Z1pjI4kEhpdordfvmffakK4jberj2FJYk8
p/NZF4ZLrwq29sgnL8Ps8veCvxMqyQiqo+UOwwjlfMT7hnm6M5k1Hbf9r9dK5PxJ
SVg0tkfIC42Dqu3c6kRQOODVaTlRA0Q+EUGinAmMCsNU1s+mLlRpaBUeFVUMioT8
1d9lABtfJ8b0GaNZYJ/UPO9dMDqrBCcHwtpBfthtgKFF1PWIt0jVlHCvpaBcoXPx
e/I3iSU/7TMqCdX6knJ5YeXSlKxVqATuJGLW+thhNODA1Pfak2HP/wnS/Qu5skD8
H/g/wfz7HnI+8x45bI4pOccoNAoOLPa8fEfrN36RSl249phncRUUJgkcbnNvQ7x6
6Gh2s2LQWrnOVNrwa0q8DsBnBlQPmEjjH0re9EvbtIQCteI10Wg52DHkQK9c4876
TdkM/QbQHKmCwFNG6T2viLiSjTT36xG40/2HOmmRNsmvFuqV70XCU9XCQmBF9YzT
n+pyaBCJJjewvbHNyzHL5IJC0clR28/FXSF8HclJqlOXqo1Zch1vrh4ViUrLj6po
Vpor4nNMtfmit+15Dd/Dgr2CusZFqLY1K0VGo4VYVJmEeqR3N4hoPR+Ov5tBI+tw
3fXEuKmpYC3nyirQXbP1D5tiiv2g1uGX6tbSU8xOVg2GTJIzWVIqZ6+/3aVkJdKb
61XW2cL3LP11lypVXgkk+kBPOkWrGNfT9rZULb/1DSfvVWSqlfk+WYyMj0ZXmcz3
imU2jTQf1aj5e00sRBiGDBAea+Oik5UFQ0GKirYf/5mHtKi3DKTpU1lD388wBuv0
hOZeJqJLLiFnc5IimVsn6u/qphgch8cbejFJbnQ5QSe7+AvVmjyYb6B8glYSQ3Hh
vYDy5aH1EI8xGbtIXO16IWeVLBc5yyufQTt4ytOCUb928D3ZrZa1H93KaKeSLKLT
iuKVuwCFWFvVznYFU6VxGBC2q2RPzPuko03LE5HDtCSe3CQa6WVTKe7NQvIMYxxp
f0oUP1HByuv+2fXAYWLILTYRIvzOHUOiCEBj5mzkzdO52SnrXKbuQzDfR4qEEA7Z
/qMgbx0AyEcFirfHrEVLTTgkP4IJ11Byxlj2/64hd+HXVu1I195q/pSF281UNQWx
m6CzZTv7noQD8NjqQnsH58FK88hZ/+wWUrZJEbVsT7dUVy0q2ydgkJIHI9fZ0p1v
q5Qhbqs+YHuOOC8StykYSFmTXn4kYAXBnlJvwwNIZUSrF8vDH+cVZOVz9Epyf87/
MSXd1Li2QMeuazWdUC40Gf4yFWPILDAivSTGns0mXj1rP0z9qqAy0gcKeDNWziBT
WS/JyeXSnwwmwq4fFB5tfst6lxH6XqEgh2cIsA6HlGclJ5YmgfNG10RRcK6sPdEZ
DXGKouFgqo2/LeLcg9qDrK4gC6eAAxZa2+anzFMm5uWrssqOxWP46x8x7eRBklH/
6X9btDupz3z6ojFHqozb1dX3kSD6vEBrhUUchn9I6eTpHfNyMIC1h3puwuJ8mYZ8
eLS/q5un7VO750rGDohKm+tyQ3OdVBJfIueBbTDrq4arCu34AfNzzLDF/jGUTW3+
srQhfT4oi/px6qvAFQz4+CfG/2z7x8MiQShooipkbnwrFhuHXdJqSp/hN4Vhp8GX
zVGPqBtCufP3X7565GVUR59GlP9bWD/E9E0UDfBKh/xboPuSih/53oknJrLH+p5c
W6TmcVDy2ra6t5rUm9SdGrmATtpHKHrEBb3aj7bpsSyQqxdjGeWTzPCcJ4EfCmOn
ygOby1eIFINVKw0zwWzDYgfVVGR0DALVRWeQxZjq9JCCCR0sJpT/KPGRGATrcPLk
6gx03eFtHduub5vAET8MzAk53TLxHkGNzznfyVcwc61fliYtWYNhVGLwhgQDbR0S
g+agCoQh/fcrD5kmcZMxU9S9h5FjyLsIM5RGk+7vkdIwb0W2OTZtca/vVwN03C7B
IlhzREQGVOPQIyeaC3c+dg7dMDOOp7ynDYu71EjfjJ6OEsM3l0f5/z9Yxx85dDvZ
u8ZXS6GkEzka8yoQxLGvgepBClEB+GIuyTJHg677rYibRl7tUWq5lV8pwCDHOXe7
mfaxJRySvnU8Wuk10588e7iUVDK0iwYdoPZCazrppTV0OtlVqSliMWlhTFavv8R0
FpewafIsqjcLklBzJgFkWz+CUWblbj/2zVoK28CxEdpjj7m9NNRhz4lP4k28+UEp
cSttzYLRHDDp/22U5IiTNpIKjGkrZ7BcX3V0eLisl0m59Moz//HMn+F0bQ5kDvWS
k9rYIK2Z0aJd863ysC3xaZg1M0GbjTFwK2nLi+M8bx9hSCjJ6+0TaDAUUKyOQLQp
ZB6uIOp7E5sw2vwEB6cxbBTS4MPkbFNGJFonPnivX/m5C6el/gdHty7tBwAn7DWJ
ffDePk5llZ993TCBQHYrNFZ84eRJAX4ghhFuft4r3rMkB/1p+P2AePIz4Z22vA0B
cJIqTuvdEbqxsrf18J0+4r9otyeEYqJCG9WoyNr3PCeBQa3ViuzvZjnQ+k45d8nB
bM/VTjY7AUiptYfRmo/ZuMSai0EExIqXLdN6lDC3PS60fSMJXujqAmqW108zDEkp
++dpNS1TaKXiN/kdptDJORkqB36D9WQ8cP7LvM098tOiag10xX97lJ5PYGCYDi7p
hA+1V/8hJKk5qhiikehvQ7+x+Dr84WeUu5UCUDWV8JG+GxYyxR0n9fkHPgqq02Wq
khyMXCDVg5JdCvCVvyhYPnKA6BtiLZiHiyC0NKhSKgCsXuqM3RtWZUGfi5Nh5ePp
T5KHASOF3GMdlaDdWGdSL4SDIbMKO7MjtxrAlDEMU6qGYSl4/yp22jmKw0ktoSmx
cUgVWNqBae7QcWO9Qs7u9ttDZC9FUIhaQzgG74ZMclXYuNmolII8Ri3cyJidSFzb
z9KA8F4P4zNxBGkjyj+rwe5Lq0dfZ07132VDrNjhzUYdiHd+qUkBVxAuYisAeEZh
2+a4BfrZiA8PRZajgYuAioYbSq5Cr55SnYk1qhf+RMzBi8vGwR7dK/EO1EH1GUHN
uhl7BO/09VuM/pQ6gex0+FleokYA4CDf9ZLAo6cQPq3ct6IAF10Z7hycGrg1RqIj
RHpztyXdNYUyCZ7toVhY56rdEDyZRu1RelKBPlt8c4/AM1tDAQZyU5tKgJP5vXUc
V+Z7hVkXksGv9Tp6UU2KzQmMiGWe30lqJBcOEiv2Tt2BB8cBy0shJydT0eZOTTlE
WKSYGh3+bf61GvzHKI96ghjy0V1DZmCUHtpQvXbxfjmkrekHG+eAISd/0tF9PVab
n8lBVfOSiT+PfFBX70PRR2GwwgOfCOWGbJeO0z39SXmzzPweJnT1EQFzcehkJDL3
Nw74XONgGrrPUo+NPj5KHndQqhUEXwLRR7B03TH1y7wLDt11z3QL5zckF0if0b/e
Mao/Y5bTyMY8+vqnOTnslDSseqByWaDpDi15WO++ByvhR/3niASMQcK/nVp56OQW
N5Q6oLx9w+NQCWFQiThcvfywylFoGy5DdWVxcTtqBUEAL9kxCzPrILo/fHDxmZiR
HdX+tb/u9/ULIMuJ4+ByFW/t61gjdTOhIxPs0pmlZ1p4duOtvGmfQs46+/EMhxhq
Lnrt1lygtIQsMF9dzjCviEezswgoJUsA7Bv9qnlyZ4yLcDkdHSKb7M/I5FlVuB7r
KXOpQrfgMO/dNLY94qezt3lQ/zqiRZisS7DsqeFiCcQpkuqTlBqe6hzr9OlAGpNY
HDriA3VGu3VltZlv6mKwUIW8ydWd5m2OMb2GAhzdzyRPNPh+frDM1LpclLZVWvPI
Xxns0k32wag7lyGT3UO13gnA7IsTniQUH33EXz0IY+dF/t4SoWfbjKfTD+jr1Wjs
e4+90oy6coFAAy4N8lDIlDQUIS11E97Ho4tQjki03PFXdtYa01WvmY3G8SsnA6/W
0o4s9kCzuNKEJLI+NXl3pXdMVg/6v2o5lMa5RkOpZuf63AWE8QN1Lv8547iKTXa6
F1FpKGyrGrxMvzzMRxyTm88k7T2Li0lgQclpcoFhTjqGk2XZqGo+uvQxNB/xi4Yk
i57xpxIRMbMypb08hUVLjog81rOqgzeaLgosW8PtbtZsjM2/YaIRGdI6N5KyCyCX
sNal7IwQhANXdqWZ8sCC+x48Z4Luz1yJgNVMB1r7YEsW62EpPOMb/+vO7GUoD00Q
qIq6Pu1LNpX7ZN3Oh6/hpPtBD6JfLwomZhURdigluTkfcC8oIY1SM7JFHSvPLjzx
xudg420CvYaO18Qkf6oIC3G6/bXNnGuW0jzdoa1jX43u8gCkgf1LJh1JMo0qHBZ7
6xlLy2oQ00qeXVoQ1m04Jz/uXFquALQq7RhkNDZCwJEOZWxzgfI+DbhTOeqbNxbN
mli8r+/2uKKTlWPgD/VyDGu8GcU/P+VL2HAEm8D63zFxlFleDBXu5Qm8eu+gp1g0
Wze/hlS/6Otx3D8QERKOob3RJ+s7otjAcqP+VNFS3AdC+41hkOAKVC/c4j2KgfbX
a4KfHOjKO6LEY3cjcpzt4zyqgTv70Fvo7CkBPhJBHt027QPeaXmGg2HaIgiTTBib
27mKSmoW1iVj+vORxO3uqcWc9aizNCZaDYWN1DefnCCH7x66uMrQh8/MNLv/QOi2
uv4V43WoAJaBNM7yuucp9rkoOwTcZQGthqKMeBlG2lvJH9kocgMXu/f7yj+QFgrS
+DYTop03EDvxvB+iwQQGN9eBI676+o2932yIMUxaPtBAj3Pjyt2nkV+RmDoiWy4F
Jj0CKEnEQwCH0QhHbucmySxEUP1/Y3zOZDTb5VTe8RiMzQLp0U2lxsrG6Dv9Gfe8
pMj2aoqcS5FMwGbPU3ndQ1AtwRt9rCPqO0HSQvs+lczzznK5oo7mTnFbjajy2LXl
5aN5Bzd/U+uTr5tmydyjCmiU2yb/4f2HIiEIl1xZXz5FMB0ATVlxO02TDQymJ5QG
nQWs3mCIP+yaBBajUbEvxvCMG4sQI/9kIgptMERH4JEW5m3dpyG7UpykxBcI78C3
a62XOYTK46PQp6zyagBxCs/x7xOkdpB9BVyPxKqs7/Yt7MfblJeIiQcz13WDSI0t
nOQqNxwgVPmzyfAZwLIBi92lBv4+AgpRb9qrudlkYCtpbGvpOfUnLg/jkQn9DJEg
2oWJc4PfPEErmBzOaUFMDtacYeIOkg6vIyq9DMPDPzGjNSDSRaaX0lFQszlAfInW
pBnTkaTU4R9gkC3rnLFk0Tp2b/GQ0KMKMvXCOhJ/Rrjfy43Gem3hLJSaBv4AMMUW
ljCBX0zCv/TERsr8Jo2YRvQ58SXELKJcVVWBNiiFsFLsEVQ9v081rXnmUH02gvOy
bvm6dnUMPPpMsZGi6XLIvaHcLkTsCwX9XkAAgkQgF5EXRQhzME92ETw3amlmpXLc
gfDK3H7BneR6GvQCwE5xxXdO3d2GRe0l7WXcVjGyxXcwRBFlmnWXKXsDPyJXN2s9
VJd/7R+FwOJFTpVSt/T7lhUhfSkq1rcHq3lIQT2R8AoqoQPoMjMFMyh/wmoISwD5
MqSE2MGCkiUY4jsX+KqeZAvmenXNBU/2Le0Dwg+ILw5oHxwt03YTzXyQCr0B3Zl0
YmrkzyZsdYbSIs1QxRnSyWEbsF/2MlnYD1K/pj42ehgOUILs5eAMrmwcp+Ogi6cn
Et4Ra5uzds77fQ3fCGTl515mKA9A0VvYEh7pDdjmXXkoe7mSXsH4wMhDaZnOypKT
Cdc4aMKY6h+5P1tJs9G95Ov6eOF6zkZ5P83CqDxGktG/orHxKZHos4LMMGlALefY
26fFBd3AHBTQfNYkvIUZht7YemPgs/gfDAL5YAyOAHDmotZdArTGGz3g0fvjZOw2
QUKSeo6ro3sRaPF0VEvYVog7IVEvilmqsRQ9mVDWsTGTpVyHo0MgoakqjdGrjleb
4SjwjjCDJITw/g/jyKJ/TD8JeHhwAwNH4YTKMik6uicUm4XrNQ1ZX1OdHyAR7HnI
MZAZ41yPSTc2gvknxOxcQgCJQ317H2ia+I72udZGwAc/yZ/CQGscdcaHHzz6QK5/
u2/lWAIKkqYmbFseUZPyUqtttyzGayEJOJkxI4I27RWroHKOoRZDR6HGOAGruHw7
4prJ+WIeYII59A5FRM53n0JQwOqCxhUtmc+BA3nawEuXjjZpg/eFIWT1rjuBoI72
FzKQ1TT2+UKQL+0GDkvqpipgccKOCRgnSGwn4ENU99Tm/reKhlg2XZS+s80wW5oo
D7p/YZR2wDyiU7BzicsMNEMsTzPyhWyUNVNpJNsSR17n8Xg+xfPEI0AaVVkd/szA
rYev45uaD+36tyvn5qcUiZ0MfQTc8LkM8uw038TOzg/foRomRKgPyvJh4tRkLigg
xVDHdjTWyVZFa94FdTH4FbFlPLTDf2yTsVVznonvETarruDGYvFNYOaDViMN9Zax
e3mUDMmIQINvgYEhJ2Ej+4V2fwFnTvaebldHVTNwrkSrMChhw/q4CXOyZz1riQ1r
x0YcGGSJcV/4dUDLn0slJfKdEOdwiCO1dLnJbkLi1cXi4U2pIJpOKlyoob8ilYdc
pPt8Bjk8gdj60mwOg9i9E03yMLhAzdHiCyghliGeX+qk8N6JXS1ua6zbPuhHU7JR
Nji24DqnX3fDe26D2ucN1745iSwhqfoCOq0yb9Cq1XKiz7j7xXPSDbkk/1YqZ/Kf
tqnTe9+P/aBzwSxpiKa14f1Cgo5Ty8Y/C1iQMfAyggRQfxVfqWBqPAsfroC11zEu
OMAflJSm56Hl6Kif5wmZH/nbL6HRWp7CuDARVewk7INQowG99UXG5mJEqiLJ4jAI
TSNxun000c+nIShdPvkKp9WB9yJN84GGEStGQp85YmeK6JCP7KYAK4/IeY6T5vlY
bWZb3cPgFd/lvUV9wQ3oks9CTx3ncxcWP2GCKmXNgIxTY2eYlB/pukhAaKvByTF1
CFQ3EEtY4iD/SfUfNNZO+U37OuKi2Wkdqa/RTxM5ck4skaxQThTrx8VdQaMyEjFO
BGT9vnx7KiTMp9SnXnGFsaLsg/pY+502bms49X9OnFOV6M6a9vLbUJxsCrbRYfTD
UQOza6YpETEywW0MIT58zdXt7t9efJCdgEWxm38J5FK6s0uiw8qJrKQX9NRex0bf
E9aAbvGOEoqbGPVHjBBtincLad3IlpGthRyD3zLaSXcnlI+9vEVYYHaEhbJ1DcZ8
pOKTRyi4hzXIT6N9+hchy8NZgEaYMn9y7GeoZhJe/XLaPg6yZxt1v8RJUYGEaZQt
mi4lxh5ys9oM26t6KGTW/xZT7gQyodkJZuHafsLk7llQXjQVCO5re1Bk45Fagn4i
bCAEICXy7m/P2BazorUZWWVL5dScN9EoBRVb7x/nhBcrph62vTkgTqDBZc2A4vVx
4z/hS7vf/MUHeP9TcCopqZAIVVRgpc2RVgGEAGOLZZ7AA1RIMvzVCIZCRBJ+o+uG
D0GBOekuHmXS+XSxhIGXBMJtNIOeqbp6GzoOFBE+w3gfgzlevQqdmRETOzLRF3Fq
L72c9o8LXxBiI5rLI8UZZMXb9NhPuXpq6G3+/TWIfAigKy7iQmXrzghxxhEWFbkD
QjCS7gSuefkw03ooXRnuaLeAM9zNkNhyqrrRukkEATpKROHi4TTW07pQc9T4A6dQ
AJIdmVjORyZFMVTwl0PHG3TE3FjxToQ0x06zMXDGKjyD1Y7ZR7wKulifI6hWD3p8
MxvzvkVVeZjbj2ubJLXWEN/JryVM+fb7uS7W2Jo6nP3Zu3M6psRI13VbNLa/KRkf
bAqCM5QBRChws93WY9mjrU0cRkdv/GSxRG4BU0yTNWDywF0/JWSIaNVeHT621HQP
/4DWMwTr9M+1/l6DErkBwpF09QkNL2O9+7JTmKgL05wh5R7pXxjNeu+6R0UVQLyf
ik9Zknv7gFKRvj19Xm8Xx7bnAJImlLye8WCG1T+2DBHxwUcJUL50r4pzIVZJNwKi
UV4Rz3tNeMlwxtPNbS0iECQ6bNCdGRvStZlA6dxxtAZ8u41366j9zmxpZTBG6FXW
ZbPJjzIfP+uN9VJdGBUgmQ+wByAHgfpY4hUSHVWK4nieMtLw9x7INSQn7Gp1o7Uv
Vj9BJg9tRUmV60xNVIj1iI7q3m1OEqU4HYj3D6rb/gO231Oj49/KirtfeL2NQ3PC
wJJ86RNcQKFGKgJdI3EAfarSb/pal7vcVKRYqmKTJAGELDIXLvY9TieL8nmCHnIc
2A4LJRw/sgZb5Ue0LlbeJ3upEhhHYhj3TvhiO4d5XlEhpaQRVADzWnfI5ImZQYXB
bz5vvAci0YxrHtoSJf1co4hGBOLfvIBuKA7SwtD/sR2d0lz8pJvKXSfTNPYtRyad
Vy7dtELo+vczeh9/2PFbxPwtjnilX4i3UiIOJmR5p8gLrOUw5tXuHnwdLgrhQbf+
0mr4Q/3DjstTM2P9ATZVj9sXvddukEcw+qxMiQ8lKXlCYhJAltSCv7REVh4oXxkL
6taE12hEYrAaj+kkeJpb/YVrL/9Fu8Rf4r9BNTCZIgtTPF09StujQ6he57LmRg5G
ZboWeVtvhOLQhUFDA/NU6ddL75wzftZ9Y9TmiBAEQst+k8otZyHO+KkSxWZFGOCq
qzXF0HwFg7XCmqNCLMSuk8tuhr6CYXG0bSGaXa6I9la+vSRvDX4UCH5q3w9WdnUr
RMoUlC+dByjB/98vQKxTg0DWy9Quz9V/a6ZdYE6KXwkDof4fbcPO2LZSxfgEPupK
E6gPqaotYrl8fXpwOackah6oCtzHNjtKmfA1hAB/ZUalYEANVNjY3C+N/2XwEzJ8
XnbBNkFNrxQNlMohvam/Ht9CaldSs2lOi9JbP1+xpRIOWvJL/DDxxF8gUkttuits
MrESWeWni/NmNEm6ONE1rSOagxbxnbFZy9NGp+V/W3FD8joP+6YVMWaNcxRVdJkg
gMDimu/+HC8qmMpC5rO5XS1oLhUGUBDf7Ea03p4SQwo2tPTcZ6ULkyrhpgjoHZw9
YTKONEWQyx/5QnqLFx3JA8stQYDbD1L+NHJOaTN+QM5VRI4ffBSStTy0VXXmhnTt
fV/PKSg9Hoh2dyfr6H1thmXYWb1T/uGrkmbgODhx6X/Y7+qSayyAGqQuNoBZzeOx
dkjewiyi87Z0S0+Ve5f0w2xcR8vvNVNmmPg/iVu/u7O9ryBwdnW6D9MOzxEJH92l
GL7VzvOfcwB+HiWsrvxzWlQXvNqR9Zst+JaOtJFeVmMpreP6APDiWayuB/g2Iq3D
G5PIJux6oSE6HHIqqhy93ZeG0CFX+Gbahru5vJIn0aiKvrrBvw/B1MpAMq+z8O31
oVtA8Cf/Nse2SyrNAyyUdsUaDuZNC3qQdAYeCReRZmW/8w6+tGbjpWjG7loy3Kie
k1vyhwenVj4ZpV6isLhgp3tYmzFjuff4677cTs6sb0L+MGvpXuwkZZWN9RaLiMfA
UvGwDVIKN/4fkKfOfd4rVDdRjmX0+pT91CQaaQsTGU0ZUfmwkOIFTh9Q36bjb28k
oFRt/Z+MBNQA4+7MFO0SPdcWpOo+P9M/EHROZGu1yosjge/EcfwSX6rCPpMQ8ieP
qCiKmJfTtjgiRdp/QaFK6Fc77NXSqPuYw7GwngZ11S+101YVaJfwFrKQi2bMKgtJ
kfThKp0r3jHCNE6/9lje6hwbcOuPARyyDtxKW0tjmUUIKuB7GmhHkFgpyt8OcyxE
POKBFoukVbHmZ+KAiPMOr4bu1hN3BM5a7chQ0tP7V0Jtdbq1PXfhUslugK2FUVIO
wboHvSuh/vwOg1Qbba7yHy7IiBDHYOge+7S+0IaReJZ4egLIDoM97YpsED+JzBx0
PbBXpLmpF4BEG8Q/Q4CID+lvBAHs3YPgFgJvQcAvbZ/DfAZvZgR4FM3q/rDk51aj
cwZaBTTymg2Ez6WAMpypoUhmG4KOnULe5ywtP4mDY+ZTQJlVuNUET+jM94Pre1J4
7PzQCLsmYcZF1vw1iXL+TNL1XhEvuPRg5loFFL63fz4F4nfwVESUfqXYXIcY4RgV
xzBZF+fhtg+foTX+54GzoOxaSNQkeBbY3KaJkjBlTPJaxaCkofPhXF6i5yjgODMd
SlaGT6mJB9wHVSgHPorQlA8VswQonHXY6WRgVtdECO4IiwOnVBk2Qc4Uj60p9nuu
3pg32NrplwfXKrrNp2Evq93BjYkUlsXEUW0QrSMmLhYv6ylgAktBBSUYBdZwn6pA
CRbnmS8NdsEIupNLfIoY8vMJUlsTh1D4+Lx8w/CTsxAStlqkOVoCRPXWp735mvDK
nn6TOpOw7FDIhpxuv/5SNT62fivwZDkFUmn/OP8ufOaNvKd0iCTVvPXMbyHlj6CV
nsJoZAQsf2i3gQbfBM8hcAomvttNZbkQEA31VByOtPJuf6XUsnqYJbd2+N1ziC5E
f09P39EKlNfGdtLLROUkhgWN+CO4WUdLG37A2NyHDRFfF7uj+S2daTruq0kJK1GP
TVQIc6jah0HKCLvvOoIAaXUA0pzRXGV73bRPeezQhtGMUHRkY/c+Bn4+nbNH2hgk
rctiQxK1e7/UtR/dvjt9UzCDZJuAOJdxqcKPa4J+NUDi44QMo9YA4+EC+09+Cxlw
/iY4EsxPGAqXLRODLz0vNui2P1KXGokOtFo/3P5yCIs1GcXthlm3+jJkX+f4Ljhu
57IplgKGlepiH28003ATlCU9sWX9wrZWXPlQVLzPImkEQC0RBBe9ZVv6TldeRhiL
N/QqL/NcgVuzkE7A7D7exPRHyF+drOKU4RSVWmQFjJAJ47/WEvzEG2RIVL7grEnW
8qu4thI5e+yaaWEGssWtcKoTCOuqL1JOwnXxiZ/fvq58sACzjQA8+lCeVeY2EZit
UmPdGenQxPDGwby1BLnDXJ02nDZmfTfmfVhrhWnJNpxTvgZG/Ijz7tpep6oI9gQI
FlAoxVsIb77y12IAYTicKhKF58wQhqmj0tRTXtnUJL8VOVdT28WKK5dk0e1mWiX5
bHExO8XKPfvsUK8Ezu+sc+VhvP2mF+xvEz4uddanZ06NORql0xMEytTII8/V8cqd
02dRm7kp7xsDbaqRM6zM1p9Mo5qr/ksHP7DVJOgQ3Rb015KC6+UPdjHq9Ib8kJKJ
QROCKXBjxdFLZx1UQWKxjyccb7hKkJqGel7SCBU3liBwh+KS3eRp9XTjxK9GrU5Y
aaRRJbCZRfw/3+ycFYxinYTxSSoF4/VLE+5NM5LU65Ohb1MNe1Pddc7igfzljl7Z
1sWQO8r+YtkCPnS9HBVLJ34jDcYUAaW7wRhzq2ox5f1ZT9cb+Y43NHcS4d9r+3UB
xugJMpWbTorD7+pnprvNAi6fmgYMmVasTV33l/tAEXJ8uUFxiQXSi81D9lshc115
XBBUpiXk2bMW2wTOthfll6jyCiF05fMh2GF/7LVp8MaSUI3PH2pJM9EG0TkLDwz9
osuuMOjxaK6dMKtxkw5QOzOdL79m0vdWw4xO8XhSH3AsYr3GdxHlJWRR+43N6KbQ
4HQClH0kJ02qn8vYuUCRdFotDTEteAtU8zx+ls0GGjwd9AT8VS+LWn9mAiUObSV+
QvHOHegXgoveH4pSANsekuu4aqzItSeMJq2BX5RmI8erKsKLi8GQFIvuJthB1ql+
zoFNi/l9Ov15n+NLFn6zHvT+uQmRnFNlMLSOjYRhCWwxVuXDW81XYiTTbkvFbPGb
mLJX0UFzk7BNZ19KTOHpBkakouvkIioTeB0AMoy9LrlntdmX7zMRhJ6+dIog3IqC
amVO/u7/ub4poLFw673hvzz4MrG5A+2xPKgHMPuvEnANBidfQf5Ny0rZyicbLxeH
xTS8QL/XoKwkOTry2oT1awf/+XZ0Np8XM1zmD7YPS06eCDs7q/cf17lor/2ZN55S
pFes0nwvlyazKWyEMn5HvjZOOJ0ikcSaFUJwveSyc18pprGypiTydDudymHX+jxm
m8hbHCs1S9ejiMI0u7tbowOjGf9i64s4Sv1QCOqUll6Z0XwD50zWz8yCOQwaa3OP
BxufjB162D5ureJHtUBF+QAHr3WqN3TMyE3Eol/2MrXaDwUYAQ9Lz8uLq+jeCEwN
6WquDJtggaWqXNdLjCeoDAGXHDAIJykiyVv4yzCjafMfET0BjYjFMjka9U3X9mcj
rde4O5YG5UM4llDtPlUJPk3QrF4up2AZo59oQm2cpkUCM0fLFiXKWb5BhURrO6md
sXET8Okh6YMrHDk828UETqvV18/gGYbQcjhOZvdq05XbHRv234js6eB4mqmPlrcZ
XVpTkc5dWG+zCxOteIQu7P6RZGx9CYc1xtQuG6CkQPDMlByMXEQ2uqML0PzVEEo5
vyPRef3edS2eZENN4a80nRQ+jTZhjmfkhIzWpDTYlSE/xlOBoEDqO1ud4u5Gzldc
GwmPgrpGSURmTT2/j4WQ25EVOZThRGnkQNQnP+JEzdUtYDlH7dWyI1GKfshQbTrm
P2L1dXzZg4GD83YEKqPBX3HPOV3d2n2MAPjnnyqGu9i3FADEMCeM20cdXBjZOgYF
oYjPnUvhI4DvalSg6U/oqQRsBkTaOdpK/ywYJ+6mhLZ0cSeP0/fLSIBsTyh2UTkZ
dAHJi0izLF7KlmmVFBhg4h4y+4zgMcrgz4aTCIXJBhzgkRAxa7FJyZStCMAT1umu
mDJBRQ0gfMNzEZ6gwOhD7oo8oUXgxb56KHHwz/tDMB0LPeHSSO0U13nw6Fu3Q1NQ
/Z6Pzk2ugR8EDvZsg16yf3K/iAf8SPvtRwtbppb2HfbhHwApZFt/TfXRYPCG8c+1
tG8eqRdT+1urwv8/Yxs9lhWb7a+VtjxyEvjaAAMjo9h6lT+uy95X+IiJqE41p+To
6OsAj2EnUG0liKzs8JTLWcc5FaSccrPj4Qm3Vf2plGDHNZRA5t6iTRyEUPM3mrS/
0yRvOzj8Dy8LbNqoIe1XxT9cjZHB2PvTF4fB3/XcUcN88CFvyN9+95Gn9QyVvwfu
MkZJ0iyZ+a3UYWX4I1+3iMkQBcyUmat9MstXq5qkli/ftEHqSYp5Y3md6JC0yrGw
w54nhJNKjPsR1LT4vHZFesqezzV65wB9EgKAiM/oDovZxS5sGRJctFwDmEoRpUjR
BKIBVxQcb9DcepWs70ooon7gLq8sjhZqAvTPRhoNYNe6HOChWOjoL3HH2ExFWJem
fJyzL+lykOb310HtstlptWOQqgxUlc6kTSeoj21CDDOoHDJhpI8mUG9sRZXpltxp
Mlilj3mSs8doNkcaYLDvJ0Xnkivj3QYtuQDCCIczlWV+VcVv7B8Qksa3tCOvsq7L
RxqYFSQb4K08RD9kgGOqAEzfofN/YbvY42i331D8LyS1k0h6IPwPbvCdnce9cqsC
+2O+jXcNNNwRTd9HK0Ci7AeMC/3MzvlmaoV0ok90Lcr9fLib0PDpq+TBWSOS6/11
AvYtRR8y4C2vdCPkOh9PBGZ7pf3aDi1gbXD0zhw1oJU715RoOC1QFc6KriWgjcQn
x0jZM0gqOdsF/kPRLJHWG9lynP3s58N6NilQ64ra1RCJ6v65+domBnfvh8BxsOnW
b/xlH4PmYmuMhLn66ALTQfopwM40DpsbWl2/uYdPK9GoGWSx/5Td8/jKoVDqSlbr
uROyCzGDr4PqXUNhmDdPdiqER6xw/MYnPptexbiDMPAFu8ovEn13Vqvgnk6BcyLm
UWsYBxvDooTKHOJEY7OS7oR/oC4YN0z9L9ZZxAIlcGbzeQK5a+I2flj8cTYlqux7
LwO4W3s9xV7FPKev8T81vHUm5x5pH6Ig+732SGI0rJr51E5304breNoObg8yYWz6
6jzg2pclfYwBB17L3EUtznXIJJ8QGsiRk85FFNZJsJmyFTQSPgCVwXob263D8roj
iid5OAJSGcTx2RZvWW3Btt7uhrsmQ1ePD1oSPk3OdyzfMWKIfU2WhYBRd8RpZaBp
QmDwtb5JcwXAo+aaIK9627RdX6s57U4K35nwiVfOf9Fn6Qfk+fU4lXZCgdu1JGoo
/NrmLZrXcYRkZ9x4d+GZMcMaxpgDenGREcyarL0tCeeXbvO73xxILGLOF+aTcBa9
VUIIW3S2Ir3jOabO4y94RrYti1MMHtyVTGrNS8InEQlz5WbPBiBzwoFO2LEAFxds
ryebrfRlut0RCsvCZ6Z0OI5BgLljnvYz7X11jvrmJ3oksusHNm8DG+9ZmpfeuJ8D
Grc2KsAITicNHIYEfMjhNGn113UFiyclnXOi6EZZOgisnm1E3MyFWQRf1caUDCC2
4qnByLf58mxSMhfTjadainw0JI9RLK/AljHuGiYR3jAuC2Bcplzab3DMgGXOqxp+
ecj4Anmfy0jDrV5KfXz9CPC6p9edh3QkOv88I0V7jbgDrjZJFAG8kFhpUe4Se1iI
7ikeOOIuLvUAj60kqu6rwpW46RYlpy1luMd2AOebkt3gjWeh3T6PP+I4f+QBMKs8
rvApo8LsamBqVdncfhNdqZcHVQCsJYO2oC9c9YHqHAbJqbd5m4Noj2DGHwyqQrHU
OTVDOEEaEFEXE/q0sYFcfbHmJntfMdHdSIbgT37TW6q7uJAzrzphwZ0w1P+gzihx
KgyzLeJMCXUyI3vTf5b1GTIfXSdH14z/PqgVVYHXADES1pTTxJESFxFa2vh+QGyB
z3+Z/8Kp2u7h9w5ZIaUMjtcllebrNd+yzJNq6YsA19l5IBOk0VELIjDXLqqWTItS
y11Dqsjf2AIQAwGa1/8HGpPbcFlD62ThzAeehv0nAiR8p04VTyPxJrMSR2B0eykY
pQmSX9BVzskiytoBKIeZQdB3I2YEuIFUxGIrJEejPmRTVEwlkSaKThwDkJBA0BjT
7+v4r6BfJ2YbgxGOg0QVFgjvw4afZvTFy8Ct6ysQ8TMnYfgUt9YXw3vR15zWbKKd
bGFQMhPyBH2IqvEXK7aVSKLyDpoIqVoG+JbzC+VVl3AD4ZwYjY+wVClLyfm8OOqb
2dcejzOaj47lw+fBDu21Y9TzbRlyViHXwhy0wysabIolw9M3plEaAEVysN8aSevE
Rbj81m79TQHt+Sq1v+5E+EWlKvyXT1ZM995UA+4oYSsuQREld+uaeEz23/78wJ75
RHlNPUCqT/Snzy99pAY/NBp6/EHozvMi2i/ACc39vefsQEcytco3nsJopIhiwJgP
CoPmZ+7n5W79Nq5fQHeWE7IO8pT0ZOejCj9QeOSxcMetdykhtKjmUgIEmumakSNT
1XW0svGwMVTnEpR9D5anunsI6Np50hIUNbb0ZYEF+OvwAV7t4eMwdTVt4Jmu0COP
fA9T9IMK2/mLWzBaHFSuI5bC3eNxMoK2GgjSJK88o//TbMhQqkgzYFEWfFuyDd/x
j1FxRCgkpFt4Uk8bUaU8xGeo/j0I/U8Nk1pNsm6Gu82WgWUld+VovfYcVU24GNX3
7AlHNbGt2psZWAIsjLH7s3OgHkU5eghdlmCRBQZ8JzB1KZEHxz8JTRvWh/4IbOfE
FeXkjmhoa1ZoS1GbzfckaUzHGldoKb/4WEhhs6E8To8VtWFtULjzb8DWsuE7+gYQ
Z2p5Zcwtf+FApoPWFalhHsr8InP7MMFJjUh1A1ODIF04pv2tbehhjo+ogCIMc+3W
KXtlpea6BWyqchUkkj2tM/Nw0KpHfUeBzb1HhV6Yt6gWG4bdTMDHdtf8aJdVJP+c
a921IhXrGPRS+TfGG2kCo1rwkMP1nJgMVTesugzvDdoa6D8cS10q4z8U48wA4m6U
es98bkj5ynheINqC/Vchfp+XrBJJr8Uy118q8lA3nR9WUDgcoYgH2KcqSWdMuXjw
OS8iSjZKeR3oP57qny3PAE7nJklfQx1qcZ0gO9EM9dZVGRKR20sipwvoyGk0mOtz
/yzhDJ3FVUD8XByyKqdFjSJmOpwPWV5lbGwnw+g05rZEwGKv3CfPLcNgX6y+cro5
GFHPf95garTAVpniswueAV50/yq7DDVNuJOl3SsLRh9DUpJRMTuM8ANZyDFhNZ/Y
cxY7f2UQmUSg4UjUX7EzjrjLkX7Uf5eNK1beVSiGjLo1dJQa4yBy3htk+J/gKQER
MdiJ0Ln1sYoBVH+Q5SP+7GfXGqaSCzSlurRDuSnEh0xSNF8BNERFqyEUHg9O9STs
n7bC6CkgaXtjGBblQuW6RoJ1h1bKqbkrvHCZzuSQqs8OOGB0KqbOL9pWkKw8lDgX
RfoS4Zsj4QrG4KmdkrXnQNoS12ysoCdSgG4jg7Z5L76hXkPLzWX2+A6DCTBkJ0Pn
kEpHfxwRyZkc89iT8ocuNCE3wqnR0qT3K7mV2RT0izzJcYvosEXNBJxGcj6zuQfo
35rrpCJpbkPh+ltjNYMk90mKtGV7FnDW6UTL7dwbjOQhSodxHXjpYbfqSPC4Xxox
XTuD9ghucB+Z41zij5zqI+JTZnJkVadQpJ3y5UqDp9mLj3ZzWsEUCPmyRh/HUsE1
rT7t81lFCG2C74TOEK4wEkFkTrkC/EPUOVw9lxQ+Q7lRvo3BOM7OQam0Rg4WNM8P
rX6azXbmLw8Iy7sypSs0FDwhIAmcW5YKrGBkspqnclK1EC/G3M0AzrZeP+5Gym05
asFE1gREw3dArU0nk91LIWLzeOVdqGUh77dal9ZbrDrKAGBFLfe99VFrd1pqWSOq
iB8fn+sIr8E/rRpzML9ZP4cVtqLUvmNRDzAh+9rvQi3rDT5qYhvyrmdQVobKUGDa
oy26M+gifrWYyqcerrdghcn2wXiWDSUri5VIAlxcJTenQlVReHASj0PgoNCN9suV
EhJC42VFpn/JcR6qr0srrQBkjLzpNQlH+QmXR9b/8l4wfTEjiGbwqEoFjzrNT0Jk
jfnhDo82s2FvauU/O5drNWQEFKzJtjPKmVMx9tO+8LwRbtgRsNfD2A3YmXZBfKoY
jFFZTsIWFpxUxHDlk7f/DPFv8SP6umOwRhrqcwkq/d6VqEtlHA8KO2DBqadfhbHG
r5yWEHPG7n5cnVGOwp++NW7sXYYdwP7acK2JSKGxx1dW5Lj71FZ2DU5gX50LIRky
vegqKJB3AYagO/NjjR5ACVZvRqQZ6IueA0WjVTG7BvgIi20IU6fCkJQ3Xiquqwie
O36HHWMJJkbvC3tnjKjnZIDEh6j1NIOCiWB8+03rVVj1K4idXU3pZE4QPDqhGbxr
2flB7aeNH/JkYxhLIDh04Ae3Jtqc8EJ3E2OqFynWth5dlWqwLXrLyuNt6Azdz5Cz
w6rsv0FOaraoNRpFQ/0eWaqzSc+6DhRFgHM2bcGlewOtj4PU7iXzEqX5RBVQX12s
FQK8UhE6moaqfwt/Kr2VlPMI3ipBsYReTN4jhDj0jhB/feCg3IdFInC8mQJm7dQI
kMi2rgfegVqq2mcodkXVvt3qkCevrjj2D5eOJReqX+VmLJ9N1Fs545c2IXjQdW7w
xbjRuQyq5teVXJa4aqrxeb7+jRKkFjF0YO8E2jBqSrlrY0FGK/VKX2hFnoExMa+x
dAxjqCtO8e/yGz8/TqJBrnIE8M7f2bxHPzdHoIECFEuha8fFs6Ha+o0YbyxVoO0G
VvZ1Gup3qzgGzPgl7q6kHfMT/2t+qYknKzb1NolY39sfxLez+pFnBI2JQBPX/t0o
qnD6u9C4kAar70/xmMjAVw3clfd4O2ha7s+7qcjl5aCHQjjWpqakQvkXcjro1SR1
KzBD4ZZ7de6CCXNtvo155G9bhbveDn8RBs3U85U91D7fLVnNPgCuaK+h6WhlFLzZ
brXA3mMi4i18wQqICCcA7HH0MUon1dgndGgg4PowzUhBHCIvf5X9w1MRAbEDbgYO
kykvtPnyFjgbU4m2KVvIvdk/B0CeiAci2/i8l709XO3TM4UMKG2I3ddkgrg9zzKn
rSfhnd7QuC43a0O947vLrd/57r0gWXmncwwsCLg0iSxCoDnPLno0Db0Qhwu6moZP
gidflU/qzfZXfu8j0J4uK/9k5G9cf9doftcHSBv9gwSJenOU0A0DMK7BdJhC4NlH
v18/MoNjNa74Z66vd3lbkADI12+PiRsmBIXBWe8ZHW+DarOXgGEHI0cXGQOTSQMf
Ok3czSYnNngOIsU2mIcgtDQNwRNyngIX5Ky8jJHEE81ZKN3kVlhZCT83uN8I9kTa
SmB6/w2xFgSgdlA5rekDo+60+4OMnrWePMYDbCtsqIOSLbrkIvk/MS/3xW3PnplA
4yRX9EGTdq29Klh5yKn/oNzZYbGVdcaR7dZ06YRhHaj84MEpxmzQpYpTx5Yb6jhL
dGTnjJ52cF9FUOcqOD2qJOKoDo2xe8eMyPB9FetiFwNliqYz84nmTufUODeQ2aQ+
seaLx5rXY4AWYGo7ejcYydX80BHkcumJJnryq9OkrFMNC/oXi4IKxH95jY3DDnVe
swTPOZMnDVM0Tqa9FIp+2NusE+nO4tp1mLQI82lmy5J9SXG8RGwhVjktW3EYSKeT
IClFi7a7C2WWZunF0KgIFFP99GC/2VpMNHkjWh0zBacnOWl/Sm0q4gJW+wJu73QT
F9URG/U9YYwHzzOIMKEJSxiRo6VHkWKG2K3FSX8gKrU0dgFVHVTz+k83sMSMb7W3
LYwJkF+gyQijZ4MuZwYSgXsSFIcGYBwxe1cZEn5mLQ8FwETTngw0+tvhCjvgGLja
8+t9go0IRGDCn5wTTA8ih0Kdq+wXebPXHWseowGh85jasmdgvrSxIZ+lURoJsFoN
Xjex7ITmmebDGcbidQdJY0lDGHoPh/aOKbVdsN8YmNsFnLKElJixP2TGhx7avVjN
DJbhmxFtEjzipH4lHMQhCch8JZqtd3e0EwKbSl7vHqff2/wO4CPX3jWLLIMZf/Vf
c8FlSSHGSPoeqfsgrhdNeNIWGArr7l6bHj75X+JnXmFIh3U2r+UMwyQeA/xilJR2
/Hg+c07nClT0DYji6/a18Lbth3DJwz4PaPf83Im7gj5oLKiNiod887ZC6vW40y3V
9LqsrCHe/AZkmyO1OE0RPiqwg4mbvXPh0cy/5yOqE2M+uRQ1YelsuiQ0B00PkvKH
YeXGCEW+82Wb+D4VBWbM1JXw1H857dfGbq8fMiaR+jfmnUUNVwtUZNYNJye7H6Xf
K+J5XDXdRikrru7yN2z72Rq8uxTDUdbmFIzrYD5mXG79LlMrimRbh2uDSNqnIqs1
tXxBt7Q1XlzScXxCgKJk+VJ2MypoTLv28RhJuEYei81VNPLIhkRM6M+9rVrx9Pcn
+3+DXkwoWkszE6c2qc9K/r3Cvj/NUiijgHAnuqRIbZL8yVfCHuleHL5KcfshNd2V
YUjH1F0MfkLICTcQpmQiNwPqUEOzJMju+Eh7w5fH7BiyYxwK2ZUBQJJAkc5KXIt7
9nDQHwfwhkZcycxX3vX7Bt0qXPccyP9n3NJ0b5wSJkDFiaK8PqP7dkNE5iUwJ94f
f94Wh6Y7f8Q/YC9jECBjhOglMq0MOUcpiJNPR/zk0ATN1JaGM4FWwXveWbO27+GS
gWtHhic3YXXZWHpiVzUA3bDgP5ShriJ/y8eRhMaJHU7mD1Yb7VERkWjM6C/Jdx3C
lQ9mzi3AeBFUdukGSXUA2xyo0LG6Z+6/GXYOivewe3+7vs6kKCqU32mBi+aoB4a9
8Z1sqJ/3ERx8Tl48w4YrhEQNRJtkPKJost2lRsXM7ln+wKUbWcfpoEqBkDvkbAuu
sa2QDHos1HUNA42xTREeZRP3LpHTzhKlgZ/HSvfVFvnvQtukIOuQkFLooh/zjniF
SMj7bvPQrGg1VAZkvIA5e+TPOQo85hDhm9f6KI5QN0+Yu/jnPjwsge3WH8VGYsFf
p/1RVbGtwHCNe4MMhfXtxindA9Lsf52AaFtm3cDqPAiA+FtgcintX9QkRYXjbyVx
XboODHgg6B0MfaC7UCEPT5aa/f/5jiGNmYaYrer1aaK998Yy6NvHWzgTXJ0EfH9d
z6PI+jdwdmEbP5royeRmap7J8EvZRPn/C8ljtBB7BlOQAbq4HhUc9IG9L4wDCbL8
IJLO8nKvlhxDs7d2g5fxuBUcHgnZh1KqJuFCQi3fBBUyHK9XMs5dnuKZFoHqcV4q
RNsYu+Gz39/B9WdGwM0oXgV3D8dYJhlgl6uJPpjzIwy5KlgkyTAtaZomPUHaoIZP
H3/E8cttTy3vHAFqO7zi+/dO7Ru5sBcvH+Arbju4zD+NpB4CGlqbW9UUOSL6G0Zn
dG+ZhnzimVpB07sSsVWpfXk2XMfreN2g/oUvhOer/RsiuM8asvDzfNgKc3eb2fqG
7gzA7zGGT3m5vz8v0DQsYiJRYfMPy5jZsSRDer1AlJmWKGvDpNPKDU6a5xuPj1PM
D5c/rg5WV/PFPcB40yqae2TBJso0P7QRCCE4W8xbFAa6JG904L1ZxcxxI0vEsN97
7VQPnr2rqiOWOEcF/J2PfoorMjI+1qvmImmz4hHMCYVkiMTJScvlEVDngSD4wfOi
xfXC0v0dTTMkGpKh7FA9K8u8q6i1XiCXloLfRWcYtW2CF4o8Z97YyQKKXjHe1vGt
OWKWa8C9J3CMIpy2BpEQ7KZP5TLg4FfKEzl/gg3j7ESog1CrUGEMu+TUis+fes8E
lqTiMsZ3CFNAiROaE//rCILecJnS2w/v6NgBFUfiVWnPJMcQgj1rAgk5Uyb/GL21
asLpeUYC/gKmJlOOrUVML3V5dIfKQlLc8Cu7Tuh7dMw8hqN05aPtjP3G/rbUPFDr
jJS1IESkq7tXUr9dU1OYtOJwsrh21CcJHqXoTAVcI46VGu+hTSDhWtiGkHx0zV8x
lgVFZu/FUT2BtM+Lujd5Uj0BUVkl7Zz/gBsnFSHVJJ5sP0Yl7uY7AJd8a6Fs5mQH
8ICqz8W+I4Uy35H9oyOHOhGy6BAkUyLYyDSex++oL1IIX848VZxcW4chale41++x
h/Nvyv1B2JR5vZ/4K02Ucb2HtjhWBfQm5Z9skFZQX6rKuZ7f9ZWrD84vw9t4FcHG
UGhU8EIpV4fFmJddvBf2OHczJXMjTQ4DUoXwp1QJl+p/Ea3XoGjI0iCAaW/Yq02g
sZb+qGCf6mcjc4vPBRJ/UOScoQBsltS8kCccE7A/koE9iDDO2iLRgwiQF+1FcL3j
u5f7dX1ppmucc4rehmFQpF4PUI2pjHu6Lx9GjB+Tikfsz9mW1R674WGTeU7dri7s
jPxt5aetF+v+8EgdN7pUDxsDWagnfm9+4T0vqR/dXC/qy77CaLERVjfqdc9oYbr+
NU9huNZjl84ItDbhKmrmx72HmyDd3vj4B3wS9VezeYZjVkE2BsdG2vn35Oxxv+tz
CmpvijUcSSkfYKqBvUqQ+dkeoo7OUJE724QeIpJu2pBtURRYMRxpCyjnYhCuaGHU
aX0ldb9rwmv+Wh7HDL6ZzIeOXUWd7g3eFLIisrZ0+Q0LfmOo1MJ32yKPqbb4Gv5C
RE3b1LBzdXdOc0kr4dfOH0HdhQpY9UrrurUxe799e77yONXn7VzTOAMIVp3RCbPZ
L7I54h3aFDmXbmCp73meIx76Xz0Nql5ZmMRsyEmfJVfzyBOItROg1A+d0rJ2z9DQ
TF39YuFLcMYSU8ehoKyg54JAcqA+E+BVB/iUptuZI3ufbMjec42iFGB2RUOgHXfF
n3/0ERi5akBGqPYNc2WqNQpGX2YBdkYTO/4BbvhnfVCEuixzPz5F1JeE1r0p/wrR
sLIUqDP34ugs2ZgyOu7l41rjnACxfw+dhAsHcec5JDUbEI1L0RfylSu29QVeS4tu
j4OQRm77Q1BfZAthXgpQAp8m/YVpZ69VxdlbMWeidRYPSXo3FtqHpNRgf8CUOcSq
M5Jq1GZ8+SlVmcpcg8G0vwWqkQYj9aLzLgXQxCW6fIBZcn91GygBotLvvaKkITkj
bSygNTyqFMylbiPcFfHH5uzsA9JoqLSxnoxjZ9nySbP2EcoyCGFNhbG7LOajE8jy
KntgJItUSzzFTgHF+F9TPwxSpP7EO9jnjG62kgf6defMowt3Oa92u9cPjeSqtnqD
gwAi2ksLnCjgSLbdN7QToH/RDAaiYYExqI0J16fWe4297PhlIj1w9z5DN4hy7xgD
LFoz9XrEUMYdK2Iol5h37Ego+MJZ8fOVnsC9xcT58YgZMFnyR/4wv0bqtlB0KAyK
sahTSrcGJtJetZM8hs1oTyQ1/LnP1OI6Q7mgeGVRmPJdWzSbVSjmjVF/nTny8MaL
gRTe1lvER1KpQKCL/FSXOvQBciwjAI7jTKIGt4nkD6AhvUI47oqARgcQWTCqhy68
+qiYY3IF/fE9AEj80GA9YjLpdgGL3N8y/bRZODop8ZVfIhwY0QdqbWkeI2e3BTd1
qTExI0XasqKZ7OuBKX8PqQ0D93p20+fdg9WiWBd3LbeSEojhkFKrK8HhpikFqABC
azvnMRKAnUSA3/AW0bDs6fFKxOOj0mntYj84Xys2azWqytQhZoX979w+UZchAX/e
VXOh+SGKSPZIRVCFyb+g9c7LRZ/X9B8YhSLvUaRgC010/0dufVPKg4/xVaRdwUV3
blJNn+t2lOzTf5uYvt+ixMw/35d+XJPJAjZ9GFUpav5Ae4y+vruapT9u/xKR/GHs
jT27NQAopo5GkiMdWs1NvZZpBv98WcZ/7RAfpyo5StMwH1buQ8C1lzIg34kSEC55
tCUDWuc+cHXvGi0y0Jqq3rqc/LgBi6umAnYKGrrCLLvR6apCogkLMT0yksj7A5cD
FZLo4OwRKrS7gMj4sf22Aj3UAPVhe3r/gSidYSeGmhwiIS6GE7/Ee41pJZpKA/LY
o+cEiDWQh/VyNDUyI+XXcIRA8r9y9EgSVx5s8jtX/BZWgC4qtfe+R7y9kaJt03za
bSpDME07NGI3Qw0K3yquuFf67+rUEAKOcVkEeXPxTDPD42UT4b49ix8a4Ysq2uQT
R/XccEHKsKrTrY7ZLZb2jVjCpzqrmJa7Tvd+Ga5mXWCze3mI38TP5oWZzJsYXsCR
bd4JMLmr4IpfHADDiRZmrWh5Nd6u0Wtv11fyPKlra3RTAOT0EAHyf5Gq5/G4hhyk
GDH4bpFkEXlYpWJwDyo4gE3nsd/L+2+VYVNpRoFz0CKPrVFQmfb55us5Wohq9eRH
CSOKYXlm9RS2AkmmUNmlJhYhhbXc2M+zJ6EvT/CgEUctD9xVBQ/+aqiOfLK/w16M
ppQWjoK0i0DCn4132ejPMn/33GYs3NGWvBievT1tKxCcQ3V1Bk7G0N/GTTw8/6s7
4zcK09GsLVa4aZHLyu8iDpqgfx9WMSRRANZuTUkIMsYDNRsbQF+x0thQj+keLayu
0oiBj+OzKdD02mMiYyms0W9Ahozooxp2U6WT9Lu7qG0UesqOd2so9voVCihyq7kC
jE2A6iwcKGPBvU30/nW9+yU6dghKSz+yluqrYC0/0YoZIgRSclGt1kij9GCi1AMw
mDrbAQLUh37ZTa4G7CtjhLGBcPFS3tWzwgdnD3xE73UZ8S5Wi1emcVkFc0ouVa8x
HSv7fAcBQ2RNO8BjwonmQEqIK6x9oMXtV+sfgY5T+r7OmSbWt8qgIZiqRRM+vXpQ
6iKgmvF6GmfLelgYAZtAgOVpwrSWya9+6H/QpSeRezzFxAygOsTi3Oy1KNXuDEMt
+eY8moDY7OISXmPh5uCzADQEYUrbFf8EPVInL5+dIo5MWqkRky0iDTjbGZ+2BG1S
zYm7ypNhd/8ntlrZx2Ntmt9eqEoz0FkYQAAGQnCoZQj0xJICdACtVS9EtcGSKaVg
agTFn/9mq2/7oK9/kt15OpmXnFPqCVptwzzb+/J2nv42pFT6h6XC5XLzv2fhPAUS
CrYs01/Hqz01GotreqJRq/WjOqprzvYLBu49s6StFq5dN9tVLZrfua8RQz9wqQ6b
RTO2bi8SBPTT9CywUzW9dmPR+Jga5hCSmRCj31JfqsPzRuX1dc6Qy4ab7zL/dQLY
Fl0/Y9dshmi3V7Lvh9Yd/iO6S2o8KO2k6ISbsWoaXJfMAST/1JEhHwrtqoI+mpZ5
9YZOOU0ftPe/9mcL1SMGJ9dxOE6vJTAkP0zxKttTjbv6VK2sfepVg6clTW5+byC1
1XGCBXC4tXszbcRDNB2QGe9pjMdRpPIt8ribFP8nU47E5qzWv6Nk8vifQR2wcuog
Y9syaKc7ICqkbL5E1PWYlMZrdi7lLRpwT9BxrjzLRqtaZ7/pNUDHRTbxIdlginjb
glE79GBbczG2v+IqgVMOpA22pSK8G+rAAYAN91KKMIYEL7nD+Tf9hofVxhwPXod6
R6ZoQei6BJAYGSqcjQVcEmtalPb3lrkFBilJrB+tcvsNnp1sEsWOAXqWdiIotK4E
zPf0Q5OwtNi2514Uu11q/PKLmVZjqBUEIegbmCmspA7U6YH6vrYFudt+M8FyStfp
pKn86Bdo0XkXEUC9NjyMmTlowcNq16rVMR4w5ZI76SSlTIJnPOYxnUnZrosMhZUl
DMg9srMLNpItWdYGbqR5wHxLvL20qPbp+lMRa1IGNNjFWs3IOEKn2EfxNJapQoDy
eTWGrBGRQ0Xgb75HrSqmm1nEpJPm+Gk9iem7/m7lLrIhDfdhgWSLA0TZNf7Ano8P
em4UT4vUSzSqHA6wKQzWKvvv1Jq/z9vroZ/V5YTXx2oDJG4NnyrpqvqFlvgkJnzq
t5CkmRSnAd71cNG4YNHrXRSosxozySNKRTRizo8rV+EIezAplOLUNPAif7/35Huz
zSAxmwyd7zTyXpbS9j3qubqEEi+jkfZL5SzAHEjm3chRoqFO75/WqRUuK49tNarU
3So9BTgEYxKad7xUi64O8kXeEIH52eL/OFwATJsZ1gac1MmSnpgV0+Q7SixE3UDx
et8mxGVvfX/tqvz7sf/DLQGl2DfHAzhv2LNBFz61FQa/yEdlyBgB5N+uaHm/e5KF
6bMrdHpa9QhMpJH3EZrRPUZ6wb6ssOhWlQ1TS1ZUGBB38cRXMGhE/6yndzb3bR+X
O+3IeSJctfaaz3aDw+3cisysDzzEv/GtZWqKuaUEoeLaPscR2+nqa8g6HkCGWbZq
aNKaLYMEY8AEafcEiPOz64PT2CSW6YI/CejwLkKGYl0T7VAhJE5ejvC+m97Hq198
EPgklPnyrR4FiX7j9XW6HN/3X2MNvo5famhmnQKjVT5gIIgPfqJrTESouJH2m7W+
7NfrMJll658jxfAug/LDY7XdV98wi9keeOIFX4SvYKnRPSRW466YKy5JzMT9vwNw
Kzc7OmrxzywS6KjVsIMyt3SCCNxbL+DhuNiHxJvWSgO/xI8VdvH0T9U31Qpbusgo
b/Q3Y6VAO44HYo55EZAbc0r13/nZLlHUa0sat3+ctlzH3kUlrm/OqfDYpjivtDlJ
Ab1ZbRPSae9i2NvdZuSFpXIwJvLQi0xbKr6LWF0adnbiIef04DOapcJy1bzG1rkJ
rcUAEa0F29EM0q9TuqRDW96eyP1hCAjRIkpnSvSUH1KLVcxaAlOp6SsUKeEz+RJj
TMo9FU7V/PrqR5jzqapkBXFD/u8cfLKoOr+8pFmQs+TUUPwqsgXfvv9YWBoPqTD1
XtUbp9IVlHbpqc2liIRltQO7Von6E4/hYmU6XVnYunjWXRwtTMeb7wNDFYny8Tbi
r9AyGcFL4Ey53Tc9W/KgiCMI+PHcP4MgOjvfRNMj/BlkV0KB77ZPDUHE/7aPEwMT
E9RUUWgNRqs6GK/q5+vR2m9LqYJ+YXT2Fn06L5glwCk9sChAA77AZ9CPkKrQVKao
qxyz0E4PsCuEOP5oc+fCqYI3uqOzr4awYtr1OZGtLA4mqkUiPNbVug78mY3fynsQ
OgeO0t/vyxWzuQ6TnFpi0hC+m6IG18XMLYX3HX35YV7o53sZE08WGsCPNvyl02Yg
IfI93DlJPk1mX9ajvBf0rWXL17oKB4KM8v/NXU1PjRrGOoDU9XjBOID/oTe7Xe23
Dmteqv5+ai9NibLELdU3Myf/9Zp3F89jFw8ln6UnbuGWhEnBWAvYlfFudiEZyEDN
8fOqmDxAeLXRtT3y8T2TKckonvmGgzs0zRMdh8DAoXOEnMGD8u+PCp3zvN0wFh8z
OopkH9EelHygdJsyHI91TZd0g9y/ov4CAY5vYGMFcxuWVlXSt5I5aLpd78OE0ffh
qEjF4kP5QLCu0NC2PdM9ABnz5/Gvik7pgV7tEhRfFabRU7X3fs8GJb5yAu2pzbNA
+marLZgYfYkBFB3OyCmmehv0Ni5FAp6il+uaZfgRvivF7MCkJnHBI0o+oawbKhZb
6T/XznwX0LWS4TyTDo0MnZnstnZko8ZF+3uuKtWKMyGzKyAj1RuCITYStYaRj8iU
ZR+o+cnoIghfRtzK1fBkaTF55KMLCVxMI9xUOPIe5n6AJ6ZlSXQ7akcLqfyKXiEG
fjYRvhIdG3ubf41qu5Qw+mAG9gOLYyqVG5pPqC98Bx/tfwk6GremKKkXaS0l6xHJ
87PrZLs8VlaiQZFo89k5eutf85CrTCiStuYMusXMlMyY2uSL9/3xcDjuqZ0Y9dUi
zyJYzj4aFBK4AGc838M3JWjp2YKmeYUQ+ZT1ueX8KAtaPEJR8IV6kETGViqbCyVk
iWedpwNBV/uvEnBLezt99Q5cG0AHDNzLXZS4SruSIUOxqm87vLNfYtDtNPQsDnFX
Rs3i2qVlnnjMPtDX8UzIUl+ulhyeTbu3GkOQ+WJcfp7ekOBdZutSW2JkPcSpNHx8
zWND03oqyrsKeXbIfJJMe4gHVTxnRfx0gCULnCZaHiOxIABH6yp3T5q4Iwqmy7Zk
zWHA64nCdeF3dsS1bEC14FcnJnKvCcXKlByLZBH8JOFn0MNtIAK9H5JyWasoUptp
I1d6WqLnhYhUuFg2jby10dJGLJ5NM66utXzQbcVabFeAiehNoBP9P+IASSPwhKoX
KrjmGrKxmczN9pA2IKXQJrsifNvSPSdRiItnCwgHEgf+MFESzYqM+UVuU6I+UI39
YIgsdetV2awIzKWJzv6FZxcTRw6bmU+S6ZO2Z/2UvCuYyMFqFyOdQHuG+LLGkWSh
1/8EsG1nAW+XeoAe8fi6FODr82VPE4Sxh5kRcIXb1KpED0TvYsXHtgDxK9AwYZzb
wJYQvzXSfgOy3T+BrpE2zR+MZLfy/V2P0y7ZcdJ7joTnI78OFHKofns35XnyOBVn
UX3CoLpTnaIb9kznKhqntN4KEHuOUb9pWX925mrj6Wl7ql+3YQ9f/qJZgjhIz70B
ZtA9MyunyQK9oAg49LVnkVbj5lqq3sGlYyh8R+i9LNVgMo9rLj7G8L843exCJp3P
rNQ8YUxTQJA/2n1+FdeN1+lrxDSVYnsz5LlgynZgSgTsgDFa7Yxq1rn277LurNzt
Y7Jh03vyu0qIHj4+oyY0yztkmkMeoasQthRQGkfL0aMTV08FmxYVhAxtttZbfPwB
AKSXPfaMNde5Tpcis7bH6uBo2VbVWu9aou7Stg8Pr6UnswusGGZCkQCvRNT1sK4W
0+UCb5gDrHtCxLT7oR6RXaUQt/84eyKgpbMZ55yHq/tUA3CTzbxUtR6U8e78Pvgo
ODOGYu/yZZXlWa2iIdpXcXxgxkm8CFAInCXIRo3w3QVIeVehpRPPTKxTcgwkHnCI
e5GRdtnkiuBbQEaFfgZTQBOSlgAYtS3mQUtvv3l9c8ypfOfK5T7ocKCnJCzIh/oI
orehfaMZqJ2rU75iKQLIzjRNsKWdzeB3HCbWxeGfvc9op19texAJthy93fEmddAy
CXbduMnMyJkkP8gSi0cSy6HFs+onD9irtPO7DfxdcxL9cIke0H2+186Iv1mkonhZ
yf65ggOUq/YC1SK495uymoT8Z2hococer9XtBXl7dRzS17yNcOb3oETET5DoGjYh
aIrag6zTe8oFDgpUsKyLx5f6+8CQ7OSSKrOd1P/yWNDUy9NwHYreQZ4qRelSgAtJ
8oUhfLlxNu9x++nEBq35DQEGhgf6aEDu8XKcNlPE3RG1W06LHmy8GrMsnh4zOGCP
nnIRmqBeybrxtqH3h+7T5yWYqrxea21uZokjmJNk99U1ja+Y1toR2VdjxdnF1ZW3
VrVXNwujB/6psmY6fyFyrUoLNLO2D1tJw8gtV1lwdbvLK09O6sA7agIHFdppMfBy
RDuLAr6/OBTRsrmqMnqBFGTfIi1EuYvnnV0wjKbCQNs3ZMg2OE7Pxp991FGvALj6
jlVJxoX1657xoNUyHS4hd+eTONX/7GXGA2Cd0yeHL82VuTOc6n95zJJGc5B4SxxC
uA6VS6lQ8+FCG6I77XK+P8uf+J1j6WDF1At52Cpts5Pi/y9DvhbwNriGm9+/s2AT
njdPa/jcEMf2y5BlmbJ5BNRStNcDGvo7QSk6QH4Cp6HN1kTbujuGiyrrl15ifdCB
0jSShdke6C+hFy7QUbgCqECTeP7Wv+LeKzyDBRgvEy/CWDFr/11sXmJlBs537EQZ
IxQimKaPii9W5VfgnsZCKxJSTtT4fnLuSooWlPRIysewrpndvIB0dn8NdzQJNeLE
1UBqK8/ytiBG6F5j/R628OxFc6B6V86aNZPp8dC7y9oMBfIrk+p7sEsfwYo3Mwyw
tlp2vlc00jksCHye4PBDo5EwAMsdImOSPYv9z+jxZyKPcBK32RpgdXblUdwR6FAa
e2G99fkXu4bFtVl36NePkYWsAkDDrMAOlcMNcB91Nb2WU1yjMGfl8P/ywvDQkTvX
bH5hIcKA+hcegfCG1U7f624adsxndLzaX/G/YZFi7CDKpBBDKgWHnvSXw1kUdIQJ
0iePJVKuWf2ifAOoPdLUvakXeb/Kz6SzrNUbljc8Cui64ahs34gqKe4PDYnMOWCO
CtGubjP0POVpXmaBVnyZccGqvoQtZoD9go/1f+PfNwPYOxS99PFIjdNNvXK9eG5j
ZSQFFkMWkloi0HHMSr1PTq6sz8IFmZbxXJsmJz3VwLFQhCFIT93juOX33IN+ILig
Huv9UwPmybly+Ev0Kh/gHTyeOsxSIubdqWAEHSyp4XelNsZcEiBFNLq+3aylEL8X
VHnpQtg/yn+fc+pKym1a68v2TyBWdiBLAY5SEYPw15v5oiI//8qkEBwcDJHs2kH4
WGkul1M3VTWu7yGZH55iAJy7xTSAfBEzvF0Z9WyOHOVZeLMx1D7CqnaSq0JDdur/
ozphEnsnUIN8VBpuDkXuhWu91rTilKLKn525+RaWvjtn0O55FjpVF2N1BQxlTH2Z
z8KxyDhZxnR360yEx3IFr2b3n3IUaPSkVbOnT8/LcdSXRQK+KsiSn+pgCOb4GlkW
HeyZ7uTTLiUHwpAfY0STtYKPigucdqJCRySV8kZcmMx+tCHz75kkuc1RSas1uo1J
oePhL255HY/MJFak6wnADg2696zx5FdE7N1mvYNYyIJSc9FZYs6wfCTfzLGsfi7U
oD69YrzOzmnJCvJvPBEDnjcPQ6aVlyk51cNxiW21BodPVU/2iW8pfWGuLUEDjWVW
W9iXRVZAuyzhd74bdbQZx8lxxu/USjy0RXuxsjMlPT5PjlEdsMhpSVgVZYJ5alC1
ve8DFwii0WqM9quqf4sNnKixWTK8lvMzC/3hexMFWlqEk4kFfES2Ir5bRmywi60V
8qeMYH2io3//BOr4UF2QhKN+vv+QNghdMOZEI1pwImvjwquCHdJpxMHvPVxynVg1
fRgaQmXtzUQTtSFRePWh1shb4KHGHXY9URb+vwGK662dHaV2CO30gWEGFTUVKNkK
DlnirxNcOgE2uHHMthIsL4D5Z2XHHu87gEe7m6qRK879wDQAc1TV27kQ+v2yQ+LF
igOOwLtLR35jGlim6z164z0AazWvds9s0K4BvZ/Sd2bonT2yk9nJOT9UMDD6uQUd
K3sC1XFx2WTaByQb9+HOeyTFWJWGeSKuF5qCH6CoZK58GHGgXHft2RZjjcCoVSF6
Bzsm8rV+actujWFZ2ORwoKCQ+80AcPNAAfP41HxRqQaqR3wKv1CthQL6sTUl35SS
WY0l0BDD3i1655fPU1kzye/4YzYe4bItug9oY4ZvIyKvH1AlgsHEO8472pl3+vyb
cIW3qQG961zs2+Jv5nd8XMl96YALXKansMN4Dpt9OBQffB9F8OHOEtMe8hdN7sa1
CuDgOZZkaxcruAmgv8nfRgMioAIm0KkYQ1tbPUYBCgWL7SRU57L2Qv2qe50hgMNZ
5z//T3vlLt2nsbWf7PGE+MnNbxmbMiyYy/gI61rnHSDrR/UlpCdFYD/HokwITp12
5gQK7gtywTI917KCfE6KL9RT5gcJ4N3I2/cdDPRE8tHGxRe7b8RtFhsNOhqHu5Os
kmERpFFm3989UPODnsfLm8M3wK6LMliDYQ46BsCHisyk6sj1kk3VdYsDsUUu8N6G
O7WGmTaTeKFZB4RIiVsaoj+hwn3aee6NtxltjNiQTCh2mz17vGqgoAYS2gnoV1xk
UuCxyjqe13DY1F9f/F+9lqkIrco+hHIIJbo5R2ION61W8P4GzdITLv8DO0byu6Wi
2GuZic/oFctjvj9XvOB3mck3s7gLJ0ns5n4A48yFBrxuu1pXnjyykj1XdR9yT1Z5
P33LmYLTJE/X7IB6fjBy2m2RVNp5OKHAUcHc9a/tObT81WQ0cGHQlpgCI7lKfifG
o1zmCgINCvltrVFGFd4UomYnaxsrf7KU1er6jlbYaAIuHc+hVymxzkHABAhUTbe/
RS8C4yuMgRb3ywe+HNROiUlcVW4x0iHOKwiwvuRwqJm71cUxvjWdIsnE/NxA+k1b
UX9g1QI6HDzNHT33CrbywLV7Z38wkpkbN6RahqTmkBqNMJPPsYkgOWBgYnxg5K+E
1/HFzuN6ZZA3eiukTxPl9bv24Hr6I8NyG7sHDiVJP4n3SEo9ho1KL3zu6nAwZ1Lb
ogz1tuopqL4QdazbWXgPNBqxnVFSkaZQXChuRVqwODLjzPOD4kH/0A2/KT3oARlR
RdOSfp0F1lGcLKqDfc/6VoqvRxenQRJV5ChFgoPwuCAzudhDo4Tm3x7Zws4+kQV7
VHtOaXfCxTtQyPTqqbqDp/BUQcLvw1SbAs9RNqezZYGyaTHi46u+f5lh1Hzy5Tqr
4Es7eAzRFUIM8/dDJdbl/rbzc6m37Q84d/WwJg+MZFR51f1xBRqaCDXkdntAX6Tw
/JNJsTRM9qZS9n5VuSGvMJUnQHUJEijvWpkAx6/h4rNa/c9/TCnzPW8jFG5BWD8+
eBoiPbzBpuqpeI+3GxsjOUPksx7QNUZemWFOtIjFZgEL+J4Edtpez/8ENnZOBnEs
Ys2mX6vvUAqg0F4iWqWnKObAeqMDnPWc5hIEZdAPQxD21C5wHtrM5xTUyej+bk2S
E+ugWsRZnZORDDBcvlKPTAT6G6AZ3xm9B16ot8YZZ9kBXArgrHbQpP4h7o2JPDzz
YRoVjNyNU2Qa7a4/X3IQGX2q/gIVfYQQVJ6t7yK4yKe27Rdo1Ssf7GyU2qxUQhhS
TTkJEPFk0W/ZyyVOiPVTPm+bZ0+2ysx5ksVl9CpB5d8t6XmEoTihXnFb18M9PYP1
IM23KVqKKSeYIk1Iek0eGkBOFcDTr4aV77lk65xBcSlFINCm4wlZKBXeSvG0jyXz
S1M8i6DxfMvqQdJP/HPyb6ZJm6n4HWfwZLz9zSvUaV4RqaK1F1wRi9i/mqLa3GRZ
piDbrQdZZLjWxcdtg3UTeKHBYwIvqLeOXxveJiYxDBdtU9f5oaq8WJ4IiV5DyLuh
vqrnY+TgY3BvicB0VjspQUhSeNn6Ta3nJd2KFoYS9natzSaFVzyW9Mg0UEWPmD1G
wnxHKGHpkuKRictp01Oo4Lh5JAyeNVrtZgjB4HbB0IbEmhErunNM6rGYOlvDdFln
whpHg+eOgt05bIahebvsIs0imh25qXFf6ZoOX+zPxiYSw1CiZWtmDEQfl3RqfQ0h
rk6pI90JtxkAS3TRzXeNN/qbqS+rikB9NzqP/p9VtwCs4/0Gg4/+oGBDFgiUQ5Qy
sTdQ30ckmai5ctlD2hmTOSSOZxnC6Gdqk9mNcpjgZqaNWeQlt8CB7CXoOehQBB8X
2d/Wh3krxoxlQrRaBZLFcwLYYTuq59L8XdYYXLXC6BkT2XrJlaJ3FfsDbSZe7Ea3
8r2sHKL5hxeA28di5gOvgmZQwspQ5Ve/rASWujX4L3MRK0nkemg2v3uoozFKLSIf
TVJiltgGrWoF+jJd1GNmW4ElrMFWft5RgCqmDu+9CQnog6JOq9hZK7Fa7a18Jcfy
lBSMWy/OEnZO0HKSTfJ1wUO4F1GGEPCXOrWqWnc+kAFPqg1yIzwC0nsP9DzcYarJ
K8QuGIhZa3NioPuo7JwVCuR0XM/ed8g5RES2R/9EILAPbX+vLSAnJM6b0QoT7iU8
Ux8FPhiTCxpWLrG/3DvHt3XBZdGbt4aQUowSsMcjL4yQfbfQ0x0r53Bj8DOww0jv
iPOQdN4gz6uh1zyqH4N+AnXAs9aQMCj1tqgqf8j/GEZJ5L7l7904DhOG1DaNq9D7
Bm6blYmnLkFsmpLwzK8jORIgoWUF10Qd0xG+42a3jHZ5pCq+Ub4R3XLhPndcsKNU
d3LCQRxu2jN31LRPLzRQRlxUBA6kVO5oinZ2MZyGkINwOPV7CGN4bbNljbu+SGvF
hLkQ6VjWrXfz0VT/PhvUG7nXGFARl9ykTwPMsxF2JkpJ30f8gzz3HKln1jAu6Ggr
MsLRG+qfuZmldPCFBk7ocDZHkTXiqXugeSL8cqsQ4Nb1kBXe8+SYhtcbUOaInRxr
CNcx0IO7W/tVoVtpWeXaV39U0FdC8momcIdbMN6jNwHQlFkEyoPtTSHu6bkwd4uw
dPysbsWxzU9Va7mLanls7ENVgLB+Bp0ZX2a8hiahDw/ozLDXtWd/sgSmHLxGJmv5
RDgvvqQiyNJkBWCtdkcrylG/evy1OGsD/mxcEnXkpmoL7MtyPjwwdQpaGCGezzGe
xciYi4yrYEdDw/rRR8NrpdcjRpD7ohnPu0oa6Wq3GsmGmXFRYeaDDPZdpGs0a/KN
JFVQgMrzOxsBJIqeLCuUi9voi6znzyRPziVYlZx+3Xi/rK37/UnUh6BrOEwWy6P0
3v6GJ/MkaJagKfu6uuzuZ5WCTD2zFsH4/Ku5Su5fs1l8hdR+DnaxmLrEsa6qIckb
Idkm6AxJQun9I0tVVw4K3USHrfBdy3drTnpp4jO+tZJvU1b4oNJtQoJWGZ01On+x
sYE0lJm6WveGcUdUBKbdAmio8zpiM5v+Njgf/A+Zmc+A1rWxlpdJuiWBncZmjwyi
7LEDtIjQSanZCUW4oquDbRPqZ5tQ0cgMkdE3MyRiP6ZHDc0xrbotr6ZF/9ucTJCE
VvuXlxSes3zl+RanEGP7jKrNoNueAkGYTXYqZNWXGrMHmyqUbg/o5XkCeVGnXy6M
Kxde1Mm2llHUzFwwHY8zfzFer/KXREdgrBiqabjutos+eEbqf7sUY+31IiLvrG+E
U9ZiJ7mQLA6YB9Av5KxDoU8yBlD3MNhF7ZKXuPlpSpzWSOjJXYWHTYnlkOSGG8uK
0eU0gXlR98aaF5OHvDvFitbge55zmoDfcyQxQKGkQrdKjbFSo4eCrh0tY9gBjWYE
5yjSj++UFl5IUDoXxvvdXC/yf9A4+U1fm/RS8Pxng32csFI6cYEZhQQWQBsk1oB3
wWorLVQCq4r6pwr9woGRqwc5TAnssZxrRZJ5lr9rpbUEqaPEtCBUXGW04sNoI5j7
VkpE/Kii7dH6710gbLwDjmwbvYoADedBYp/d0+Ok4rF+EP0Bgi2Ic8bg49Woyu6m
rJZGyb7LISUT6kHIdNVoHSZbVFvO9eOJ95M/9DraiLoZOavgNzr1kmmxgfQBS3/N
RYweqKYRzBdF0rcga5kxTht1hjySKUmROpSTT3Zqz+2RqoVVMA5btsfrUXRac8Zq
Bpr2MGNHakd8BMcwRusls08VTdrBLpVNr5DNYSR6hxvNBvtv+oC7ljvnPRK24yGJ
PJ71p1pF8RdzqBEMPjo/gPHICmcMH3ADRVr0kWgHdPwddkBCHqKAkh33KeFurrIj
zqgAxqrqitM0kMoHKr6sI8grb+u+DdxUxFY2n1uKQiqD8vue4QIkUHXEzlmCpc4A
bDq7MvzBBw5H54nM9mRF1mys1GOJO9E/CXedEwmrKORyCydzW3Km6Z1Bf+mVIl1S
YbpWA2HZaQe4/Ye33MvNRIVD/ITs4XDAoY6/wMsmKcGtghPBrYaklTrf93IBSKEQ
/EC53ntUCZGHaErxrD4uyWzWkAGq+X2bgG0pyM4DXv3p/L/YQdeAlemKv/kcPG3G
5ULEfKSUQ69xblKE27qjofAfX27erkuohvENUqtQvblHpaYbxsj452Vntg377D9g
WHMQO02bl0uKN1ZODycJl/JzgeSYHF6EDv00Hhc5rkXSKMQ0OriMwVbjtrhwhHCv
U3eJmQJ068PvMRiLHXjlhEySZqBtvtyW0eZ2XJjAJpZuWYYo83uXCn+sB3fMiNXv
47LvSaTgIqgS/5/siVNUmFLpicJaUrzzyFJSkV5+WAjL6Y0TBckY8MlOfxBq8hCW
EEl2SjACpUAf065vxUto5OOjxpSUi5TMEuCxVYMyGowV7MoamguPb6ha3+XqtvrS
HiRlqZG+cJ2KGFF0YiAU5piJQ/3w7WwQL5CAiaUXAM66VtbWpnV8lTwxh7x+r1U+
SXkpy7ZsHzf8qHfEyLj8CSQ8hoO95v9xQ7Jmsk18zGmETiTKUyqfhMcprOZYhnoE
x7ZAPgW4c7PiAFhlxYZA5tenqc451eiBkJ1BkbSgvrxxuZk+zm26HjVKEWlRLZR1
c7wNeW4/WgcSN5bw3itQXb7T+7AZDypLLLqIvg1zR3Dq9p3eMouosaCbI+Lkk1vr
aGYx659EOmImpyWK/d0/QIq9naFVXzOKZXPQ++7sF7qEKlPKmIMPrzcmwh0j0P5C
eJ9V2RtFvPGhRAV2E/Ck6ldpxuAtT4e2pVGgjRvEGPfyEHv3UXnQmXhwh9EmFYTG
20otIgUhtWavuXEEg8Zyx/iJU+hSodICSUdcnMvujFLIpOrdVqsZ5ofRSpNhpNBi
ZUVxVmlyGj/evEeuqf5yp53L7ocBvG5UOtY081MrIdCm/M0z4SdHi89JT0Ndfv6X
kd+CjjaK6sUAMoEcTXXTfrFDA25NHJOF4egToL79nWc3i3PsXQEaRwZoAb67ihd4
sAUTdxwow8TTFfADepf8gMy7KhwD7rRG4leHdKWlFUhrrzrXY7YfdCYPz3OTFLkx
4EqSKAvs61VnpkygF7vF+oxSfhRkojhNXAdpHIuocGAoD6IexhiAb6p0kTDViiYp
wGlesU56d0LvATSyMKFbLm/PbqkSIF+mrOaDO1vLQHLsKpe5Xbco2I/JJuMk+NW/
DJgHfeQahpS5tdM8fMbigEJzVdP9BY6uQdLOOTaTduTrvSETvKu1DkMD36xJRb5f
YDlinqSWhlaoo7hwkP7GJiW3nNs4PUYIjR6ACFZ43tyFWca4GFLwJBYELL2Jlmq1
drQlKGBYbJRprfZS2914CnjORCZ9sMJFznQC3cbjby1O+DYghuDMuhimOGZdz4Eu
HqnTfisBONfqTbGgS3YuHepjZ2Doxrh6TdCC4CKUEqWsepJo0ZO98ZKR5h+xOVZk
R84t49qvy2NaLhJtARkK5CqBQ0bFl+WjjpPtnhrV5FRFyVmfzEzeljh8Ec6Ibo77
uZgl7TasA5fgcysUUi373hrlQG1H3YmheOYXMXyNXHsFkEgGVFOPliUdJ1tgnDEL
MOCi7qxk9cYYWyN7pQCWVskwdbJN3YNOmkbPZXSvgaQy4eiMclXAAw3VgrBCzQ/L
yez2JfSk3U7Y0dyRUIrCqg948AtU4hhbtk3i0CGIVABOcivqa4MM4pNAuOtomasY
739AD5EwThBuJ8s1iYzi26iYNUqJji2e3QFl9TX8KFpK9v0BHbU/5gM3jOsfNiPR
F8LJcKWdEPJpMOcrwl2+DCyNC06Q/W+uxP4ows52NcZX9tPjF0j6DxtIMq1oNIwT
qxCbbGI+CjjaU+dVomk5qZnPHMcq133DGOCF+EKlWy9dRunKcpZOQr/TFNTMqhY2
2pJaW4abMn9x3pSfSVS1GG/lTD/rz+hLgDIeFogj419Ah9lSgEEhW4InmLusb19c
l0EXE07HfiV/3g2RPKBjrNry6aiVnye529lGjCqUsns0rHhymmdmVmB9g+rYot36
0altILO+dMn+DraUarHk0QVxZRMXM+BzjepZQmV3DkDTCiHelLfzhd+QA9d2ocJD
PBseUuAEHFtgD8KQFSj0cgii43BHXjbS5r3P5yfn+Zpyf+LQxsTB80B9XO/Jgo0Y
M+epMfYHrEBxf83WvV1dd6qVn9qivEmBpLlXIzOpbpjYf9E2EFBLEt/2WUV2WupO
QJ5P6xcZcAKS7E80ZHgmKxFUaV6/74BNmxhKi1ooFiJOqJtZPQiH4JD0eW4MFS1I
HtynMFqLKvWzUt+Z7qSjZTAEcOmy8TmkbyZLqqv7vuEtXl9VVQ+TSdItwlAUCcU5
e3ZREJ3wSqIql16IDLbYkNhB57Jqe+CZrzw7UD6jCNSfm7jgFUxnZWEC4xUs7tbG
Q7itZ8xFNEaG2eyrwafmXoPLNgxPbqI23ZYiLFvxLBlsZvRIvGjsOm+FJx4Y4GVl
V1dhapZk32ueUz9jeeh0m1Zdrw5DGs0kByFokVK6Zj7eyuaG4WveHTYUqZaSBx/r
aKZOniME3ZKYn/yCGetXgXnxCXDVrQ0Y+QUTBmZ/e4SLguEWmQuyNLoOP35GfW/m
eRSqjS4qynJTEbsgCYWYptP7OtBAiPcXIXxU2rGUfhAIYe2gYmJOwaVOVW+Yau1K
3y7phFLfeww4ACCNvnmB0tlhUhTuVAF304Qs06+DKpCYtqIh3K9qQnRCJAHrt6FD
abIHM78eISQyXNiiKakaQtWyeFD7V/7/rsuu7fB0cEjg8g6Z6NRloC3YMpB1tCHq
m41esSY0f4uXXfLI04WOUukb5unxa3ba8yaC1Z80yRoZOBhnif/tV1P5yDuu2lhS
sOjLudZt1kYUlKiAdwNPU70NYv2iZZcOgooLv/tFerLgapmT+zcp7Plovqftornn
NFQ43sRA5SMwksoDnJRDVq1VDteN57rtagQ6mcymB/6/1yllLwaDU8RwBy+gB1bt
fLBh3B26kAkVwtYVnujGffCcl8AGUndl8kckexZO77tj6qguG1qJZo9+5Him5VJo
3/dwteuifPByio9pp0ZvbTchAAh8xkfwLOv07jjk1mkPtdMVgF2sFNfav7eW4fIG
xIkWW6qHcWsXs1zU/CeGJk5r7B2UtV8G+XeT6f03H2mnacatfrF88m9AbNfGY8di
/PWLBFocEshS+UCLOyvIBe3Uwcgd3OD+PTOH47wbKZY3i0PDZYIjI//wL/mGdmC6
LCG9a7X/RyMIyhRKLS1b1FRV5gwgxZx21zHiYT9ulyEEF5XzVOG8F5i3H1j3kuUP
9kJFDYheaT77gUoTr+wOI9Mna6RuKQez0KGorIFKlTO2xUmyrHk7frlUz+0iKXds
rdrttNaI+/d4ZDWdHVh00JhSFHtLcZW53f3SIC7rAs1AV/92WD+6JVOBXd72451x
DSz3M4PzFNxfyWCLSpEaHiL7WKrlzazRkyEP6ahFsfGJJNq86E7xom0BTlVi1uzN
LoDOMS1SuSJGsyd/BeoJh361uscO1RXG1yfkKgJ9hpinUGsYZPbTnCPfUxlyeZTF
q6DwL4RTjo5UlkKmfeHKXWMBqnAXOFKHrRJz7S+0DLSkGIk+mN6ALo87AVvYQ9Gn
N3yvSRFXrqGOv2KmD4YfzAbY93Oip0g6MZDs/95GdR8KQjufnS5njFYSJ+GTboc4
Qc5lt9Pp6IhBgBAQBi4atv9yQ3apzU1LR+PZs8v04cfB0z7xRhKdj3LFANRiasOP
U4Oo01AmX9mdyOyjArPobsbplIAwtN762wm4svgLt0mNyyEkqyDl5+3UCHlxMmRe
GNItwK+qTf8YgYHoGDwlCO+WKA5dIQizHVpiSD262B6LSKgaejEJXMWYNNUBUOTm
ASzZnX4TIo2cMGWNFN8IEKeT8B5uq40150WU9vvRyj7U1QPorAc9oNNVP6seXrnM
Th93Eab9WxGka0F63OkPlofp8kzCGCXeHHhlh+R/5SEDEvccmbH1MCV+SnIvR5dU
jTitAx7Qm3MEvu6Jwyg5N2SB+yUrlYej5iE2+jKX62wIT1fdhqYkTzAFADC8PUpE
5dXuXNL5Sj+0sx8Zf+DeOvI1bl37Zuc4s0M2N9Cfzzj4kipThviE5ZRaBnrPRpal
rK7DrLjL/c9MsQqfp1YwtfcfU0Tw1LoK/DuK059NlFFqVkM6/RjdtwYPDq0/qoTH
pHBRNu9rRoUxDeQEhNbQ0mPch24VedoAb8t11lJyJv1maFrsvGnw+kZqLSU1V4Sv
kQk2gAfCxGh1PqffDIAJlMvd90dTG5yFg6ZODVB/LPVIVRpSIZha9NWg6426Eass
WoJ+oIVOaPJF00kkieEn+2Dr/yXGd94z8AfQ1+L557A6PIUyt2jVTxIyr800Iz0L
SZQhjYjqEplBqffotrjKHPIP8uCuMDe4b7VW/J65ZvWql43Co3k6epob9hlOc/iJ
WKlvHiPnuXmmkh/tb94Dg7oo9XEHvpQQc7OPFPVeBhXRHNQNrlVgrHSPI3uvOWjN
3a5NHuvdfBm36QrChavjMZE2Y6176RR+2MWmc5+0vFfqBbdG4EVIsxlsT6/wZbUB
EZH1iXIE3Ko74uVR3t2Z+IG150F8tu2AtH0HD4T3U/3OYfigMzDVQfkhkRzNOxeK
x4zycZoXjDEfJpXNa7IHch0aq8VG7GXASJndhnbeDrVdrdUXO+6fzaprNufnsL6t
iRUXaowsPgop7VSOy220Y2LNpUJ9cVFi/a2DQh1j30axUgQj1ziWlUbfu4pvVd1Z
vPsndEvDCIkrKQzFF+nDtfANydblkmYMoOhwOoRk+w4RYHwWx0Sigfyuw2EBo2P2
qjy81v2KLPdlyh7H7R6WXeOi1tAWyCrtdeCbMdEOFMxibjhFNlVa+XzzZy/86Ltg
ElSk5oOtn7A03DwLKZ7Rpen5eo/t1cbXpVJxQnuwb/ibnxYYgBMTj+oY7Xj+VQv+
b2x0DsJ1rMV95VmPNmm22oJZC/Ik7dlOqIJ0Hb096On5DBB7OwLrcBNw2gvymWeg
o0pYTwwqrU5xzFe9dAJFk28HibTlM4PdjOeOTJeXVgHolwgAgyyN79nDA+Mda4rM
GgK/iNGKI5bVQaSifHtwYdSv6lK6FoT5tQmyx/4JVxLQLw5r+oVx0KJHGjHNAV8u
n1ZmPCZDdOg+ATJocWZ4NVQYdwRYHLmdONdPI3xZ5IpBbjQnT026uWDrzoW6GUb7
yR8QshTqqrD+pY9gxmJpx0I1Ww1Yqn3QE4Cy43MxkmWfjPmuw64Pc7POQD994C0h
mwC2PMoj5+hqu9Tz97lZ7m6Idr503C38SkVJeKSkz9SLQiGxNLexhG+hFB/ma2fW
jSEpMByRTDTK/tqqMEvKXIr0c0dRGhSjYj2Aumf/aS7LeVDmksvR0pAsDHBbFTOj
F+8G9sPQyz91zziLOEjmrILxFcBftCXSBz53CBB26NaQbHKy9luTDimx0exQvl7/
zKmkT0MFMjVzu0+bq2aPG6gcbce78t1SCvaEKVPPW83NInPjjb04/whUsiKBGJIT
ro4HsukWqMabAvHy3gU2c2WyMQvi4rjG5SwSqxGl/U7JC4wBYZ49a7UQtCmjIi17
Ey428Kk3tH/9WPoQBmCvQLgVlUyWwT/rf+wFS8TgYzbXVyVkI/FfMTGfltGX57FL
4jjgYSANpcPtrLMuxxwaEI8smEnWe+PaFXwkK/1ZxgDuZhh1AdfUvM3c8t0BdMpk
oAASOe4GWmme0S4gWkR5DArlSPFDzf3r5Djqt6oAup++7Py/XI5s6yAECd2mPuyb
ce9KDHqNImlQvZqRB0pNGTnSR47gBB7Jqa2VTHH7kwoSQMuSJEqlPxaB4pJg+JjL
Z9LaJPf1KJPTMpRDfQLJ1IQ0UfwDCoz+JUm0Lmp6KPqFGryQ0JAY9J1+VSmehxf7
53bBKEHbGF5fULWJ6g5bwgqNy9/fLDt4AEY1CQK8z+Q/wtcRcLeCzDeQakXfv6Z7
/sH/6gVK0rh4Hrhqm08ATTkq3lQNgkCHAlsEiF5kCQSLFDbL00zhZ7Gg7sO9SEIf
pI/CntKyhq8tyyU9XIKZBUItOFYFIjHypLOjWfZoI8qpOY1WKa5VEG5i7dsCFSBs
h4/fIWPrA3IUYDfdQDuTTxUgEYkTU65YuhROS5EzjrMqlzzv710u2qKfE1q7tHDe
xSks7VHsJXyJzBiaI8MeiFWRa6FYANRQv6fU8qHaIfV3SBH7M9yX3qEBGt5/dFYq
vxd435l6KCcIIgFOQFWxKv0lNLVWiDsMB6wLfCh2BCGhTlMBa/yFkFTrse5wTKkZ
bYZlDnXlHf/e/c99c3+g+6QO/II9SxZkQB05wM7t+omGGrPPCFfXQqCkOt1J686G
N8wVjbBPqTKTRX6fFh5pFrNTKTBQDxotkkTeK3IZQFBMskNjg00BrrdNYuO8mcZy
0ezb6V/FgP3iICt2G3Z4c0PcfueuRnvI+3RPyE5SwNWhwZtmQPjq1ZluWn7qE+zB
uabUZ6lSy+O62A3ohzHJc1dTOBls7czABkI6XN+YKoTev8oOZsQ0Ps9yCRDVorRr
zI5UZYLKFgZR6CKs9oczKS52lsDfFrZIgqi8puUit04tPDRtIReZTIqFLDd4Sj76
BvDoXt1v5V7YmX8qG5NQYDMOp3A0UEX0j6DsdwCpvBr6IXFlvaX/d/0hy/KFZsUx
07tuLEVGQ2rzQwCr7cJUreQqYr1pV1YzfuE7KVgUDdwxA7owk6/FKNkqaZRr9O4L
TW587lthpPc2l2b2UBgtbQeCEflAD8USt6ymNccV6T1fEU1tQR4dNSJmt4O/Av+4
0xnEfCgxLTAoH+a7ICWFYaODTLToTAjWpIbzhQWaF4H7kbKU5wFzstZJ/gUqcPjY
uzP08jbsoL/eTRK+S856ulT43PAH4+FI/FRiEF5zFNE11X4zMZxLAVm4+9FPKUU5
wY5RU8/UQJ2cfDmQZA6LlYZvbLGui35kTrZ5jH2Ukonf+nX6ruefMPB7Z6a/vJ/x
iDY5gUKKiC9hl2goXJ1vAUdWI4/p0Hm3Y6Z1sm/NNs402FnQ1h+3R6StOJzUY6Bm
PNo1nZ1hJ5GTWMfo9Zzj3/eAgv3fdbT77ND/jsRM0yIRBly+HdF4pl5GIRHZNhVs
QL3YD5t138pmAK9R+lOkG7bPiqc0aED3//Dh6D/y2CrUe66NTaN0zSGB/zGi5Ngs
sVjnkp9wARsvUpaTgItlDRobz63dVUmM6/Kg+4MkGrE2T03JeXETSHVxOjHAiGvp
wjFitmNu2/8EVZO0MZ/s/5rN1Csp4O+vYjRwo00H1U8z1v+D4/GAk/GV5TB6pYC8
6EbH2ePNfpQGLFB/kJSz0UT/krTpGt52R0HV2PJdoDuf2+ScMb48oI57oWuJxXu3
JN+Xh8BKk8iYmI87V+vteRAgA+XWhJvc8qWG6RXkX7nHcf22gM2rft211G9SMp7Y
ttq5jZFCO/kXIs/9StpNYbl8qQmGOZ9M2+rRk6xnxOsgyVKVaiJUn+d5M5blXSWK
73L+0lf2CtWMQ/hFuZwcCwFMsMUKFeq4bV3LPGolqQMj/FymNt4sbjGV7heep9Zc
hzgAwldZHLfIiYjA2gA3efQu3xWUVr0E8b9LS1vn/XVhCSUIKpjgsQPhDIkqA8bV
THI0wImGM7QAUx7LzLZDHcOOIykVjYxixBowcaUz1QDhJB+WGYHmoeSx3yKaMtcV
6MT6kK/RtMfA5HTrSEgYslRFmrpvqGctsy+n5L3IG7194kBbnOxqdiMWMcvX+LzA
bsDyarhRTAw3n5btmjWM7qXIUi6TQx9w2iBycEjV0kJf8Ib3DJP1BL18L5WxGa3D
t40jZ8Cjs3mXXItjn/k5MVCdwPTGKP0Cl0mhDmmT2IGjU8jUVlCg/sIXjYj6z+z1
iYHq4btHMWvJFgCwPEVAZXYocl88rwQT3NVVgxkF9e3turcGA5O3jHPJ/fb7KObv
hq4Sh65c/CeH5YD8+lAPpXyJYd3PC5ark7HG88qzKQZbFlby69JGpApc1hSe3Oji
Jhfn+r8fFMNunpN9cwm4gQzSQ01SBdw+zdE+72UuXmKrxE+hILsqn2FNzwpedR/W
JIrod64p00I2l7URB5imiwmsj3j12Tg9cDhqFocSi/o0ZUrBGhu2vpHeqWk/ShkX
cSFHgj4N5BSdyB/QmClKP4NLDKW+MelL/yrt5z8pixAMPxPXaQF2sZAQ/s0jBIY2
zgGaiz6OsVRlsVPfLK3LGSDu/jEm/7+/SEpim5Vg7DmYxOk1pBf+qu6dRnQTMTn6
xeK44Eouz3fnbhUX13As2mn3srYRMTElmUdY2HEPalRYhbv0RrHZjHjvjlzFskw8
VrUuP6H+eZGrBt/16Br8Sl9ZHZwwAf3onXWpxyFjm5ofsbgns7HHAFF3ONw6Y7H4
Lt07IHmuBIZFW21LDWlf0rnXgKjqSMupdVX2hO0wWD0jI1WhsDwZb4+L3P1LF2jF
Tw2wCbdHyqzPuf7jOrPiHXQDD6kfmkD9k8AXBxxsTk+3KnQmhG5aN6sKN2jqGHpP
wfhOTffGvfaTInbR0jylMGszfCG5qLsSA/ZQxR/U23zk8ZLIA59ZFFLz98Lx71bn
+RvxCiKPvryE2raXwe72dLnbaPcJhsX4lRi7+QzHig84UFxNdclswr2pq5fPlOAT
bpHatubDDxzYyWUkuA1kqq4Cq6ae02sVJsOqG1R8o8WG4u/LuR/ElKZFRQozbeku
HeZOCLfuKTQxnCUD2q9torMrAgs+z9H1kIbIVJ77b9IUxPvXc7Pj9Z2DJ8/Ig/yx
wgEfc/gwVREwnVMsJkMxLnl7RNrRPGARGIKlUk4xYaT9cvAEuyxNDar9w8L28N6Y
SzQ85McWK38lFwyIDOTHa/EPnl6ZChsdWXXzs1Te5maI7SkVCd92vcxP/nN2KQL3
pj/k80ckxCFZHHCl9Uhx/YMMqzgbVOtj6PdXWaVfAVUebRYzQHToegcs7o3LoYb5
M5hvtHtdJ0qoaM7/quOctkdrDAXKmRnkQ1iT0/xjymQ7hWytx9hRVSDs65pzmWeZ
vvrkZs+ZDkK+RudIpsD4hbiGSZQjg/dRkL3W68BC7qgjHLSSzZhpkUJh+c21Aafy
KCC5ylTnbL7mTIJl7PXdNYXolJ4zdSUdxpsPBgRIfdJM9P49D04UMKKL60ogAUH4
rkhtjAe7GaWdxP46PIyuRFKW1fzleBZKdVaGTcSsrQFQmNNZ/QVJU3xhTUbUj036
liG3TeDC3LxWyZ/7F5NtwI1xapdTmfy1ycH8dzJt/9oDFdzsCc/jaK19xLwewluH
elLxHmIqxyo7e8Mt0b683lOXghyAxV0APIE24ki4N7Rgxp7B8PGD/LaAu9Kikes/
BJLR687nA0geR4U618eO7oRY06qcplgj3C4wZTZWvdhdGR7TvCR1ldFP0ONxRnkl
nP9s6YRdBzPta5mq0+3t4hljd3r8zQpkC5GhFwvMdP9pVGxCRxqDcGFZDhQRcCbZ
P2oCQr+Jz2ANk41OR/sdI9zwaYMbGx+yRY6qpzsTE0hNqtbnag6ZaXFTTDJHecda
334ElvVd+4gXcOApZkAZdRSLUZpdeS/SgqtJtdYEaAnkZmPAV+NYPVHIfmhwfjNT
UXfYxg9Xf22wRDKbqOFojq9X3di0YXNJR7Z2R/HmFSyiB77fdU5GI8xn0rrDrcgr
BhM56lseEuVOFS/DipLTVcoHDxo2MjTnNXMNabNSOlfBMUi6B+3YNHOvzQfZACLv
Z/oPzE/c1LKkVDUFmJRbGU3DcO/j6Ny3CxQHjCtEbemOdCbq6EgJfrlhEd3ErEcO
XyKZ37i2LdP5EbnBFG23sSWsVEcp5+vp06CIgHKCaZu1pyFO6uh+XVmnAkklwbC5
6srDoGAAhGOMcqWZMQPjLlBfbfcnakRW1VWA/iFjYODC8AvE47tqAXCMoqRTyTQ9
rF9oy22zjUs/wtjKJCpH6FMdZBPtewiYuqi8WjpCI2HuTR/f26VFflj80We6i0/R
VER1EHL7Qjykan1VyGHe8HQVrfdll5eCiLtFFUZIOavjRNoTGfNVzBUG6+iHTfPH
yR2xtMoEncULXBg7tTbSlulmnC//JbjOYulFpUPF6ATWJV5Z6sD7Ot1Bk7QH7/yo
/O26r9y3MkryQltS01hf5ZwO5UE9GR1JN5ar+9AsUbtTTazs9EKUFtimE5Lu8Fxm
CkZZ41O0D6Z05/YNrX/7YkDaYm2YDaQNprnZRXCFDED9rwn1lOV9sgiYD3tAVWJd
PqcBCizuMiB4CxfdG9mdZWfqKKX5KBxKnv4rWp77nLSqUWr1VvbI4lLocS+DFZ32
tsCZc7nMrueB+Vxx9ciVKz6WbC7Kzkfi/JRx2BFOqR91Pdy5U7FZF19KTSoaBqmT
KncoAxdazjIkq/76Ej0LKvX4jtGFGyijH1M1YYpUJyH4xhOV7Ee2yrzxXt1qOiu8
YFBH+WG+RJjZ2i/GJzl4oYb6VbRnURYP0XxFn9/FCT6nr0h8Bl1nT31xdImY5t69
+bVi0u5i73nk1F7EdW+iaiRNpEPUnmRz5mn2KaAXISjrx7i436finY5L1d/XlTVa
H02J+sq6UFABxOodFQISjbALx0JuliF7dcJve4XddNIHgpNFye6o3ZgEUJxLiws6
ex5pY5IvZPw4NdcOhd8Aucs2P9bwHoG9XDrei8hjSI3dQqG+j0H5XOF9dyPHCExL
+uISg9MiRpABPl5ezhMirn6ReSCxptolQ5h5mKmzuF59sReXueSc4ADt6AMCQ8+Q
qDve8YiyqO5ww7VWkEJmtShbliXuS7sXh4RSQ1/aOHGZB/05YefQjzFa3iFyNVrL
AgO6VibrG3phIp8VUlEjwG2pIqFHVEvsNr53rk5TMdQfRb1sh5klM0VSCPPlIidC
nCpp+WA4SbYsqNLtTEX2xbRZVoL2WuG8wMuRnDrxy3ULsWPVwtkoCUB7QmaqwyrV
Nxx3bs+hqp3OvqwT0wixvctXafy337wY4uw3dmLlXWjDRjojsP8Ki2yJYO+Zyl63
8cxHaoRFs9Od2cd5t9wZJlnkrb4Ll4uW4nj1nqLbsGjQljVKR31iEKvhLrB/adel
IH3JGMnWeeriEkC/jOPA0qu/5EnCRP+drhdoj8eQUQokTkCiEqo1G13t2NsXBOim
pvnorO+/BeY3/zPRNhCd/I5duVOsL5T11keApDPcK/d+Y3na1emQgwM0/px0jmfR
G0E2Fv/2uWF+KiylQG8HUgsSKuLvOgbGoLl+MmvGB9+cH/LxhL2oks0dPo6i2LGN
sABNt6DX0n2bYjYLOUYGhSWE8yNabxPcFx7D28vjRJdV69FrbkaO1q5fRJJ6LkxY
0BHnxs6Kr2zKLFB9NoqbmEqL95PAwHPaVh6tVBegCYz+fRwVH6EQzXv7uejQO8UO
IOolemZRVRSNWFzrOgwsEdoK9v7YcehSdqsmfB2/gCRCy1M1sViJ4CWKa8LuZFm3
FCwochtcqN3cwsdvnWuIljnQHmXLjTjM8rSgQgLbh4Nh1XcTMiFf6qaOdR7G+hV0
L9RwONAZM+9JY3JtkAZUkso9LcLh16wIIeCOvBHUit8dCgbBVHZRCxJJXEo+ceNM
AJ4KKy3ANp1cLrj8O99gLIL/HOipl3aMCVmC+kybfuyUgIHvr7OR+bLcdBpdD4Qr
YdVv2nVSNqxfzgiylKRmvkXfwW2u2RP0SF8Mui6f7grgcR2pv8ZGSu+fuZVYjY68
oCJxdoJyzoWI+0B3dSj95F3iIIj/OqshcCBeIRcmuL1hc2SIqzaP0SPUslYJ6q1r
K8t/UzpOxpYstt7AurxIZPWEynisZZ67kvx7PcKg/Ij3sceaLSrE159cOWrWnIAG
ZjbSQifbziJRkjo8ryd+7UpfM3MYzGAlAsnVfJP9CF8wwrT/jSsGmRxwy7pSWhQ3
BxJEGb1oIDaius2skbC94Esp9qT750kax0q9VOkCQ8PJe3HVsPRHMdor0zuObgPr
yjU9Qj1rUY0jqL8iXyJZMWJqnx68E9lPRuSAvhXyUEswk6M6euaIsDDLPlfkOeCJ
ZlHMq1uy9aiUpZB+NDTdV6nwVkw/QBqpTw6/mMclwL5k8MhJDrXtKH3ynAhjFLFb
hIrh+6fepdnPwJrjMynWCfhXbdavIFWDGdzymaw1k2qYZk4NFYqrIRo92WGpdy7b
weI+KnPD+uB1DgjG9AIn3aSBrtLc0trcIFbmrHTDPdBRwIGbIAjp/QOhigc3/wjR
xYJLMOc0NqZ6lcDlBjo5grK0oed07oxps81/Kk+rcYRsD3t34q07uRxlhKGfGpea
s4Ct/P86oO3RhuymO5a8462qi+9fwwGBbjgtd/4I00fv3jZJFAHbi//Ka3Z3bAWh
VZkCDTcPtxV20n3GyPDr9M4fS9+DqLZR7yYGkvsh89Eu7aZUGHQ2EJewjDD2SKVA
ycg9TXj7DvPPxtEkr7Gchmb4J7PZRncodVf3mRSdbIfYSibPgKPrtrY00q+qwEYw
b89KTYkekNw0wzIqzsrSOkA8Kwa6R8uKv5gjHa6BPJ0aiNqW9c4oxxlez7g3m3EO
PfcJ8bbftChlv5XHxaK534KhKY5q3V76qevu1XMdmFxRYVQYuUsKpvrHeE0Tw6Ci
5wlTfOEb2YTQw8sQlcKHUcc+DBFr6vHcIlnMxXvoONVbqOT9WXXzYanjt3p6VgZx
y2Pi0d+l74tWnGBOSK/iHtdo4e9jc1NvFF7hmCeNXZuKfZI/03G/WXgHb9T0NtqQ
lZ69W+rwsj7vc9xPPHdJouHt0jBGj6kTTMgxlq47SUXbp2EmdFmsNyTpZkSubNpe
P64ArvhB9XAhUql1Z06sAdSX4LxlH+CEZ+wQVpkBmpIHgwNsWtjygSyL4uRSARRc
CSEDwvXE2mD6dyMLTyZnJ1xbsOSjs1Jt+zt5Qd4Zx8KpG/w6qLBkFhimE/g+GGof
0OcYEcMyCvM63BnKQmeY/n8okZpmB9v/cncN1k7SDwienD4H3YCoPvUrmrGXf9OL
1fRSslCsjrIZjZrUrUro70A/BFHjEW5er88TC/dI7fVSqbZCMQc82Tn+6MlgSrIq
kXA1+u6ThYe3PvR8fWC8T2ny3ZJeJAOW6WbKN8XTWCUOSZA4PTEz5tEyYSA3Fq8A
56aECU/bdF0n94EkoQocFlcrhXxVSvjsnCoTIW3v5/3khcsdXet63daLiKxQktHF
GVcW2ewuJRIddUU8bqmarMUy9EmkWSXrx1xD4JsRJX6i0nnn6uljETd3BSCfneVV
RPZauawLi2nrDTBfPzwGDdGqfw4RPj2z7IyEa89xOl4YJqb6ZGUHB9gtCOkK2e3O
FdkGfujfTBYwdfNJF3tCrVl2zh32s9l/7LqY0TL5gwOlAGyBc3l0YB9nEnxhxkY9
PFO7jVE4iKLLcecqrhkElO6KT6VROQKBz8MFwO0roR4clFCgMjzNr6Xs+LDx+o4M
KazeD8hNSRdlIiOu81XbfOQoiN3GFKSGV75sF2z3dZnSfY5AMOx8unNEzq/i8mXk
PU9plKpWY2GAn8xQQk5dKoK1HWW0pxG8eXDSxAsOWLDm1aYXQFJCH2G59vHJ3Swi
79rKZf2KHkv2mrOWr2282x2RKLQ87+vWd7qCwWJ/xyQZrO1993IcIXYfQMx9sGHt
ZkF+Br8nEDJLfPss7MiMd853nSQzfo1MDYHGGasrVL+G7cL8ENl2zVrV8EMG/QO2
/4Q2PIaislBD+V8k1ugWmY48ZsCfOviS+9VOeIDl6+3Z/nbc2Et3gB/ZOgkb7Amu
bztkiF+K3SqUYbDP06jYVfAAoNdYPvi9RbDLFx0ruvDi4e64Pvi+RX3uYC6BKxUT
kZewXPYnDB4W/5TZgZ3owOtzq2xVUv2pIv83QutpbPynjarPyppQnnUVQ8zaLxpT
wfKvbmLSnrGdZHtWbxP6Tr+88LvytfJDlVkmvVJvudC+MLvgCKPplfJmhiYU6ME5
V5s/nDZL6HUmgoA6kTZqf1RjPjbYCtsz9ZLWuhc2ybZ3IEvAWnSRcmExP8d0IXLR
ABpkooBeGOZ905HErAFU1xSFS7G21ZPZ/ac0Mgey0zQ/jOVxHCfsyC902CNbwm7C
Knv+BUwP/Hwe5t5Ia2a/FGx7tX9wE5romkfxAT2y9rBsivaO55uXCKsBQY2D2Wir
ILmiMSYb9pK0pZmhp8xRBJzI2WXNACA7AdBdqSjKH0Y+MjRJb4ZvFMPD39vDJb1Z
ep8lluQjHcmO/ZZBd/0SwTXtXPYPTrqA+jWuyBAzvgNZZKEGpEVZaUZmdFaK0Xnu
SchxyRJ4Wj8Ua6dCSaRNB/xHWeP3C1vh6JakFovDrxat53fmQdVu0v4kJX1M90Sg
+9DBaw1BY4XP7S9rE06Xj/9WV1mRQ/RcbG8IOBBukZdrYeCezn5LQZ7J0dqCXFWG
cEDXBRyKXpUQNgWScKiEbjo3d/wU7dWSkkwxQ38vtdbOJRQ6dp5BduwHSBZOSxUG
aEFw1DoqXoPixPI3EtKNaRMnNmrJdzo0Ffse81PEDX00qLSQTSUbDjps/AcTvuM0
JjROrRNr2NlHZtToL3edSZpiapSJKff3JqdAhBzixvdne7dMow7NFvyEDRUkQL6T
jvvMHWKPYqMuPnjTYfuE/FCmHRnMsCu8gb0siDdxVsTiD+4fBxhzsAcCZ4diAWZi
ar9OHeSXNunr5dg9g0vXuH8iADINBfZ0m8fpfwsuMTLi2qpaY0Z/rQDCs19oCM6I
yvwn/7kqhMOLmaRYE+75hESxKx0OsooAV45o/WHXRdecWn1QWrPzitwbtqKBCKw8
u+Zt2tZ4Ie34J1+bilw8SdDKhaqSzI/1E2EIMGtsVpb+VWrZOmJAY3ni0VTRC5jF
7I/NBzgx5NE88kOcMusyHVWF+Xb3fQ8hZ06waeowZiYumB/Fd3vqdAoDiTpvPKTo
P476aTQybFh8gKfTVIegIN8l0bxUvXLCQdB08qdlJTCloBJLraAYgSTHuOy5l/dS
FHUVhRO8peHKeqyRSppuzGtJihDzJyBodIX4dn7CwMO9CQ6kcBKbwTMt/+IWj7in
m/uw8F5G8B9FNEU3raWp4ag1811n2jTlS1yPlcoARFDOn8DTdlwBzbI595zuXbQp
+LVMZ0xaYUjsSBGwcgYhWVGxoliQPhJpBe8t9VYVKAoiTw1gQ0QttTarVNV56ron
aJCU7QOF1huOCdtSYIqQDoDOS0GqXFCLTd5yIWAXi4A6wYu7/tFXFzitdCmbv3k4
uwFM/bjkJ40CtEpDs+yBUjYnVNW2jwgUj/1tIY0vixKnG4Ky2uUV22QesHtAzc97
2zp1iDv67nOOK6bVmYOLGM9eXhfyTuom/kud/9qENVJgSZeckWBiG6jBRUxb3BOY
ocasCFkpSI1kcBgSRW2XyGi5C1ejSxsVaFJip0+gkIKejhJqXkhD/f/tM3r1yjdh
C7+1Lni3nxhVo8tQbwJmYV13fxkn0f4uJOd60yy0R8DEdAPuIa/Hw8ac0hbxa0Wa
9WAx4wk2qvT55lXnhnMqYfk+bbMUYNtDg4LRw1EiD2b7SGUgt1LA9mtIWKPYtikc
Tdm502N3l0cQMKuG1h7RHA+O1gmuCpcOBMjH6T6kJM6mOTzZgoCizHzn0GASF+/1
/gFD4aqCHbRkey9QtRYR1XOmGyLl2UBmj2j2zpM3TBPTUN+Fz/CVBpFZjBnF6rnh
AZ/q1jDdNflzFk3w9IdW4KHAjvdTHiNtmYDbbU+6ExyxheSFIDuOSL3V9SJlhjvK
hmJxB5aIwbG/3JqyZO+jJFDWOjT89ZaLmpNbkq5xDaJmhFghMr9oo3AfjlmmxsJs
3c6eLNPhwn4b+Ti4Mc33Dn8q0JtOogkpQ7gjebaQZk+TcY+sOW6EAvN7Ur9Mk3MP
48N6INYqmjIb3aTEiVhGWZmisIdvxejbQrbucHnlNB2PqNVsfqbiZTP+3VP4dNwC
A+YTqJmzQ3W2kbOMd42+4+v/Uq0lLKhCgaWGOojLjH5j5NrBUgkGbwM9oasLEPN1
HolG0AEpoRUgXTzaLiwx2ahhVl4nFjCMU6EBnFFwA/Ar6tlghyZGvBfr0HEL+BmO
pdYOI9ZNbEA7A1xXh8EGZ++vmOgT1IqccPGYDdUg18oZoCJLIUSUMmMjvW22n3sF
hmsQjwENLpxMbAywOSkJDEiWk0E7j0y00Um1s+6PxtGbvJPpOwdmDE71+d+Vs9Tq
e44nsB7T6Qr9zV4EOM7s/uiDHXhhnQgPEa4UgRtk6KZdV4jc7iaEtWUN/gTdn4G3
NtvHj7hTcQoxPACFr7OvxjPgXiDib7zW9R+7DEZZMhp4iY+hycMLv+jMRpeyEJu0
cYRlms6bnVpKRsH5q8mpHh/7p4/9Ep63ww2oGDbZ2J56bXmAoGTzgz7hUczcJ+z/
t4Ot3Y6Z/szk/ygisiPTXNmW3eVNyDWbzhkTe1yEdXBvhR5edhnxihiKhXDMJ+ab
P/1rBz1/P2wS+zkmn64/Kj6yFNnQX1SB1attHG3CcmZDfLOJ2Be9SKmZAC9koqtw
mm8jpTerbbh9j3ZPLghP9z8DHribIanZv62N/8nEI8EcX3qvZofU1EI8VpKRBhNm
y/gshBlYZOBFp9keBRV5YzdJ8GQ7BIYY58KGUpdeQCY9nnonvCdzOAHNrj1oXNrD
QrSz5xWjv7RIpaaRHZOBx/yRya0h31rJBe0/iarvhwZQ48kklO4S9ka5irklKeyN
Ndr6OWZfvMoC6a6csn3yO8MTpdiIJq6863FLC5cz4F66B1raulGQTX/+feb2ZK3c
hz8F5tJkcCvZa4N7zuIGR+a3Z8W9WHJk9NIKRiSEHLRaOtYgaaZgM7x9Df68JgWJ
ytmqZKMz8HRcMYpp0k6ZoHmGVF88F5xDMnNUErxP/nDcvVeLtbr8eaAB0ZEZYDV3
8XWeTkb+cNHDCPvLDGSA50T53mR8QQ+A3H6IhQU5XFV8tQcd7th/uuiQkxx3OKtt
VzQQ8QbcL82yjULuYOu83O0gPI+vix/6FypCBaOyhyi8AUJz1TjCa6py0bNKYxER
IoM57WmddJc6EQy8J4jMxoXDdzqvG4lP/HBdywWBIPORfBRwEBU7ob6LK4/WfIIu
x1bqBABdf+/yiRD440JIt0wj0T2pCL09DTDS2wrJQndgtLKuNx63Y7XXRsy0goIk
tJ94x2tleWl7nn5Hg3EsrlIaYXl9RBDVWQS/U3/SpG8MQ8J13YzIAiRb9wxWN3pR
KPzNSP1caggLA259ZY18IUAfp3KYc9qeOwIBgsIiesN9vNmo4aGpvUmk0OrpabnC
RapVEa4HgXn7VH13nrMBUmL9p3XKGLpiKJPBmMYpxUVkBP9Dq5TE9WM0w221Q8Md
X/9S17gNDgVCqcAhFCCV4TC5JmXOO0qBE8a64deJaO8+fCETxhJG9Qx0By2SAEfh
otdyISgSX64vjff9licAtJ2IBdojM9RhsdOsYQ8JpBeJUvBqU1YsilEhabapkKI8
rVDyEH/CJizCBO2SiPNVsjKfRnTE1U1u+1/RDkxcNjXns65KcfRcpspLF4ze8zS4
lWZ3DEc/oao+UjolqSsdCgH8Zy5dnbnL14VN6zspg0IZxHnebHlL/DL17TCU0AcE
AhHzarqR2+SjL2ZNbbb3iyW2JErypU+0pDH2QluBBBge6/zwa+XeQLTBh9tR6Yza
cWOznRgTaEsBToax0+hBjsvuT0JsIVch1M1zD+RKozvRLK5nHZ+fO4I0j5/CCSUN
POw5ug8gjGjv7R6NSv4NgOuEgJrwzQ7EgsJm77JI6SomGUR3VVnFKpSOMXNsNDqb
c02myy3mxET2v4Qmf6GQhV5EBteTirnVNdWqoYt/E1o8v5jozLLiZq3DAqtLwVRq
TQ3PSmWHCdlvtQnYbpcPA9GlgdGqzOFqYCxKE4kKZpW0MrbSTh8ziQk+DPweETvY
mHS2HoBZNH+wWWmCP8u5IckySlcQYqjDzD0Sz1JUV+Tt0zcazZFpP6QgqrO9o3zk
9WlHlTlkg6ystlV8WwDDP+nb+eb/TldVZ1SZ6064LJUKen3o6jIpv1e5qiWHh1x6
BOX5tgFVXQd7DAQM84YYZlfgAT+ujPMHXJx/cxPFSMn45hriv6Lqzo5HATtiJJqW
49QUYF+tzX/iQIDp+6Mg6VDUeVqfgWXeqKM+36vwO0iS2wRQKyzxB/SGf2RzIhzy
mHyNuwPwplHlXgIAjz2tYPhDEOE3KzP3u9J4vhEkYEQbG9MmeuTuBeum67Pzz6wd
ZgnL+eOICaEjh/qu6ibmgTdfjcQnoNRiPVja9FYEEWF1Xy8eBpuU+fS3m7/hohYH
oQ4Cf+ugsp7tfHWi9tMeJgs1PNsD82zViVY4THnsbEtencz8xfeXrsFbdoWiv4JV
kjI8Pw2E/o1npsoHS54GRz1eS3unLnG1dgcUs53BoZpKmAPk2no6gxZc7jL/zQNj
5kx+BcDGbH9OZpXwnTbEqGbcz+d7ne84CRjF+4bMVEPxgkFy3iKz0yINlHb7HjLu
ytmH7pTzaHw/km2G5hTqY7nJBumXGv+koY/KLSdr6HQmE5qGhvWS9k8blNcbX5Q8
Kx3FbdLTxJzQz1lmi76gpDd4F46TBI57sdjuP/XjPorbJIJiyl6pqBHJ2WJ37lNl
4DSsLFj22Qujonq/3Lp6FxtF/pL6l+Jaxc6FgvoUYVV0S/oXq9gVdoy0s1LCk/7P
1m6m/rt4xo1kqcNDO7hV1ESPXi3X8FNRvV09AgLYa6BvBtH30XaLQXv2tm4/3FAd
gL2IHUNqJ1Ukz1HEBof7ULtCMrmHjHtP/3Mv02T51+EXb4KuLbztxTZMnju+f1bl
LH5k89Il07ERlEmLEYSHFYKEyZq4iMF6ri/FZmLXmod4D9cwf/ZhvhJd+JPUMYYS
DmBavSMDzZp7f+ay0Q+b3vkZkHQOE+abd8jVuJyZiA6N/IssqD1CdMXQk+nsJW6b
85GceQ8bEwIi8VRgT/QgzxV/EEBxJSH/Jkx+4cVLc8oyJnzwjHjUm9BnC0uskuo5
gZSM9jjO7ryKwvLtRDU7e0cjlPI5mE1O0vyrtkX73N6dfuascgrhkSX935l8sRIJ
8o5CjSfqGXCcVYD0DjaXBpH2ZJgT7ZQzJJVDtLXdvPvdcJloM7k7ny6cUsoH6+ux
lOahn8G6rPNJmbfcxxvoODK5sGcrGIxdnptL3APzGR6val6ZWl9sgQtndpvXYas2
cv/PUJmswqQ5hy2f0sXx5HbsNqOI+dcudskDVWu9Q0ShMnT54nncSra2iSe8pqAF
RLzSyGeKhfVv293H1/0/Ks+U5Z/xZPOkT1fMMSCAPosClWviGf/D06NftVetnsP2
nW6gbk9zYDccalGnEQEcY2CxVc2jbCL0AUu1bXxHydaDiFVhCT8pStYTMhi6JlMP
IYEwrVF+xlGq615iXZjIBIofC5CH+4tpZE1Ot4Hw/NHxWcAS1SsXkV627QRJKkOJ
sGm4HHYF+7ySFGEJZCan/BzNsDAsEsWpRBUYcXfujOmN2a/6lzeFhwCJPxXAD/lv
k3+ylcYQEQNhN3hxpewo39DWzj53PB2d58FvH+/SqtY8FyD7lF3I/Kr6BxXy4X7N
bUxjPQhepDlBclQFTt5V2tPV/+ogDeq+aTI2W4lW79br/5J8lo4Y0yJ4Xt6XIZdF
GPKMGZb405yLv7lReiUOsLeh6r4UHA8Gdizy3mI5oH1luxmUlbe5ot/HyzOlIrr2
lqfKiOWgG1gvRV/RSs9uPUwEgWXZsM/+52dayMdcJNTpIjoXNcxHXSmMCGLP+Q+Q
uTK7R3J+nHUxWej48t1w6mywHdf+OQtnG1phOyL8NTrRTyzBL94a+gnRZ/U0Pk1J
O20e7pBD9k6/nwdP3BoM6slRXQQKoDppcNO6K97/xlZAEvV6AnoKYfy7gvHEycQR
B9l9uaMTx7odYej3yxoTsoP6K/60CPae3dsPtXTpu9dcVhb0wr+7XcdK2h29FCGJ
UcP3G7HN8bP0Eipagu7i6NDJ6f+uJH6HsE7BmzwCsqNLh7ueFJxQtKt7bvRMsWDX
T/zg+CyBLPltt/BMGiNQmzncX2CF+hSC4EGtNgB2GmtvVfrsKvl9Q+igSq3FpjZ3
S8q+aoxuM0mtTo2wL5PbviBnqylVE7E8xlHEh6+R9nNtAQxK979pV2Q0cFpv8TRp
lWtTUojd4a2o5ZmkVggbIOnbTcbhELbDWP3ZkiSb0t2prpGLXL6U56XfkgjZyNjo
8J/gx91QlBUtBnTAfCq9KWLs3YGTA+UgZebWWluT+mirUdMhlXjNBLahnD1ZDZDQ
R9sWUNIF8zEAG5uRlGAAKyrP39tbKzdy9GzTROemtDj9DD2RZFXhqJi7W5+wAi89
E16KyAjdHMUJl5cLDd7BFexuTtnypz9PTG2j9PtfuS5egkXe5APfx8tKI9nJRsUN
ToLLrNXFjf5LL2+lI6Qb6W5ca+Ru/12tHoyzpArW9+kSWeKfbPk2dSsh/vQ+S6O+
OzsItBvVx50UdKAOn9+7E7/bIBpqJV7cDzQZJOuQVhpISHLwAlLXA3Nt9rWlnkXm
r1Rp7EBoG79B51ZXSLdAymuMWBeqPSGz7lRmiui4FXaG+Oa466mb8+vUukrfsw4k
yjVSUHyU5PN5u4BLp2saRLh7rwrFhplJ+mgmHPKPhNzQ8IIEIQ7CrYok0kkqyzaP
OJ7daBnG6GeNxoLaNVlkBPw6pHeExqZME9diGHGN95zL47JNG3NK97MoqaiJlqyY
V+YXStVMDNZeO3D/ahcUJwQirBSfgJ+a6I/uZ4rXuMcD7EnEXYFqMV4molQhCVxw
M+vyvywB+5DhJK3gpXeXDC8tm+Key3ZNtplp2PdtOPQLkL8jAXSXNHYHPrSLlAcj
e9JzV9hjfouCbpNSwMjIYNZyV07y1iDz48LZw3cT005MUSGzwKEtxrpen5lqi7kV
ian/zqp1g0uj6C+a/cpT04pfjbIh60DVkL4De1h6ar1q0p+4lHa2J0aAHv1iQIPo
aHTrDA4rkRqC4Dzf9kLlEm9AGbSgDBQWD7eFKzbHY033LnMwgrIJCqNLzPZ60EOF
rjrn8WUcHwZDF4BXIAJZx2+iUGtUWvXjOh64Ng7qRv6BRxe7By7BI/MILH1sRmLy
VVquW5WeroSSUXGHSJWk9SE2Txf6ZHAvYOyFkUHQyYyKukoX4Q+spZGUz7qfUpgQ
/KyGy/r6B3BXpgW6z0EpzRQfYrfgAjYlHV8LQrkx5k0owFi0BqV7DED/R2Fc/eG8
b3y2V4GOBab5B2H1/4ZhFNBAdgVI3tHmraAw3RQCU+UXxldGQ63yOZmVgYIx3O0L
Q298Epzj0lezarT5ZGgLl53Xg8nO18vsBYL45VF1ohUdg3QwcUtY4+NTHboQQtcs
f7eiu7zMr8uecPt7A/LYOEck1zMmn0aclyAi5C6ZoL/L0NmOsjlYNNnPqmKMMOh2
chGsBS/dSbW9x3zlleQ+o58hPJndvP0ZzhM14YFuR0QUT8GBKFAzUkIZid99E+rX
719sgEOq0l1Hmswc+j0Wu6KG0LXBBBR0Kc3KdHjLT0++2MpWme1/e++snX9PGoj0
HVyw3IV1Ls1JJ0dYnOk8Z/TeLdHHngEwjcVvz1JzMIon52ER/3Qq7PJYG/Kr4rrV
cMxa97Jww/CpevX054i0eRSDbg2NO5Bg8fRG0SRYG85fCJi49ZntMEQFadCcqaDu
Q1aIPXd0qPhAfmk918LY6pw17Z8r2W2DcFjY8395ZF0djtYk1o4JspLdG0rtNkVr
1ZHHqNyWmBkx3ZChIGWxsMx/BzjAUOqc3kkQaDLpUU/LuSm4xNk4r/a1Vt6/3Drm
AkcuVUfQPGIxMpkz/VkTJ6SyifaTplWI3Mq2QUj04yeinHDuQZBQajvxQ7rMzdEy
TV1D2f7aHRRnN7oOVvx3ROKGBx4gDsP75bhXIHdwYb0H61U5Y2n90AdjO54anOP+
aR+Cu4YTMK7zFJLrUTGsG4fHui9JyyWxKggIDxg4jaDh5dGkByu970WGwDIGydnV
4KQrShcCX+bVIZTWhUezieWzbcFWCuuk6GZPlpNIrI9ymCZJ4Fi+ZTTxIkCQJ1HT
/w2sgOA9iHM28bvQkzkmXXnzF7oMwNZMzXDimyahYbFr4SQtTnTulOV3HZIwyaqc
HH17s6NbfJqcOrhSllDri/hJRb3bJb75rnrkd0002P1XckBKTQG6d/60Ra2BwwPC
FYwR9Fsf6I9jqmEOibJIZZVvcZt0EscwwgKdvpi1HBT+nFIhoBDKls7i/jfYlPk8
hUuquAFqX+Y3/GvFmNGIIj9dtF+aRsrsx/f/MW/50IjNUPTkdmGtMJ8D1tQHpC1x
rFfmqKfoSyY5Q82ElFDoV9UVCegxJ56Rq5iaGzdDSNt59MS6q0VgOjnzDs2/Eptq
ZbzSX7TlVGSpPW78Dzg/dwmn/QBXUzly5RnYnJbOH65DALR5ObfVp0fSaTqTK3nW
E3GCdI+9Xz6lAdsBAqDKVlOM3K5JOPlPf8kg+dg/Cu1a+4gDkq+BqJn6G5mVwmtt
IBjSf8hDrTXGa7flXpaWKh8Gc502yDlbrwhG87Jw1bdraZgkQRbGsMQhxaN0epcG
sLqjfisSpr2FlZAyhPRISiJqZmk+9BumN/aSXPE8kbrtA5kvQBCafV5JDkW9o9PM
/QvnioBlgwuMesfBB4JR3fhE+CKTWgiUz4oqWwk84oLVo7cl7InpXtUvpzZsfa9J
RD7cxixGXFpRGfYEHBnUpyapdXH+3i4wX7iLticuSWorgXtrSdbiefpnFTjjdh1Q
jZGWuQHec2rXZGvaZ/Vr2VBVM82aTrGJig3B2WJrV1npxXUfv7m3jsLSomBPOSc3
2zPjUaa/RXU3LyXPpVdAT95vGADPTc7KPm5EMXzkxSE2txQ+7MGWc4ecTYqIss9i
gHWyqUisVrgfa+ZhCy9vhp08YAL04xYmixLjRVypQANmva4kG6cVmnMfUrjszBa/
DCdbXnxiaCZU2jAz7DdF8959XRYNy796wIzpTgPRKn80pkkHbxy5YwEHSw0Lc/OM
lVCcrD9irJwvRUwVA1TDYXh7M65z4S0hcQORH82WxjdKNkrjS6lg3xsJNjmzDtZy
gH/XanuZkk+QIncTKQAfuYeTnZ3RMGsNyjW4IV5+vss2LgzhnSK80rq1EG8FWVPM
53g0SMExQWdBNGoru3HhHEV0RcZG4mhAJZr/74f5/fQC3uqCYxVdhYqDQnlYhWcN
wDjlpkK5rt6g8mJuYvlntRUpuy45k3fIb77OhrRkO/zvOw8czWwCnuqri/TtU4Mb
8zYNTH9/gkLxVBL1R+wEkICK+hxYT07ADGttKxcGvhhonkImvQKCYSWU1QYUKxiu
fVFbKGioRARVypPPObp93WjbJwPLeqFOs5fbnumo2n4LfDuIgVnYzk2v1KhZuPlr
rzSxm5FGUfZRh7SASNEftGQ4W+5NYarO8bUOazpSKkLjaL1hiUm3jKwXrEAXHBaQ
+p82cMpMEl8tHdft/YVW/8qHSKVDdriQvIqAp5F+Vs0NcbuKcJ1+jgoUreg+F/9B
96jexFsNV9RoAzuzbfLSx2guQf3V3tKuRHDcBZukJYOeJQ4HdpP+4oSKUrMjW2Bn
Byj6S4jlMBKehyUlHOi8TvxpvzRv+4+RuzVphIA7dhAXQADealvIloOBMwcDenXF
4kDhyfTEVk5ibukZ7/MpftNAzpQvuUnj9uR/r2b0HjIU+uCf/3ICNnrzs4s1lG0W
c/uHwtbkGR9F63BnrNvTR8mEInYJG3R6DbPmnFRQ9JcDhFZKfVQMnmu3PBO1N6DA
V9vBShyaKLco2EwzXgadlR2jyFVa6QaMMLT6i0uc7dJa/1mtRlMn+cO+ekVGhzIz
EBnR571pS5cshO6fFP+a0l5EHUwvKi6LnANeaeORQdl7okUSIFSh2C/mdzmlmJRf
7kQouJ2HnAZ7ab0HRXvPOwGzeiK2twqoDBT8AKcxWqJYVAPrwOUJlsLSaSRI+1df
GPhUpXxvHsfUg5d+87i1ycOIJUqTJupUKpRDVEv5durT+LsdEsesO/VoEX4XknFJ
3gVYtg6DMwtPSDL41yqx1GwB/KcxN6BiHrrAYSgInr5XqQhO+AwjcIaeoQ3jggD2
k5DJiQ5b060UY+wczHS3MWYSi8PTlYHjT8u4qTPYO4L0MpOXq6sx+lF8uCAkvFoB
ddvMuLVJsKfXNKsuMjkGQuJavrSutrMnxRrq0rnbLrKtYX3yNbDYR+MAIXQNycsj
6FUmPkVWTP2xb9P4mPNQddmH+AjxPneqsOjvzIHlSTL9GFT4MgdPeUUlt75V9Wc/
i6XTdB/k6vAWps5jwyARVPDocexxKSKZBTxwiI9QjVo8/bWzUC0+Z5gVjB5Yhtug
wHGetJyVAtXaIq/MuX99s8KdvWMEBj+iPGVbOAPx5EZBBHOSH3S6f0H18HgrE/dD
xwZkVEJKuKcay3R6sOPB3HixrDPJ1apt5vqrAHKGhtFg6A/eB/13YNpeYJOTB5e3
qFhdYZY9FYVA+oPk0nbfS8b/UJMYZySf+nRF1abksrYl/6Lcb/t5DCepqsmQ09yS
qp959YTpOHzqHZbAUaWWCoL6faV/pv/GLTp8gBqNve7wwhjEuftMsdl6C5+JTm0u
CuoA7rdrxyZo51kMgPkBEr9EmPe6gfutlmZ0STgORrCGgbF2iEhD5ocRgJ4YiIoY
JkAM90UteBrJYgqpxzH6Xsv38mpIkPO3KRJ59zXBlAG8f2pOMxvxqsH3SXkMZnAy
81ckv7mcgeiBW0qz6zNoo6QdDmAwT5Glv37bCi9bKZi20/Y0RvaqfD6iMnDOIQHL
/ec2wUCesrrmL2cLxzdRjlnaaCRVsNvdfeZShkAh3nN6D7yn/JganYxlWGaRbD+8
0ih3jHSSw2S0gmHpv9CQhkhnQ7FBXRMBRoNOv+qEiOjF7m4xrx6qQ3vQ4Z99O8hv
z9icPkSsG3OOh28XMWccSGmPM1/omajPsfkydC1F/Xu56FJ/aGsjPv4JzSt3mCWI
KTXv1hCBny8qemp1JCrMbJ4bInrj9lM+qiQQTzbAOAvP37oa3QHpFLXrQKVbL1fL
Gm3Yrsa+l92PfF2MJHJDJCHzsV3CRTNUM1uqGABskqpvjajngUFDxuflZZgCMWKf
07lu8I2j9AswJNOwCQa6WnKe1sFgIhQMigYIESCcOff6pIxcy4X8cqTr5XLMQhiu
izk/wfn3m76r+uQMv6Q8SEaPad3rbPo2PJ/8O+pRfo8VpgdlpFHCTKwvpZM0WXHR
SX8ZYDOY1mxMP/GDGBdpVYfZ+7j68B4/sbXKsbAJ7Esa2KALf2T/tIElimngO2vJ
5OKG98mjBg6OvHVxAWrlLUwoisfFwRIj9IGbFmhaRw4YvCj89i0ehISz+HydvQxc
zMZ055gxd9HxH1mwzFTAyZ7tnHIT1Fo1SGmQXzBqtskw2jyEXES60isvYE1gz7pP
N/9I/1JUp7qvi0/U25xi2O3pbVKl7gL8mSwKlALkC9oSTCHLysjfnkgsmy3On0BS
YAjBa5kRE5TC/mUCvjb/KK6uw3Zb+9M9i7d9T6+unhZzaq3UFqqnDu8/glVzFv5u
FLsPYZoVkP/f11G75XYoy7VHijBQIw8n6dP9WYWfCnLynFKH1HUKDQUzNAkKQ5AB
2xdyp7AgYRy1Lt3y+yKAY5EP6s0QMJTzdETrkmwYoVH871bvCR7XMtK1C8bihauj
Y+UysElvurs/tmnD8N8BM7k19I/v3vceGUEaB7oo10tH6R79qT8xHOCh0ImArUio
1+wqeUTbOG0J0boarhURtCiV9dPanUoV453QxOBZnpag7hGxtardYyvOFtWZ6eYF
Jl3PABGqyXNQP641JExw7SKH2suFVdqVnkvup4XL2IExBqbvXbT2xjlkMX+VdINt
qrJk5UeuYdLGNovEdkxBKDCjL8QeZhtHbyvsXyP3HeojF2j9RzkdhvG5oTYLwbpN
iBPUhHsGXkBtp5SOdEUEQd+qBWgHLmHtEPRM8n9+hW3RQCckEK6k9w09aIvQ73/c
NV3BGCjR8lSRAdhP28TF/Cr6/Vmr/Sfousa2U6uHhu4mk+YPMR7FmQg6kpTiRYEk
8i497RTZTd/IX3Nrl7wevnAdx2IQ26msL0kmn6uHi5tFmrvF2ALpubbytG4stkwW
tm2lwTykBWAkNnlOpuMvOVdskAttPBUqq6oratVWIMshOMwVZHi0Oz5iyvNaK/S2
W0ODplGzeImmOfc+IWbsbu0UNxw4c6+IKM/e5xyuHh22LH74XYjpSctRGogdwE2c
I7AnpO6HZegv5A9QOFypravFqiGvYKNmSun3YjUxaWOjJI7u0Czje8+k89ZTOsjf
0HJvXVaH7G1WzzymXAJUMTiDBUpR83E+k826eerwHaTGx2di9zAayrzZC2RZFa33
4rLP+mVmrY7PMqGxfFqJSP3Et2iaWxly6tLado0tcHpwFSB4TQbNes9jEFsM+CRn
t9TANbzAn6X8EwLeG/5IHM6NBXFdAow6PcSw1GSV/5jBZrNhf3WUd2h3VkEdW33M
T79hoor7MkHp/3wXnjceOM9RupKSVseMdajUvnXWqkL/Do05/mUZyig1zaCEPdRy
4mTQqMmLNqBb76kKARPttYeYPL6WbFHrWaM1Z7jstZuKMX9T+swKqAFR/IfVuckQ
QeR5z7Lk1glqbMmgDG/1j7DhlJZDbOK3UTUeSgmLW0WwqFcpZy3ddq5d1VcvP1Wb
d9tpxXnXwzLmxhBLVvjwBbw9+BBmQ2YigZAb2bTlVljDg9iI06wmz5Uw213zw+Xr
FV/uj86wW6sITdYifoqDsgLZQfHLZTE728WDfGMm8gQ3lGbV8a1+61GJ0/0YstJm
kBy3ENvNZ6C3bhyIminoCqaoAPjN2+teT8iGIZSdh2VSfUdp8z81HlZSJbiqSaD4
+ab3ijnkuA+uSg1hW0gU+pzr408tJ7bGJU1EFPxOva0yE12UyoemrJbSSfmeH2W6
WBY8VrGt8W+4GaB1VHxa1d2Ky83UVphnCM8l141+1xYijLjkQRk5esMCuK0rOSgh
UpvnHqaUvuoF6AfD/+OKlHR4z54Rc3tacictCIWIWFAT2QZvDGp99VieWC4ckEMT
ew87+PS8mIF1+fpUsozE89G8BDDsttSOrOTjVFVu1W9nuSfvFAatmAlHe2XeRESR
CjaSkPc5vIVArdJr2pUqNGcIu2tUyNSsW0uOeweCcGdin2L0BdUm6xpCSpqcdZZt
gkOYoARoEYlNoNJZPS2L1CqGVIQTymtFK5la5hy3n6MJYcDg1BIhijRa4hATvK3a
GLTiLsVK6NnsmcaxyWGB74o7EIGajvOcGfnB5oEelTJ6DRaSWHMGtSwNEuHhQU5u
P9BE02PkMqvcR3XR34tWT/fuX8oN8vwRBGaTu4df8ohEsWVkeviQ44uAUHOyn0Aw
I10Joy/mnjQfpjiIyTp2+bYdEK1P3cpoubl68SjJq2FLM2eR6HOkwW+HULIOW4CO
XRm7z1t3TzY6MvaSVQ1BLNZTh4vC6P/22AdAZAwiQxRGdGDaN/Y3sOAQNK/c5eVM
DkKGwWRmnY8VvKR0aOUoPWxMlqNdGBC572VMn8BeBUD7KxfWrapnZWQta+tk1PWf
8UM476So6mPgqWr0OUHvYMliUyx7SvLwjg7DG2oeBMXdiG9SrcmdOVM3G+7bztL9
DqSNtcA/OtCCVn2XTffcRgBKch8pPMUaZjviE0JP9uMjXcshHsrzMH/DD+57416A
gUhvY7B12ge6C9noD8bEv8XFmSCABuTut+zbPwrTpfYd87tF+Ubqcu9aM+QmHYuI
nk0LdRKWMiec6DAT3C04jxVSqOrUMKw4g1IKIvrbmZH1v9TB60yAhpNAaM1EkZl+
ZAZ6vUXO5pqUoa/oXzeNwFIJghc8wJw9Nk/KvcF9gmdm4YmeFgceXeeHev2W2eHW
ikUQZiteLqnzMt1K4JsWShFshBogZeLP12Ws2DLlV7LILB6ciVlPO7Ncmisfpixg
BeiFrpN135FixPWnZ8HZ29oabvKIl9c6hH35uEZ4uR7LiQKVX4ApCseUDPb8P5A6
kVjw62We2KYu0f/dlAlFztr67SKdnhnQRO6YcxdOcJvX+IE4HRE8DgjlNgMI3iHK
mnf9eG/pEuCzXN7oO9QOC7IZFofla7qnLI3VwnbrZ5Sc6dHjpuEXtTE3HFQz2dwJ
4kwEX8YzbluwnIwKwvAzzRJt4X7L9xexGwh5eqB3z95/hMdzKeXT7Mm4QhnGxtjH
OlAPIc/bYzj2F6vvsz4+1pnvZv51jS54Bm/FYklIxeeNHITuXWCo/sJQiAV1ZSo1
GPsHRmBPZbm1J/RJMtRC4jYEWfKwcbaUZBNW7Tf58CBHSllffPmuDKISQ/wV6lZC
dDiU5R4uhGHZxiPqqW5MpuNk7X1PV74dKaZlejmgTnRG1bY7ZOGUIxNNEZsz+APG
3r1mUSikHDHYowtCsfVTl3/2p4uodXTo173o59rKbPKTNfNqjr85eWhyTowUbrwE
wy6IbV6uqCrvD8hNxyYhMUH1r/qtFZpEN7XpMkg2yykIU8V4dR2s7Gnrn3xj8M5e
OWRgX8vZj3KAWFvrRQXTH61Y2pQdLK63YqMv+gB5fnJUzAfmLfM+iGDe/IXPahBF
dWfhbd712Q9KbOIAZguIjMxjS8NyJq4EN0et87m2rxwUxVFDIxY+gRASkwY6Bnbx
32piSFfgPmvvjaXWz6XEPhhrcVW14Iz4OC93AbDY+nX3Am1U6s6YUAaOQFOQHTtg
ySTDlOnp7LDhsU46TIm3ou3lNr0wYFPSrEXUoNnT/zItBmAFprYT900D2f/KuXcL
RKRLdMoHVZ/wgd2jvO6vNJRcvMJXLggwySoW6+Mc0JeOQJtpHbnoPj4Rt6x9CJVL
t+ATja/mc1x7QqkGzInxmY9fr7xp2Z89oiEnin8XtcvaZqlsF3vOu3HeRT5zIwXr
dCHM/wO6fZuYNdbc6TVV+KU1QkCAeYUpFqX79s0kUNryuHfWWUDsZXYhLUtErKTC
jPU5HIJVyeMv8NSvjVK4a9CKZ54MuBxI8BFR+sYv9UeRqTyvUzV37zCVwvJuwmkE
4RUR3WlsDzLVnjgMgFRxNNhSabgArQKo3Nh6W8A3Dqmxgdx88Oq2CRo2fw8liizB
j4rS8U/0ZXGkY4/XCRtLmKcsbAvfTDUAWoRmYSp7hYAtQ2FNPg23k9Em/p1ErJs8
BqOI5MpIG+91wGVLhB/IUiROysJRPsc8yTZrUtC1GOZyXtX8KgDY07GOsliM+Z2F
25rw55pCqGrWaAw3ZRtXi3R/TilssTuUlY93OUu8J1UTuW1zt/gKXMOyZsPDyulX
l8dTi6zX09VfA/6PbmhVXO0SOLVt+RnO7sAWqrmIVR3cP/0mJ8S5z5Xp8gVvcXZd
d3VKcKu2ykxlCA849n2QIfyt/2G0Spe1GuHWZ/N79Zgxna0Zs0j6+mUASnXCw3Bd
5pl6JgQt56J4mUeXmMJMQvWU3Cj42PhW5WHLfD8yMXdqLKtOdk6WQWsf5mPxBqwm
TefCVLw0aE9jfzg81Je024KV/fFUh+i/w0NQYhQHVikL+4qKT+zM2HMXKViAYNwL
R0n82fyabp/0+ZJ9Vc5ccNUKDjpKHh+wk+UBpj26XMqzkv6AHl7bWMEIqIsxpLNG
SPwuum8WBSjeLaKHK24rLApOkrmmb5VtRFQ1Sd1VxJyXC9sHiWe7wc1kNRZNL2VL
p60NMXN68zDOpH5fH9i6QLZIAn34L85rCsD77xVtNAJbf9xL23W2GnN1K0RtjrBL
SQBtc/xuy6c/5d/cc+LRvcsfIEk9/TTY3hQQrEGSqamaDFHMidKLWoBL46wJgPEl
6y3QYa+S+tROWzMQPNxL3VKixenkke8+tln/IaZOUSTjO8jyCRNok+XCAWGkrOpa
DGJhjb6i282keWPNuAtmkNC3GpKMgbxiUZZmIJ8+S2DkYxMs3LxvoSraMyPsmuU1
96jMWnQv/zBLCF2n+r7ZNNyce7SE7168LtNODal2F1X/G7zsIUObuemve69J0KOY
176SU1HIT+135/9cRENu/w+dKa4zr/sd/2LCFIFC2FPxWA0sA0/6RA80SOFYOr1t
5IJHWTDxsWEjkHf/ad18jHUBoMhb7rbrlDyDB36XJaD0uz/ILyrC8nMgxY/nwcKU
P4DFaM3Bh/3tWPzLEwEFmaxOYl5H2Gnhq+jHTyA/U7NsPcoxQ5hVZOOlc70wHz8k
InZ1basZNCUZPLxcOH5rr8v2fwPVEAyLqcnPLtIr0dtorOb8wq4/bYl4u88d+axM
IEBDXrzUboQqfaFj+C/DfvlHL3DGRcgdn4P3Q3SFvQREeLB2yk3ftMwNsA3YHPx1
2Fk5qHvQWOEOvesqmCMkI40s9iZcyC9QniGwTVF9D1c/j1a4uhERFak2I9QcuiFP
Ue1mXvoIj+pkx9JTV6NojtHeLtW7ikaEmZLV09xVJNxxLZ0ZQ3SxMhv5Dhqa/7am
9SQKDWd9QE6jY4oyHWRw2dA5+2O1eBqus9u6GvOQbJd4q6K4SWVlWzCA1UliEIQI
2SREhIg3L8HDbb2SVrKByDRehs/FZAT5vdXa1/b8hHthmGthzSKtNy4jYEPFw4Z1
VXAr+eEeJpYJ564BQUVVUkrzC3pGYsZ2VSqMzmfKI5fSIhidYRkB6SwtVFSJ0mvS
7B3FyWOG4apfzTteg38d4m48iBeILnIhA2SAtyJdg/rbTfgWKreg/icBhZhfzXMW
rCIt6y4MmOzUJCALQUxFOkw3Ab5UHYr582hzHqkuusTPX9bIROHXdlHnO4LhwmIa
6pVPMcYRN4rCy6ren4D15I2pSjE+b7WtT0eteMxgzhCp+04QLiZK7/APMZ0iqNSH
ZIB/jG5aaIQVGHDnA6Hg3euRV0kIRAWb4xmjfqDxY+GcF4+/yxrKmiILVyCYTyjl
Yv2eQE2uoL30AJ5mWdtn7FTgsoosMKwC1Umdg85QhiNBtMgJXFiPlRh4iht7ehdX
g4dNo71g/mCXLBs9DJwlV6BIfK/DAPCjzwVKdtOSNkoaYOn3zYH27AK09z14/1zk
uGwNTFZFpSjhApQaDtb0+HJk+67j3Z45KDiXVKPq8IQPcbH4BdjIHeYp5EB+BfyF
rIYv7ciTqMYbXNWsz3orsyWLH6tZ9FcBFxcnU7FOMTbvWNVw76F7QOieaqhJctmv
2E8yVfNnQFiJkJutL9OZ+aSkskU1tCH6U5L7xfvm/u5Yylr3q2+zDoej8geOJe4y
1VMZOineQEU6ia6gtfD5mDL5LbKPA9Gp+eaDll1M1EguSCcxLng2QhtIHxy1SHpK
0v3CcJXP2ewkL76Baw412JbSRUMeqTP95U0XbKqk6yL0rXQOhc3oHMAnfa0yn158
fl/rpzOgD4BcOd59io71V4Pj0Rp7vW9ghZfFd/1ulantgQVdh1fbx+x1xt3+Ng+W
/na2oiZ6d+PtSfFerV249e/4RrdkKIMbHISvaVGO0HcYb3MouyHPInKHON0VJjMI
JD7TPg4MNl8Vh9gFN3+520SNnuCrJddgWQZEqWCUgZqOF+ByrL56DNe/p7haO4/U
uPlW7CXQpbjIOP3Myv2XuWWu3IMhOVXHQABB6saIXNWSdVT0oKjAX9TO+xfkO0mP
iaHhm8ou7lqQYv+DVMgZhRczbuAIh8F1vVVTe+MJopqmuKHGG1qClaVY6zaeDSTI
6PFSJPb6JBDhEWBfPip33SgOhPztAQ24PEdojAlqYILY4N1OUS3KBItdiPrLdF1A
gFUdJTE8HqoyIwLkp2qNNN0ry4nKpj3WTTALGEr4GqoO4s/03wVbOuMqxP0UEIOZ
cyc/E1uQLxK1LJrWKOUI5YdVzg+hP0VcbcFFIXzz6yFM2bjvwcv0tH6Mr4qV7QwF
u0tnHkBBgMP4n5DQtgnGCk44aOFJyO6TeaZMWjPIqDRHc3AeqZ4AE5fvBnmiPQZ2
a8ppCMfuGkSn9vjAz79dYp3BdtnJEDxXK6toa3jIzH6XsU4W6c01HRvkNXSOiwv6
X4sKNPZRBo7hm3oDF0LrOgi5joc25XVb9fbigo3ONpoHvzYHtTGDXZelQ1PPzK3s
uKG0eoFOqyszaQmqafxhkRtq/jGMnMss5mLdXf8OL0FleH0MDv2B1fmlONuaP1pu
RF89HcleGwCX255BYZHZp+LCyIS9r73wer8AY5j2zz5WFmNgBBHmPi6yw0Jq837b
60QKt/Yo9t+uaXwz2oztrYHW3Ags44p9oOXpl1aM2QMnJxkSIvBhnSg9Httl6+D6
WojfzGzt+TyMVMwpqO4x3QNE8nklSjxavgt70SwoCpcShuHSi4l6/imuotMg3+05
PeUbWZsZRvRxRLOFFSOHSacV34UXAtR82c8MJyukV0NEUiWNcy43JdmplmQaOBJG
p9WGVMGjBSFKccqaa2Jnjft6ygLLUs5iyrssqHswqAWeVkM+RNUXnMYyJonIizaN
pWMtSZfcrjdQBxmwXsuffq8ImOP+M6wDpDyV5nMq0EGsftmIYEx51kxDUdItn8v8
x4dHAvTQYP8gqNgnczQHNFp9L9Ztv/OwIca6S0venujegk5D4c4NJqt9SyzLsP7k
C4DHSyDzOimIDClG3Ph4XqCCk3wkt4igVmd6dBzp6rf1C2SJOUnvy99Y/DfQx8cl
Q1KpurEsCVgU4U67D2UJKe4ESUR9SkpHdEgOh2lHquXwbdmVcm87EMUepHr0LpbW
et331GtBl0j8XPinRwRMmgV8ga94+hVL4PbGEPesa/xN4OW2eE9nUMwe2cogLldX
4elS/A9YcHUyhUMJyQ+FGk0fc4OxYezsU0u9B5zVcSbX8ax8K+Y3xkZOkpxlLREm
mCQTI22ajDaEBcONJhoa52tIB790nzCn86f/Qb9I41ea61I1BhObY17z2rYulWC3
0qLZ0kpXzyJX+3HV6WXWovbrUwqclfFRqKVbDEKFC9PyVNJ8uss/88ue124Q5W3r
t6+vf4KBb1BGXnUvMr6IJYQvrIymD75JDkcuDGvzn5iMFbqAF9Lv6EcNUTSfYWta
/ziiXqZJfFHiondnWlT/8Cp7PfcL/dOA2fQOq1Db3UHoku8zhVfgTDDNbhngMsWY
5bjaKPmNwO0JKhJpOI5qfssvAUmI6q41Iam/BjY8VNL0EpVhJIihCYrBmx7qE1s0
YD7pV7QN2/zs5OoVn1XrunQJmp0KJjZ0pkCUoRM5y2ke4MbT9g5YR909ez+Zriuf
WPEwpvPQ9d0aI6uDLqMHyFh+Sr7UjcB/sV1sASpjvHrgvwJaX+WTEarssPCJ9gRc
rMVNZs8ePCQVq1PsB7Cz3SZlYHQNpxAHQeIhZFNQiOMu3GSnefGPpNcBkno+kRf7
phqh5jwNG8/4zP0zu0FhWXGy1HW6K5EwuhRhCDfbcwPfd6Q1Unb/n40lNB56jmQ6
C8boDdA61G8XkoZ9LZK1CMV4YjoFDaa4osQpXjTGoFHnwYPPXNQsTprVWsCJQ3AC
l6aI7FSC7A0G9AEXygsZEOXgDlMUGoba9kcaEXcHLD2ulKAoQDBV+V12Fc5vZoK+
Xxx33NhlBkTD03ArhwcNDKY0gC2rOweVstC1t2NDnq7a+xvCuhKep6hD3v6weXEL
KbxhCN8cXG5UdqMfyGo9eW1D7v407DuwtKKUAounmt4+GT9Bu65IlN5vTCU/cps4
XAm608qNMl0fSGWTUhAJ5WPiKa601tpK0tcbecr5AlUfTCC7r3LfHGoJBYNhSHyQ
N1MYdavvwYFSz8OrpGz/Ko3QlsBBfa8W7HEmjS1nVmy7LhK50V92ROXlKnrfPHoD
Q+e790ub/T+wNCl9cLyve/J9aDIZoEuhD/rHTzuxIcSVhdG83sL3xHdsWooQfRnl
/LL+VQVsfrMm+lKxxfqERgIp14xTw/Get9/uO35EJ+kaoK6/UuZQ+dYQM3HsdGSn
i5L7GRSHW3stMTIMGqUD+E3PCJxpNmQisSw4gEzfEw5mo/8U7722bsfZfToGymS/
976ZYp3DYWdvgvAAfHWdQO47XbqQO8WMqK5YeG3yYxY7pqlk/UVp3/ATPSLLRntu
GNrDJM2bKARL6RiIbD82H+tQ0ZFSWAIgbwDAfaSbTzcZs/ijt33bRHraBej55HRD
Tvyjrv8GGDlDcAkwkYHr0MVoJlNz4+MEOivoYyUsOtUv1tKlQhzcY1/MinHwfHFb
vcO10jw+yf5fnkSpf+QSERkKRHZX1JKml8lIk2l3lBGPMueKASO8IHyHV4z4EH8s
2rATXj37mQG8WR+PHiz6/Dsu9EA/jNnFIRek4wU/NzYDi4KpGvjDzU+F3vT33LgP
1MTWt2nSJ6/ic3+uPu9W3/YDYS3kkh0cdxuwHA2xfKTjcUG4r48YCf/j3GsQMvLL
rXIhrv0uL40qWBcZwTgpYV2GPWjbbNUQO64knuAR+rNyXnF5l5rkjaQbPO71PRLT
5FzdxA9PuxPNfC/4UTV790J8yyec9Z0KLeYGoyeYupWrxw3D3yrc+hpEsLN5F/Im
L4j1ll9Q9kYv2seewkOmSPB6i48WMJUaifu0J1oF8rCWUoIfE8oJFDZ63dXSQV7l
YGLfE1lKzLJ5r/NRtjcMks+LqtIw4bGo73kRi+kAEEiLvYLD1a9lrNQDOyg1TOJV
UEj6zbBc/ZZgWyCj3XUmV+1wGN89bxpaYO2WKQdF3q4NO69pTsn/C5UzJhysxI5C
qxJUPOA5IYiZAPsq810t60aB7igkRM/PdVgUT8puA0PIcMpAk0wR5rgs6LtfGonW
wg5Ns2O8n/2ZvmTRhBiffvRVmSHv40OkBs9nrG0yf2ddySzVmgO0dTQ423+QIV+j
eHOlr+wJKR4yk6eQTimv+50d0L59wW1yGspRNJlq0BpPKO578ZeppELH7aP6YtzQ
sn1tDvlx52tEv9sUAoV7SO60UjlBLhiGB9s5MqidU4vjA4bCjTKupGPVGVYnED/e
phscwMgaw117lqCVCtiDLLJtPvHnRsPe/9LyMW2pXAr80vsn683c/eQlpF2x8ug4
+rpLpzLQdU/SQBt9eThjTpnLtiNSCt4C1fBCthmMjuXsKJDXwgHrRiglupOHPO2h
qF8BKMeNekgtM9zxpUL+x1pRPXZIyeT7qVE9UowOFQLQPQJVOHb9bz8FkeyITtnv
I1Nzv5h2mBrLI262Bn9dK4LzlcxPT3QVXCBa5QfPtURjsEcALNrp46j7F9zSt5SW
h3C0d386ZeGlaK9eM3tXmXUCVo6u7RAj8u6E8tHRg3819yVYOVoFjc8+b9DA8asC
IfMcPi5jZ4/7iLf6AmKIBWQQA65Bcxw0qHfOVEzIqxi/F9dPLAMxF0Xj1FWm97s/
wNRhpIKIJkxRYn3WTRHoKmHUK72OEEV2kSlMZGUck/KOSMrjs45KGZSEeQ6baW5S
CxbBqpje/8PNZMZRr+TOtXxKU7K9duORu2gCPt06hQBouyOP29tz5YW324qe0ZoR
iv0JmBt+5uTij/sfr7FNdRNw+TbsiJyz3IewmZvcNOTZvJym0Telq0g+8hR+fN72
VPkI1hCFZqC/LaROOgIngmEGJPKRevpZYOpDliEWrwoWoBClGqUwFcaJ+LMzXz3W
JAhQWMwYtSDvnq5fK3tnGuYUKQZcBONtMrC3tWkzfxvA0YzEAhWClJtel4e+HqsW
ZrvSE0N8ZlNMtE2New3HeTjIn82aCa7OeEGybwzWRD0uxaX8j2zGD1YeYJ5Z166p
848G+pCyWP5Cx+5T3akNmWXFItOSGXD8AzuYvhly3DWQbA3pJXHFSHG7OTDzzfoA
9Io6lt4GIxi5wPkwgAbLF2JzQ7FCzLgCOT5RTi+hE8piB04Ne3p1YMXCnIo/5LF7
Y3VhG2mEpYJReN46KjV7UY601X9t+qfzfzfa/DdkzH2IDsdY7YLW0ZPvkyi82MIA
498tTXW5/3/11iIQi8Rm5zWEywT5vWllxFWUjot7QGTfQciOc+yU7J9MSDWzIatY
9YvI9lRnS+2FWagA9LmzbIDBw9fVygT5QLRSvxgTEfKTrd7Z1kKHZNDRlpBkdeyu
0QkUF65jIRKBqfKWZJhJtIA+0FmxSEJBu40H3BSLaM3crEXxqTrST6Aj3djMuKry
hce2MLvESbw45ti/qZn5bIGBpsPMA4OHGVVW+ttbKqLs5uGiG5a1L6Nk85WtlOH0
meSqL0MdLK+JtN5ut1CQHvZVL5YtCuvbAAskJhLLpy1dfCHdD9m6DDL7/xB8tB7u
AZlXRjRdQqRG0FlmWWE4r3QtwZcraaiQLwLfT7+XrjqLPshKVKrIS09ggmdOwmzj
LBSrXPTfd0JvtakmP748CPbc5Z8aUXGrdcByq0KAqqN0VCtDHvfYHt4C0AAe8X6N
Sj2gTZjJxrURz6pwOXK4jBHsx6z2K0JbavigbjdeLHdVXUL6PJ0BVi7eDleHN7mI
BzIObVgS/YGXARo6N0HkH31KnCJyzfqpISDuPBndA6OkvB+51DQZuAk966PXOjFz
Vu4uvHjtYpwtXDYIZpV1oTN2RJTfXUeZq/oyvHHprf/4M9L3nbH4VOiwoVFrNDYt
Y1bwInUUmIuHqcIJ4Gewwlr7pZxHB1bSv/DJsmOFly4K2qp8njv52LYxH40nxJTj
IN/ucFUPCt8drgkTUMndQ+8EdNH+jZ1eCuTGSjnzjctTuUnYZqd7COr0mPG3VZiu
d75GCRryxvcRaa163PY1fElSk9pb//PIgbUyvFZwEICHwjSF4/baJeNlemxkqZL7
jyRvpbZvrm8A0ry8UrgKBURKLOzoP494iUCQNpb5muZnHnt7tHH5yy0QPcvVuPDN
sOCsq2ywVrCBqy1wQeN/b4UXG3ee+kzGS/Zm8Jd/MH1o5oDrwEdBZIMEY0r8nMII
Uva3IqT0wICb7hAVSAOtOVz2IX1SzjCBPOsBOvhVUFumcS0KqQou4kPCUVbbJ1G8
4NSAa50X/CedTekeTyS8iaaB2w1G8Ym1GU19iWkNYk9ZEzQQKP6PZKkV8CHN8BoC
INIpJAI0B4dU7XkpNSBum40/f6u1TVOsBJBjdJWjQCOa2pCSUucfUNSH8YXgrACj
8mUYrnlLDQtumRORtZQyfgXYBlCS36ywN+vg6Z25gFVh4TVgAEiIwcynZrDXJLlL
22OKiNnuTYWyU+xkBL1DgutQOnTuDjm3kwfvQogfS1ZSH0SRDp7n08uUsFIKw3S3
Irm65wRsQ6gMhxjYPhYk3HmgvB2No+6L1KAzvDplxpn4NnSwhfq73+vLPOPXauWW
UVJCKWs4BxpWhqPYO+57X12kh3e9Bn/q/sak2CJPszRCSQXz9Zaswn45i4vN0uwE
bGb6n4UD6IOLdrEumNaWWkRXDrjaSQthH9K78J9cZbQu1KZRaqewspxlJHiXuFQ+
caad5xdGW7OOMqpP2vQbQqTQ5aUwS8dAjMACHCKFgkW2bStKoY+Y1lPmVcIdPdgc
7y3k5oO9zpyizCr23lAOTiA2IEqnCUHKPiLgI9eET31A5zQ8iF8BKDQkyNCcAbD0
jsf2/QABjcpMFOgmQ3M6toASab2F7Jd/qqt+piU35MIT3iZhsrCf/foG6uZSebC8
zWuoGCT0avJ995Wjz+m4q/ZTRqvX3FQQ4oACV3N4lOjyL7BPMAi65NjmSC7eefFz
utivQjOlenpDOHiphUbd8GhymGuelUkQwTKwyl9edu6KvymEgLlbBHySqK6jb72N
DYVJ1mBeHCU0RueiNq249Uf0lcS5lN4AI4m5mwf64xnsn/h7BRIfJBarkG4v5Crm
yMlJm5b6biWWJK9Qi3PMWe1Va8xBcCayvHZ/zrDzUO70+7hnoE2p+5e3WfwAS2Lj
rQoDuZR2gALtWvUT96jAFby6s8NVVw4E2cS20884hLZXuIL2hFzmuWqKBlE9m37X
HKIp9sWFQPnu3Sa2UO+ztz7ijex0ec5kG7DhimVScOL01qG/qYvFjHrUEC1pJGu3
Bd0fcWER7WjTczoG4cgCGJjdGF5xGbzZ4PfVRs9uztXpHW6Tg9H2BvNag1y1AQvN
0vdp3YqemB1SKCupvPpglXyLURgugwoFfHY7V4l9QbB0UqI0RszqfzOTR4wfzpsE
DtWfgR2ChIB+fhLyzcq2MFNiZdiTlcGlSiZDdvbsRr2UnXMDtgypHit5e0I59Q8h
uPyOUbfyTwF9TnYm70EISLTxoaYPzEboK15RKtaaryosFIpVoDjFcN6hGle/4pa5
kfeobJkc+TbA1mwXxgd2emW+GuM6+sFL+T5HLmnWKbQDsjIVW3bXV1i1JdT88iJn
3WFnzDi27lmIim+K1pkG0ztBxGelzNrdmPzgysOJTJ1dlzdtL4eFNzgmBp5z482J
vBGzHDunIa1nLoidRyPPC9k4bXy33fhNo5l4zb/Rk57QI0IHrUr8OWEYuZEIV1mR
QaWa23vyOIrJMHnXQRL5k44zHHPFUJ3Kuncz/r1Wtne5CS2tLneedOTKWMzdkqAg
KCge1cpnHEmbIaTmNK6qMl3uKPpLUN6WQ2A2LKxFXzrQ7c2y4ldTzGClXiN71P6T
QydtoMqCikEVmLShtBV5noulWAPuZNGqTmo9vx+slLsFoyb6ngrnkuy3uBDb76oh
dzd3PK6aGEQWA/2+39BmErOT13HQ04A+58bFj1i5VeJl7OYoG+NjY3UPEIq9EQca
5sB1NdlJP7a58i1tFdFuibs0+xTg0WBYCO9rC/2aktstPvcEPZwtwgf4dPE4b4i7
TIv6oaKc8c6pscAbtI8ho10BqjamaFyqIT5+Ev581il/PoMJfTRauoLjSvvugGVX
GngrqPjMJcpyP8MBLoyb+zeiMvu21g9PTfDbveXpBezoBcVaZSB4e3dw3W5HCLXF
Gu45XWywZgm1nf9mIs2E3ZQbPPCqRpMuRHsf15IKfzATMhcVLi0lHM6zgmxSePa0
Dyqf7vCbcXZu6RyGlMMa5WslDyKF4mLE40DLECMhyKKIPDCwZGlFT9B+qhHCnM5r
gA7WHoG2jTdI0iv8ZusR7riQR8NDwyUy+nNiu0tnmUvBZmYCSboh2YsxLIxTJDIw
XAP5toNGCnlxYwfl+uD6X8SULGdb9m5CjM3M782r/BFPRUjaEhl+k7oQlfyvFpVp
xXY/89/j34VoKxnQO+oUYz+ldKIXXQVk4eUt/zuzn2ASlHgmVlWXKiunHHnJnSkL
NilIqmhOd4FPfnO176yfEEHa70oPHoDhNbdrpJ+v3YBQ/+iov28rAiUBhOkNQ1mc
bN67Ptxinn6yDSQVcwPJWGjOJ4RhAlh8DQq1REf1xJ6KMiL8e2EfLMiWMHRFvSZ8
nbPWW/alT3GiPIHdWN13Myf1Cy/ulDihka3/RA9BUskeZqpMVHrEe/J1X7jqq9J9
nc1158uiLX9Y8RhdrU614yhfekM7efI6KR3XPz7hHq56ufvG0izA2e15Hiem+w7Q
FytYxAYwTnfnWq7LIT0bOXVUdcK1JRccWLIS1RpTjrJKYRiEWDC3ZluXB/LP5FB+
YeKDRH7wNjGu7YUbYVEnuLEYDh0k7WUJfqs5sfrQsASmz3BO2KCZ7+r4JaQSYQAI
62x23PmF0yJW7eFDpnCwdYkUryeQWqu/yMbehfrxe7v1Vb5X9oGKZl0QOZTzef09
2dCGZtCgSsWgQLJeabdfgOIg4xVViDNlok1Iy9h6K8OTrbHjLOJf+jR+Ghv61/+U
VHnVNlCLPxLCh+S7KFW0PG/yxCgC4peksnC/MbKAnQimMt+NHZwZDhIMWq+bLxvt
iKg/QrdOn7qp8+VrR+eb/c8lYhFLKYjlRwby+LUyVvfKcSe+8XQdEL7c8Oz/Qnjg
lRotOeOzsBPk33RHY3c0CiHKAiGbSS3VBn+Wn9Tx9v4h4OeBgX6GGzPhxnH3SD3n
l1igLsbjPQSowDo0FRd4nDjrU2KwAssbOEeJJECqd4Ztw01y8XcOPU1oCnnyefy1
+U9NcmKk0HFDMiwQxrUAc6NLD0P+f5IviG53vKS74Dm4u8JSVOiqHa+yff/Sw+88
z3v6Gk7f483CazWc/tZLJCY9CwtZbO/WW1oYRDgkNgCZYxdbbYC0qmd8V4XyxBoy
gBmor2ECZ+8XbqbndMONWkDa36VgZ4nBkw9s+ePnhY11VvvnBnC1YK8S1KOy2KxM
IOw8oSJHG4oSkqGqmhYtqPuiD01PH4OGUftdQ9imQho0rMCfyloMpwX7HmnGZMmc
xiYayiS3kD5ifoZs7HwlPtuTsRqcXl0G6XYtw+ETUMmnUkktDih/CzdtQB1jEexj
dZQ92rcj1hX9eqkexQnD4Xj7TaYbjfZ6YWk05pd0qJ1aP55atKKj4quY347l9uY2
lUDfALEL0/Gb+d1Z2zYDffsY0KmVK31zZR2optS7iFAwuev/xWcaqM3rQXL/JxOL
7MpMt/pc01EmnyAWlY9x9utW8FbF29SxgY/scHs6Oc8xv1c+tAgqR49NLmqublNu
UYYYt/JG+l4hB/XqwVg+GS0+EXUtSV83uOPZKXRJXUtIXkQBW7EdTsB3BkNEcKEA
zoheYP93gHeRw3xbmjmG9gmkezjsrzFR3ndtyNbQtGxPGu8E1bTbi/D/Xd914gDc
OYUPsva+9hKdW+QpaR2nT1cyaiVFC/AxKMV5LpysLHGu8zoit4wduLMSZ/ZE3y05
YYb8t6DEbHqMdbtDJF+Ur7lKwoRBReu4KdY9eW8g0eHJsAykwRltYPJ3x5YkInDF
5v8Td2LngirMBoK0iemCfP+53c462e9ddk1JlNEEuhTbAXRit8XYp593zUGU+YNH
tjGaEPYlHpXFv5NNdEc72UPFUO4kW7V+hRUryGpLBWUDxTFsY9rYJYuCBJB0etj0
xjPKiRREzy9l6RJDBKf4k8PIMjfrFofrGjH8KftooKTs1Zlkz3vNhguol/XabWax
/XF8OIdmpZa5NVeqCzme9kqWMMiBacpHpMokoQ0rQSWpegVnbq1Ecy6/5PM794OH
Ms1TYpowmVMIedvV8av0uvSviUhG4w4f/0Qi7PBWGtJUM+du0L9RA+zVlXBRu09b
G3BzALVZ5D4Nie6I3cu0TtU9VocOv0TVfeN4s0GcaQbRalkT+gMlf0FHQAgPrg2X
Xlw18VCOsoapp99ECTozPhf72qbiSRtkVqxRZCDWDEH9XWYLD/GLSM97lYOTQ3iS
RrYAeVNdR8rKDqm6SuXn+Q2KjSk2Zc3VNcg87n2BFfz42U1QrvsarNNia1zh4h5D
drbtcwT2vRi3uYBnjvvMOzErQYEjNzHG9ULISCqP7WfCE39Ls0f+4SUtHg9BIUvP
WGMZasrPJd3aPG/jLeDlomQdZdb1bjXYhe/DxypNf0tQMnJS39fajkUBfKFK0dLH
na1BfCMYNe9P4vVHM35Q+rzINPY9EXRWPbZNFsmrJK4Z5vnB1tVfZAPj4LqCpcyl
WvWHfXGsVKnkBcOW5hYT27VY19C6LzMZ8Q0HUQb4nDkrSJbj0jTsPse1ZqaG/1vd
vvOJ1OHC70nstkcIZRqonuNwIFIBsLt0V4NjN2JFI+RtAaYPHlkJOZ7zUyMKMSii
ZVHlxgmOjj+zkHMYA1jdyetsd1jZbGVMy1ifzwLLwpDW5LEuPegtjNi+QLpUjXlg
VOe9N7t6HEwtoKVOsrlRajfWHBWn+n2cX66jrqrdC+pLyfHXtXJkP3AjTio54iHy
qe8uLsMqAE5RAfsDOSU9B5U3HQ2nUQj3tfd8mVucTNGh+RyLNH+p9D2hHUsY4yTK
KPrKiE6XdHMYephdvkVBvgYdiyf2gsr6xxivRuOvVoMat/3YiI4pHTJXRe2kcCio
zB1X3nG2ihDuG6RIQqMoxVss00fL9tkSMT0gbkcGkaz/OViza01oGDwSjfkIqiR+
BURlm9dj0ikXQO/jgDCCDLNQbR01GK5O8V9/P84FcB5IJk8t36z/R2P4UwkYB11y
X/jHfGLlKR+6Q7wGmdt49OlhGT6+lEZgACgc1/YPB7sogFMtv7kp4bkr8+W9GOGy
ps3uIKGZPAWdZDMI/DEf143/qZT3mMV1KjrjRgDmDgovzSFAxVu/chLqJQOGpwMs
eEoPiSK9sGzC8AauPXDD03/d9C7s/mhfobgXReYiLoVi+LzQst7HzeWHKrXaHx4O
ASQA7mX/mdOFJimBoQZwATXVlgnHznryGVNhIyv7PdSDjwqpzP+4IwHY6tt75ePS
oMwalQdZiEp79mZIQUjIjhmXpwm7OaCJNoCQU1kmSTR+dGuL+gXk0R0S5KSNG3jK
CUpAG8sGuNQMgQpLLIqbogiur0ikhcpI8TAPCqMsASUpQ3Bp7Z4zYM7MeFdde1vm
XQN4J1HnuBAwO4T5MaPYFgAGMY37p5TmRm8/y9Y/2tzMVcX6sGj1RPuS1a5nSOJV
wFhvkUEXpCROsRrLgcNndksmi/2aYmp+2qJJ9LVbMgp5aFsTe0dzKqt5+EF+pdVf
RkT/WsUIWM77hS7FuvWRA86Q1ABRwWRKlNrCsU4CSjemaYOq9QUkFfkPMXbgzhPv
ZMq1neQK7fRES3Eu+SUS0LL/3PO3xN5/2qON0Ic4Bdf5dZnnodNA020zGxanMONp
k+oqH7fa/Ml/WZQHGK7P6Bomg3UQnEMt7h53o39FGaEcN2ESuoNixW/fcE2UfZKa
+LpLNkcSJcoIR9SlAbn3ILetSdh7Sr83rYhbKehlAhFl6F9qPcFoglm/iPpSwr4S
bbll0pyaHkgcwAC2t0w6BbQagnCGooKJ6NjO3cqssubJk54gWwnvLKqgoLbLBu9P
n/xybWeNURWo5CkGXrYLZ1nnEeQfqzYPZGjJEf3rTiCX0rYccbSk5zflchVomn/2
TlCrzh/OmqOOEEapGDC3NPBfma1dcw7pFqjYQtLe4hvr1LneE+22TSkG4xEa5TAJ
nKuvGoHZv8qJoxyoo28dwfTX1C0W6hrjHuTVhdpdkm1lb1JDIGJBmPOIiPHqFvfq
JAPsfqm0xGO51iVX48DWAUX/0T6tXMl18vOq69uwZ/IVxD0YjMwtqoI30F9MtIpK
eCm8g1A0ghlQbtJIvms80enwpuqe+VsSgLi/od5AnBwrtYMCRW/kfgC17+VdJvOU
MJhWgamjKGJ+gkcU2HzHzJQ7EdYvYBsYIX/eRcojmVMviONE2iZLEGe5JSuxHyEZ
DjK0l8eoDROlk+knXbzHK3UKCV+QRP9A6BygwQS3mTqHZ6OiweV7MlYz7uxkS4OC
t3+0KevOaljrTkpUfPh0je/ZjFFBsdviNGGDByHc3Qb/Jgxh8tbBajV9mcofQxik
avvxNduGFpktlX/2t7FnQzPzvcsWQR6EMLmNAPyCav9P+iokP9hSmqKvbwQWDm9y
QiTXNUa5dsGipL7Gqxw/7EtP9gruBVzqqf0PyW4MmBhhWEB8d2tdQsgxuytrCusK
MjyevMS16gWLMNrOqSW6of9XO2DnrD279FfCgpd84ay8ZKtY7FxYGctOE0ucOu9K
RLuvw9FJbZQATni5RU+12BhVSuWBHTs+pembvHkKdcKtWnHBQte4wGChL+AEhE8s
U8iEkreJt995UGoWa+kUXnPxcWVWrrR+t8eyop22ao3sA3+k9TEXY25AiEembRbZ
HCKrSjTsk9+Q0m0jitKZObcSfa24NL6lVwGrDcXpMuHKpiBM3VkKeGlXLeHDkCjM
KS67zFMQ5zAkaSxptCtDh2dAEP3E4sUUTOrvnjkoUCLXHzaRpA2r8Nwg6GZRYRG+
BXYRPhQLyJnrQuFL6r7VC5/Nez2OHbaeeFanRgMVG2D5DzQyNv3TpPQYLv+/EHhG
95eLjxd2CpQO8jRS6TJNZ/fyNWTQaKzDzVsVsN/YpvrRNKKHeD96w7UChNtcgHyZ
CKJWyY+xaKZaRExFFBmvjxIKXAz+SjMmB6zb7ZkyAffcfeWF3ITDyT9Ddtb3Aa5T
seybyT/OlVmvyP6ji/bSY3b2OjiR4jkeWToVm99gjITTELm01Dc5bJUxI1SJyXyT
84N4d8CKPgwiIXdjGzWHzg+CmCM13k+AaNpLFVtlrxLlvrvRY8DzJ19Iq06uaZyZ
mKOOxxJtMa/jomqL1KbNaaWgGtzLfh9GIgf3KiXiVimtFJzpePlPRR1IPqF4cpo5
bG1uCoqWRwKrXc4oufOc8+3h67X/VBB3IAgTOYzDk+p/Fx85EOEfuxHHNz0VH7WM
nvZMNlyrtqE31ctY5l/vRfDIw/GPePBNY6wMKmxBkBS/SF6h79An/7Mzqsr6sCz1
LMTHUcqLZt2qhbAm+zDSshHsMCFWR4bCxfRz6etDOv1hw/JcuhPtThbPCS4cgvYQ
Lf+ahta0beCB+/uxISE5I0aCMNKU9K8+o14VBlXZWsNBw64E1/5BBnQQIqGsq4hK
iXWt/dp4QnuSOSCcaMJFIH2fLfNvdDbFu7VyetujVoqfNs0hM2BFAoR+x5yZNG9j
MA/SnJWEKeXMJU3shpK0Wol63WZFOmRbhXfV39X9KvGxsaefUSRH9h3dC0Nu5oxu
S8vdLh1pQshPInpbmM6tQDNJYSGV5phC1NDupPNiiDxV/6xxricibINjkmcglb8D
6p/rHcOHNjg1LWS1M7g12viCuJ0BFCbkyhZShpqrBkUcZ363yBlvPTtBfQ9PmOiY
2a+igsCtpvSKQJBMVCqvkGWHAkqTdeukq9nUjxj/y5fZ02zjdwpXoEDxQGMRpPTu
bCVDaGQaZ0Lh9xMQE11od5GwP43eY+kUG7bw1qvLdFYS5vSLczasbC0nLRvXRnfm
ykrnAly0YR6JA1jCEV6Z+JFvmnSzCBHSztQAQAT6JrgKtAWMHzcHlRwKKGtV9QrK
otzvAgz5EXL4XkC8xty5pMIwbNMMlXVCOSbVD2jfBHl/vD7w1mHSLCLkUlnAzLmq
ewW8hSntSF8+iwyeI5vmB5KjP5I6bGypRenRTMPmHLzghoAqSMIaTrT24RQhrreU
3DcDPsY6DYKlliNpPykGMJmXnb/NVggLw2NITV1BZSnNgqRgG4dJUI2wO4bvBL9A
uWu5ga5jgvf1SEEZX4BWqNOqh0zOTM6rmTiG+CdO1VuL466UydF3/mMdgUQDTQvg
LdgXiVd92HuYT61mTJrJsPFXghyR9tcQLUXvajQ5ct8iVcGiigxnexXSExPbuLZz
nIx+SzMqvD3H3/un2Bufzakd3OEHl0/6eXkHCQ8eHtvFBX6lSZURT5bZgfgPKos+
RikThKAc23N9hFzo8Am+qaOCHcDF8I0OMKZWTajSexdcoFNJPr6v7QVzwgKbb11B
w1vbdiadT10nrKvccXxcRH6hpQNE0CizIBGWRDd3x54S/FbBMTEh+bzuxHbr12RY
TBEQK4PRgtc+9vJXx+NktgsEiI2iZhL6Xs9sVypjBJLRELwL+2+Q/iwBW0iI0Ukl
HjhEWPCpq+IHdUt/M/Wb3eLp50cHs4SRNQpQp6hHDcbEb7L4fWmzDywhQ0+7LJ2N
MeDjbkZldHfN4QuSbAsssmbGT+NCkLCk5PWnls5ZkejPiMCLiKUHz2MJJFS2IrL/
x7w/0ynfFVBMEaxvEiSXEskRd6mpv+3RUj1ZxB7KFhzyJKhUl/q8lFfT0XYkhU/1
YdIe/7gIjmG+KX+QOYGQVpOXkutYEVrd++Bs+LFQAGtq+1hFQb4WvS/o12qzrSg1
3eJQmaT9uDGnL476j9WVmiNBsiPUQ44kdnVWBg29BobNkUjX2hQ+HzvgYyQLkAHy
81yWRXlv4RsfUtpPKeefnLRY5hP7LK9ar7+7oo170Oyvpt//TMLqKUA9pLiOJLSs
hIE1Mockd/JB5l//RPNq/X3AonVoLbykptcVAfE2mzc40GcPxxWIBcjTUrp0RxUJ
0nqYVhrgexYhIu3CSgIBgyWPRUlqDn1sSGU1YqhMvfMZxU3j2/tBTfotZ24fgbxT
OXiWGFLJAXy4sdJl+fpeD7YuFv2Z0aDH6Yb8qmlzj/riBWyjmMGQvlsqDBrXvC5w
dZn++AMjyJB8nD0rXLtcRWsD34aK3HCycwCnEPm8OeqzRJrVj9AfBs552ik9paxD
8qC8xjLAZs2y/pgx7tHpdqSbzIiCf+p10sI7RzIlz1z0xcwF9IQKaKPTF6RLONbO
KAJ6k49SOtaCp36f2dD0/5ZEdYtkdJTh6O+luS3kYGCMhJ0rfH5tTm+hTpKczYtT
qT87tLA2spqHUWDrocyN1w6vmuVlLLm6uo/Ns6PSAs8kQb6M0vPW7fmWbGjbofYs
HQTwRCYcqo7+BjKWet+hopHjQTveEhBJi/nT2IxmLnGb1ItsoqFV936HsavuilzP
13dl/Jm+kstzm+BxyzVAfkDLu+UmzpF325SO96CaoEXFnd2eUg0JtcljGR8YkuxW
wvp429785D6CsPKPnxOz4ZMrw0bbMQ4JHtHsVA/6LdAsT3JlSmSM6IHWzf74eSTG
soVZHt5iNn91P1dcaCtEbmTpc/V5Ny5cbrTk9Qqf0jgw71kAmsTiT9D9LB3MIu+c
4SDtlOfKgplmmnUSY16DsXGD3VKujZYyUn6uvkEbSxTqZ/twjoA2n1nKqgeUpi+i
2zNfIOG/rFxKhh7dkGB/Q1rAbknIxsavs6QqLZEUaPshkiuKm4ef+zmXJpKJTA+l
25hdbljpPzDA7bf9PykRCE19VG62ehBAu/AigUSX+sQ/er3Z1JsNF2ococxntBUG
pemuI+Dl/ufFR4NKd4CB0HJwEbfCtGQOh2/4ow4djfv/yQIcqTo3c6WaLTv1P/FL
wSOcEODy9+WFU9G4K70yl5liG8k+R7cz3314hv/BnNIwnuWiCErft/7Va9ORpVg2
EwDFPaDyxEgPH77WxsHgxcXMoMyMKgDcjouL5JrO5gD02pOHOfIIMCiyB9fuMQV1
HanObL2KWUy3eAlaNIj3VE1JhsVux/OGA2VDvQ4shl99C0iguK4Un9tAzHRZL1xI
cpuXmHUW+UbgGWvKQKIMYqhKix5gtNzl83ZXaCCy7qvPEHwp4vvsO15CQJ7yl4kf
tleck0pT6XpT80TBE/nZt4pZsqcgtpCKVkxBvW1QSuxXo14KnqTo79L/oXcGBa/U
Z/J8lkVtcEvmSZ1PsijU4lO9cY8ddgEShCZ6EnIDDos9suB58Tljco8K0YVfO+Wq
ja/LvIoIVLGlakKKvN+hl+rQT3I+QiQ68fnKgaH6uC0qdQXuKkn8lqVG287jpzIU
wgZ5d9P1ghoKwwgdhXFdhriYJhWkqfzVMf9HbxGxEnGLx+F0sWH3+c0EVYFwGDKx
GN5O8nnR+h1YK18hMP9KhrYgL234MnRx3YfShx9npY/Wn+BBeWiH/Md1GxBAqgpM
ThRE9i+/zhT/cR2voRpNG+1EN315IMnmw/EhxzBAvIyAHLlqpRDZkvQI8SSUvJhu
f4HUetmMRL/f9VZIuILMSe26zUScL7UCBRXqLsK7lbBUtHXGDNkFnKVigHXBjWm3
lRU+Tgzq4bzESiCL7ZVP+BQDa2oDxAVgIXKSHt8ekrV62zHtdt6evg7T579JRvNX
/LF+MbO1k8AY0BHbD7C63Or9wag9lHskQIKv1JXCb1USmMGFBRCyDxb6DwgywvzF
FUi0jN9fJ39OnH5eG4DhfrVVagjlIrm6yJq3FaBhc8TU32LTi3IeqlrRZbrYto2r
s5vrWIYudDF5Rzmk8aYeMH8c9G5IIeoXsrufigjrIaH4K8Io0YL52XPJn124giWc
J9PPC/3eNtdXQ0yOh3kcSQstm1jXQ82KfPn9IS4z5xonHcnEZu+GUwHddbvjbxNe
CzPbslDq6gv13ZaKj5SvQk32Nfj1suRR3IR+8jvdNFW+4gzjvxkRGjOOyT0azdrV
8QSlrXJLG/7AQE5WKBYr7kblPguhYpN312kSGXDUmvwml7p/nJAzSADD1Qsp+Ojj
PvR5AiV2GvYR7yCUx+W7HWakQgDtLcYiGQu2FU/rtR+vpIEJ9p4wKu8hcZ1EuCV1
Qk14bqFSpO3GtyJQM5yK/VvHglscjM98km80FD9TROkSEEgCw8oJeULPkNG/jnBk
Ld4wRvMKwl2cgzbdKUUcoH7vFOqQ80z7/B7Q8go8+V9g5Wy6yDLLEp6fQ7pWovTh
kp43pOKtSyQOrA3p5H+kibUorFKR5kFGhAnXH/0rT0InKTHj06Km7djXc4jO2QRN
2thy0FVSGKIuidgQtY3fFgKlEVR0ya1jOF95c+brAUEo4dAXKhunLMYPkVcYhTtA
AQuyxlIElV0OZzzNA32tSljqjUxFoVhkPtl22MprbyQAWeU3ZdqZYvLOaVslyGvs
8I4NOUSQ+cMCOBPItx0KQ+ltDTcemgzh3JsgcrkBIRABOt2TCm+rbtLM6mHHCmeS
qArjKdlDawVpD0mGWHhrHk0mmmpbqZLHl4/l3uUChrrLKd+MiMHOXOE7Zmw/P2/6
JJeZE5oH5ya7kKMjkBpaqo2B/W6CTUBrq7uGWzm7dEZFS/Qsa0qIIq0JM+K6yxAA
Zsh7JBkWFy5VaZBV6YMVEWyYHRn10vBkmqvtJcQnWl3Ha/4HokwbAXm5M15an8bh
+3RzYHCN2QVzhrtRbkNO79o3ER8K3LzlX1nJ3lA+dxQFjq3zQU6O8EVivyZxDO4Y
pjiWGuiqfdtw34YEXZc0Gn48czDdwkfIf5P1Y4HL7edv6inNpnVtbSGxJrE7M04E
Y++X/BIxndEhpCAH8crR9hl/CSTjqIKXehuyLrsTvYxFiZEDiuGi2as2JCQ7mQGP
Q/qYtBkIDxTZdYINisZjyD3OtckE7T55uf1oPXghtCN0LFQGmbQwX4ttixEoFCbg
hDRbaCobrXukfnXlX9ZD4B6MgEBgsC6BiwAlJVewpTtQH92IXdBAAq9B1wb5AEur
Y9/IPPrqz8/fpYU9zdb8QDh9/6Kx4V9wjubhaHetzBPOyMchUdmv66BZgD5GAWsJ
9MiKVbAr+DRmjr2spPrWeWQ9HvD9WpnlCmx4FtxLSHZcjGaPXGo9cBvINcpjpTJQ
U1dJUm8v5dCV3S1UEYejRQRdP7MqaFTfodQLpZ+ERg2qwh3X6Z7EaKZA4aD3rhPe
8h/BG+ZI4VMmTzMA+T+VJmkpnvYCwL6wnDp2I/SI1+o6oavF0T7KvlmmEYBrxvzo
KuqHEwiQW1wnRr7m6RHKXAKbKE2gROw9tF6WsaMePU3VW6/vQ+1JUsVxybNKhrwi
twkS8oltbUIgG45Qr+ZcR7YiyFcL8n6ooOA3vvNQCeWdi1YPIPz8kbHgCZo9PcvK
5Nacei6tN05IdAbNpJw4UyylhIuwRFYOktlrsZ7Bd/mIuQTK6neDV5wuQTpEWPfg
4V87z+T1BS/3e0VP+qAMRFGCJ35isNfBpsEEgGEkiEBNZJLrukUHLvwU+U4ghtHP
wmMGbbc0no+hvXIsfVrKHJUwVfeL/s6hEyt5ZoaXYvH1zOM0htQmyCoBtRhQvYUu
uZUhXRxFULoXMx8UdO+bnECbElbdLnuc8w70Apr+iGBYYRSRL3o0xgjED5dOoeHN
vjFrKdJA1kHOoCfO4Qn7wmawVr/OMYPcJHW3pKXoohry/DTKZ0/hoiVWmw2iDh4V
6qkeJQOTpXInCXY/A/5qTjalZgL/oo6lfK9mn8PX+5XLasVuPE3TuS/YNJH46ycE
ZvqJi+oCoOYloF4jbADgXbVfeg2fO66Yma6/oLbMCR1TLMwckL6+ttj4/3yM8S62
OcYKXHd/pxKLKNk6wWTbqgL0ua88r0Bf1Rj8PWxxJKeQujnYO4DD4aN8b2XLFwZ4
cb10s/zApO6LOsP5mVSBDv0f9Mhk8NetjzLFA8roInj2OdEoFpeYb1q+yOfBke11
EuidUmTBRvZnNnoVdxtRFybRAQzSs9xemrznVKAQR3y/IHuzjSzAu3XGihdZvC/8
WJztT7xWvPapEnXcms/xKr3/zmCXkrjM/yET9OCtAOWScJih8+uJMJSKNqTnPzk7
6fFyAS6ITHoB8XTOXOMYibk5twvsJTBcgzcfMD6k887d4PFe84IhIIBuEegzvuVl
4NR/UQ/y+eSLF0iSPDKZsENJadkBj/838Um3m351pdgS/F0T+fEIrqWmtMzvpRgM
qbNNbtr9SsOhAkrX7iCIXpBPPx1py1ZqotkVD5NZTVAI+Jyc6qC9Q5TOoEELWiMt
+vFOKaGsfXRG/2qiQlZ4DX5cLqLebDqusEJNfXCKz+8QwCcMLShsv1vQiQnoHm+e
fws3k83O5/Z+/9Tk1poXp8QqVe8tNNOJoCwA7zbqvQif848/iV7j7XZkWPY1fT96
Z5bIbzXHu+grwNQpshyCpSEzAZfIfIWg+GQwxHXfvNzfF/eLyQlwzTPHhb4uUiLg
GLUox9DACy0Hb+1TMgAsKG1wKbI71OLBylyETPHaJTDYM/9EN72xq64h/FYQb0Pe
feUWAaA3EeEOwUETesYW6EIEJK9Ron1QD6+jndn8qzv+Pu2SZp0gn/i9aP4psVx+
6EFoC6jgFyIaoT62chvNlInDpjt4LIL5XtQ9qEsRZUflwx1TcxUAF3bagnMrhUEp
3CIshJjMSK85w50KItdQ8UizoKbEd7sQQf1gNKwPNgAEFdBc5iok8NQE38gIUT+T
P3pflgNCS4E/Acx470AxYDQpndeMopP1zuHhZtbl3Dm0dw2OAFQVDyuZFFzprQKV
L2erXwC0ucBZlwVAQTU23PFUnEWw1Q/vFW/55HV5Dn5ZxywqVSmQr6mN6wOwYKDq
Gnl8cmyWciHJ2YVd8GHgZy3Q5V9dAaS3lfdWCgQycHSZtrcCNK+L4ni34K33VP8c
SjcQ2ZsRmEn6lWk/oIRF7oyaHVaizIiPFGEsRXAW7vXZ0umr5IbCwGXJHLx2WTiR
4auoLi6G9fctXGfB4A26anstiLFSECkQDtUkBBrYkRc2tP7C2oVF2hm6NdaSSz2P
NmWZxMkxS/BZV4mmT0Ai3MVX/ItdPrY4lxQfZEixr+7V/KuMu75V1HXk8viRkYF8
hA0TGnWosSTCqFelcyMh6vEunGGePiTQMReOb14LaOQBmK+r0FCZaSr9IE5XIGpx
uCP5oS9YO87NYMmIukXfsA9KPzXFU6QBGOZY4eMiz1Rtv8SHbcUJhq0Qa24i38vr
D+l1UVNiMD4uNu3F42EMl8tl8ZfmpE5A4ygI4cMa7Er9Ck2mIUjPaK3t82qlhg/q
tebqmYvgTXxJ7HQ2Ww9N2R7gJTY7H6KHXhfKEj/Fk0/L8XiF0GMGlb1WKVuPkW9w
ta3SO5KzrC7OP5kkhfzEoi5evNuecQTLPmunV5XxDSNXPq+tATfpVVctUXeZ0HRh
d1jzWo+didfue9mEBJ5RIgcu2ObkYIcOZTfOlRxW1W+AhEwdY8XidwcedrObZmXd
SurQfZShwBtj5+Ck81QUlrm2xcinLlwsJKXgTNLm3fj/G+NDLyZ6oVojr++VOlpN
0J7rVgAlDNWlT2HxZVPUispi8AEhhU4zYkHlnkUl3HES7vEcfpqVGq6Rk7u6SI9Q
AUcOMvCsFQIHbi/Wxuk2vb0TitUUvnxQAMesKX9riUfFV+OI9OA/hlZdUEyYmG+v
cXc5s5EfvdKKoflJS1EENI4BaTJ6C6MclNiCuOw1Xy9tIxFfYBZguBh+zargwRUZ
XuLp4OFwI/WWippnemLTtI8B/T17ibZsao/cDIPElxz3Nst6x/sQH+yXYH5qGBKm
VKH6p0M9fljwazcH312KqfpjTbcqeHzY9giH6myx5XMMKZhOOd2UWgND1dvzShos
Vd2kwlmVN/Tr1k3AdBe3nMoA+tzLRyrk2m576ty7JpZLXQJOa5p7mXrUQo6Mm00e
zYG4PAflPm9RWGlH/IEDVRh/w0vXlGgK9oKBk/EThPXLX2pPbBFWNYzqhTKToeUh
EvOkWU0xPHe3n7OgGxAAzx4+cry9W2LOcjt3kQVn0RISe+Kiv7aFCH1q6vRhJePC
UYb/pA+8+hQfpvsfw62VwwmnVLRmWRMZoHAmujyLjmqpEHM0EHv/AnTLYvHxX0Lf
QBC82T0ZqrMBaqaFzHa6a0vdPqTKE301U/RaIRvNMl9RnDBi0V2uB/m9BpLlrshH
GU1SxGvVXuEP4wV8G36kuZ6RDbRNdmwwDvDw+K9KviTiA7ZJPS0Q2mPJbUmy3EgO
n8S4pbpHR4jYjmGE7DbsUQUi9sie0DP6gUDSNYP6zvBbScKxF2Vtz7dA1wbs86WK
HVJhoy1GllQaxnVjd0cQVLrfNS3nyqpDbxFfsl7+RuVeJTjtIUuGxcl1h6f07HBo
0ReqMJR7rmCZZqN/PPBPzexpxVgaBUnvprWLvCSnrwGL7b04pjfUB3Oobf7G6L31
FS8O/X8wPcdA2YB1/YhTDj1HWg2gcjU1c7AfHeka0FGtWk0MABE+qucsOqYOdXbU
kdPVtY5BfuQ8g5CWPGMKBSwk993PLL1S/kO4pXrilZKV3vFoOH+++CnIKPnx40H1
/nbfqtoE6eSdHBagNU13fVckteVxGmkW2izCJ486NEvrnb69RZhUPjEbr7egrsaz
HEXWkRlH4VNtlTkbE9CSOYUYzFZ4WuwUD0d9oq5h+Z9z7xCJAcXjeqKREjkW1g5f
07Lr9h6N27+SaFRnl9SH6HPEOUldfOJsVEM2JSxT+lBfLe6gEsxW4Zm2i6gK2FOK
du1+ps3kbjtK74hLi+g5lJRRIh+bouK180VtRMkIC2hg1GKXZtgyIbwEcRfhSgt8
dqlKLcfVZ8/Z1/eaDRZ4VLP8oF1mRIR4vVdg/PPF9RKvzOM1VOxfNgkvMFumScPr
G0WBhoJmlfTix14jyqYYWNCzNeUKS6HgeYnr9o38d10nkO4ympVcDDOSPLIUuBq5
pbhIhmdclArrLrXrOWKBXQnY8B+aHiTuF14nLBILIqWLr2pSNhCVdwC+AdVMQND/
mni391AoVWNMcL+cmaMuOwcbuOqMgIB4iY7C2H3EfFbyGP480btb1w8o69/EEA54
5ckXQUCgVGhfSuWqlDzkPFy8x8o7t52TUeb6PgwfJ3zMFQrPajIR+tAP6clVwsje
qfXRU5YLKuTFjhNc/b0/6G0kT0c0wv8m6wiY3b24HrcrjTh5RGnsFBYpfJVAcrX9
1sCB0IyjE8Hr6KZZ4ezqZqPC32PNDt+RqbXnldiHMKZzEhjCziXx+e5vIRQO08NN
Guv+3JBqd+MHDBBMOn3sT+bt0AbVsUa4XIuSce8CdDpDH0lIV6hhmx2s/ewl73E3
Wo12mMmxBeC6pz1+GlBanqHQHJQMIROCFtNSG6EVolMARGuE4qYrUJTb/n0nsLFq
LDnQhfTojKTVfyUmATOf3yiUnh1L67jiltg1jt4xHA5yZCdET7TmBFTvM5nZt4vm
Nj7UvaF3kWdVESq2rb79+RaYIGHlJAu4nOxUba460zpFTrcHmLxdek78QdbrP10u
LcZiLMQJJ1EXfUAA+gifniSW5JXmSdLGpjDLgmaxwmmtn81rJ/Gn2V0K+oCY+VDd
RjgUiOvVnpKziQaR/+v3j8Ndvq0u6xl/CoZbx6F9FIAFNAvrd5H6MyMNq1sBQ8VA
HgfY4Y3X91/COPNGPWI4DGW5Vcx75rM92Fz3/whGu3s2bncEEBTaDzqA3IHDyblH
lFMFqcLJ4dhmbBos+8ZP9AzSEYnj3VveegoWmSH8Vv20iE5z1c8zp55DO/bEXXoc
FL9IOtq9DcZ9bRuSro0Kogss+o6yRQEQJk+tWwoGQ/fZ01QVJzGuTWhPGtHwCDKi
wFgi/5FCu8LAGKWwB7NhO3mE5ZAK8Lo9Uk6bHdEqGk42BWsg8hVRadIi/pfFoafl
JoOAytxa8OVrLDHj7bnKeahhQYB2h09Sii4RGrURuvqrxZp1ytYcoDfsVOFMdW2n
B9RWJcFxZ5FAge7TFw7n4klcSstOCWkUGoQAgC35f5adVNnfflBesREV62SKFagh
AM/FI44sC7qZYGd4d4AT6zz0ao0TKxc6WEuqndw6w9Ddm6ya5OjwiQg4CqAvMT3y
FzPSZ9FhoQZm3sk12w1PUfJGRM6ZLKmWVu40D7/tOlKfIkmmBIIWYFyRk6v3GrZ5
o+RNF7EZen2+bgl04/vQjRpP3m/tuhbdDSJjvzy7HYC7kxFdmlCwcxPumYl8VtqR
FuM8EW8es/b8o+aqhAWnJuBtwh5/MHz+cXPvYyRLLmAIIQmKAjMOYYG1nD9rFapV
wgMNKFzGsoyQmdP8do69Hnf20/RGNWf2DLYVPQwH8V+H78IZ/CO9Xa1RxwjZwMwk
7qDjPPRwDObGXim8hf+m4/tIS74Vp0havkKCTqfAL8HQAdhHYXggTdiOERBzkjff
wUOmNs0QqvvAoxU9TlSpXBzKXkADRJf36zKK6iqtoXljYXQeGdh78bpWRPZnyleF
gsZ/2AiLW+hs7GlsCI589ZIqsm/GRYhbJ2kGlU7CWzxmaycu8s7nqKNawt4omSbB
C7c2sdhZ/0b70L3uRDG9+/yHI2QhbCfcxJ9HZKtbIF26t4XuS5Wt5Rp7d4772VT8
MIgieO/zfEt3quyQ93xR40Fc6euEzrAtsThqAXIS5rCHPCklnzw6y5Gq5eDCsfSx
NRrEI1QW6x7sX4WjK4pCr2LCgSSgtnXlbvhORm20mJxFuVvkbPOArwGCYJnBzF+n
7f5IUU22IGc59GFQvt6XDOvyNAtgb3rVWOVUsrOlMNzW7iW+J0LEBFvcYTaH/AhM
31KVMKWFUw50tBzhhYNApi26+rDNPVPqtEhtxp3rABXFpuZOGX5/m63H1MsAh8/y
NiAbcRr8FVm173w/7hye2/eDBsCOCzCnDaI0Zcw/cPC3pptFylrluAeKOvquPwnB
7jtMijd1WQvpe3CTBhP5yiAGPP9z+wN9rTkjYKvrIrpjdCdUW1IiGdNvIFbdqnV1
aIZB0uzMCh4Of2PnzpcalsAX/09yr9XVsDJ1BXa8011WPLH6szPyEmPwAE7iVTsn
KfrHG6HXixBpE/ecpOwDBCWs8KGj+5XLXfIPVcbkTaPsmjqMpn+Hps6eov7hvYIl
iG7UHSU7YPlAt4/o2nB6LndiFso0GV8yNqmNO46v8aUPA4wVQbzDgJdFAd7y8OD2
TS9gGHIeMoChLImzN0CIZz7lVzBBa+iCXzvVvoARh7vWnbSDrciN2lM7W04QuKgW
gkWS0jvdqSPEkK001o1jsml515oRd0A8IMjMhMCkb6TiSMxYCEKSoxcxPwswyhC5
u+4W7N4n6ixk3n4x64jMwbtWTk5meXRFG71ZxpO7IhGhWosvcTske+TcDHRY+CZz
cNtW9xszc1PWpVpfsUA3CJbFZ88guRzI7oMIvRsYQBm76R+8rCEKLiIe58+VZL6g
5DOJ017zRmDIA0QjqEW+ClEcxL2YfBRW3PQivMUXLUNWTHRBVrEU258pjMZVQ2yy
PDAdZyZ0BnRY2OzUCt0vEOz5cUEoNJVo4t9n7yE6e9IeoaBwWWEX5pgyIO9TysXk
dwKTaUVjapaDTMCuCudWgBXeavSvNdhEOowhvGeIqUYoi7TaFaq1xC6EQp2NqCRC
ykvzUMUT4Q4B8+NDEBsiL1zm8ij3MAsjbYW0LiBDo2uH7JKuhndxOL6mMoMQrx2h
dsJzSbSS2kv8ktgqbL2L9ZSXMtclkXfej0/OJCw3A/HRllewO4SZQmPxY5zuoHby
nd6oZw3pH8T5jbf3PfmC5dtq7wmGcaYr1ozpMOLTp82HPdvc1hMtDy8rr3xj42fB
gWj4k1KkehM5ar16gl8qyPVsOFcDWhSdnWLDmxSZSRhIXwXis8YUxx/tGdvbZNvi
8N8FkAg2yNVN6wbSkNvOeCgsSBrbxxza/NT0DKW/iUbNxF4AFRsi20Q00+jKE0JV
UKmBhE+M3BQ52r4vb9NvWPepz7KQNSiURNt5ie6TJdf56tYV18tWECDsw45EVK9S
mEGsYBz60+bTKFu8Pe3UD6yBGkRcAAibxc1KnJzd0H2a33wcF6jDQXmpZJ2YEq+U
HyyHnZrGXrXa3D0MXhrqDdaEsosSJdRyF/lHL6rSwpY7/7PDycE4uqYdpoAm6uL1
6xOO5oOwEbnjxFuJhMJ7ImPMznhJZacj1erQ3au4yr1R3qu7BVlYlj9a0NBTT2y5
Zf/WLO7bD/QFJ1r0D8ZPpV6SCbZlgrCMJwZMVfKMjrmfmQP8duEyVgjdBcImdLti
2WkAhVvznzGYvezyO9zjrsPKnhj9UADRArJKrHVRPV0DhtkIwxWm1NrZFH3JPVeL
rYIIMKA85QDcJd/TdJYzD+ih+UoXmhpsrRF76XbkmuC+KvhAp/AoJlC/8zcrTw53
/0so6mnI70uAQDd3fwwjYy4avKEdWGc0tkkx5OAmDNosN9aNRu5fb2H3yl8vVUqu
lRH0+IkitWa/wJ2jKel4H57/flcU/z9p61JXEMad+4er3cth4/tlToEZSSGric/Q
iDmhJvhqcrCj9JYRKd3f+InHi9Fg4w8cykUkPVu80P2jkE5G/GF+/SmrWCyL+nal
zl8B0JI4Sa6AFuWsyNZRWEoXWyUT/ufQ9F/eNHWE6xRgUOqP9ESc9QtFl0Lb1xl9
JT2VTKTWb/VSFN2liGmO7YcTO0eYUUqnGjAmqizvDhZIAccK2pNKlgdSCmfAjmYh
GBpjSs5gqlbdHgwo3hf2pQYzfOu1E8r6wTuQpBSex8z5uRtFpBaMJGZ/BasWoBkg
/L7/iB1B0xcGHZu0FZLUfCIlzud9HmlV+Yi9aPbGyD6J4VjSiInRFdPo33PfMHCR
WevM0zuuaB9DiUN/ZwjnEKep5ZeRvIWoERKWRnsdSNNHzgau2EaYD4NJgstMoboS
LRwnj6qEZYMzhtdOY4U/YiRENpIZeXL/Ab5lux0dpi4Ri2SlvU1XMlk1H4qBOiKe
Mib0oxj5qzFEeYogqVIsBypzqUk1erc2rAxqXBQa6D6c3JgdATpogh1i6rnr148K
4criQNFp3AF0EuIGvObDFjTy5g5rqjIIPNCSvG/cWq1mY9BKqY5ZCew/b7ULWavo
NFLdBkWSp/Eek7Az7en0p96x1F0OI75FzQTZcmgYHpHziWzOtvwEyOsKLq+TeXOA
GhQOFsNrBYFoyZ8kxEKMbOAiiKWvp8twQlHZUx4003PWb6z5BDp42WF/EoqUEOt/
yPe+ST3knHYRmgRRoJFg9Ky6p8G7OpoFpzjmz2Mg979Zp+aaihpyRAu3H9XKTVg7
BugnkrTICTbKFoKaPTi32HJFEFWudFhmXyHH0qAfqlIRtKARQoVnFdxe3cjyQqPh
f9/+fCI1tF7Ow/yjznEXDbVDabndnb988CGCgwtUwsIVf8n2kXaYpBOp7JSdL6kq
JvSypln4QdBW96KxiNcNCibHiJJ5U3ip9i9q4a0hdQzzqH6zHQrTMc05ZQ/PIUmv
/olUUZ7ABA/VjQtz/gUOqvFJDT3JzSzNP12oJCg3XdqwpSaLNWaRf8bWBmsRzVPq
T7RDALvSJmBSbf4/jgmGI0KMTcnOVpXHSY4TPgv3a7RxAbVmw0E9HQtAsRbrII41
Ip8zsQ/E0k5tcRR6qlprBQTQqdE3XoxRrTnsZaBqsz+PltON159mb6uGUTiR1CZW
D073zO1mN6SeZHJXspktRAHwmaZC4KvS7pdnO/VzxNfOWQ4lyaM/FdG3IrF2j7ab
f9OGjk26EZApARvhzJfJ/eIZVMEoWXpmvGKdt8T0IfIKkXdUr6f4kgHlzk7pYqCd
j3JbMpEDOK3Q1UBifaoUuYPw14Po7vYmB3EU9Qcs/TK82BGqeaclQPql1WmyeyJi
NYY1jQ1L0mXMI1epyXTDa9eZvuFenD8ywKlm82nxJnEXyNF0GsoMQOfyM6+mjt33
/bMA35J0dKucvHZOQzpY5D69epwxoExG3NkR2KrsDzKMC07kwmAVzOY0MIS9xEZz
FWB6Pq9mVjDz07Zgpwh3YlS2PP7TkQ99f2wYfcH+PIhMzEoF9qsQUfT3sH28PH9p
4Ugsjk5qzfR4JTuHWDHqmRfBXMXS6rtbh4iwUkI69ZJGnXlznNrs1qsttz9oWg4D
a28K69sAulQ6k77WgsEZ82nL17XfOkyg35zWE/rUbWmHpgYS5K8gq6pKyEu8SNMV
2jK5HXzwYyeCuGnfBT8DLdgZDvLhulUX3E55QfLbQ0AvFQS6ogfPpCs/gbaSpyI8
DGi6fxr+AO49oGnyAOYIuGdbgwKdrNBgE1U0LtSXbS9UjS5bjvEMc5C+oBQk4mNy
Flmklr3H+xAuvXTquPd/g5MMNTzKHIJWuF4ya4QieB1K+aw6zBpOj6tYf43k3zS7
kFC5/O/J5RpZXNNXGL4ibgHnLWXFVzmJbSU5dT4wswU5bGvdn0jwjmfT9ZTJUmES
ZD3vV+W35Hj2waqSh/teEIQaDPyw4zG1I2LVGkWhu/dNLHTAU5gVZTxSxMFQj3oL
vzu7DntlIKblg1O/oYrMWAhaSquOjtGNBIdToOO3bDSkmz7IBF7IbU/QCx6JrU7p
jm7L8cvnlQWjme5QC9IINUTPG+ZU0ANM5EPR3Z6MArIASyAGpp3Yf72IThj1YXnD
Di9ad5oREg2oG78HPa/I1d76AcK85dlKygygH/s63ea8naiGpX3wKY04mDalVx84
m8HIjV15X4X/+72WpuIlM9pQ0kcxiLXnPCsKsNe4kd7mTs4fvo625pykjs1veVpk
RrgHKhpexQx1q4B8xcmgvNcu95wqhxH67+haOTKVAEPhKMv6wopT/DBe00WmpEgV
oAb4TvMHNmqD/A135uRygI36lYSIjjymNkvncgxUlZYRGlCTbqi5e3W5NLNuJTfK
9g2qvOYV3Kz5tjcQ5C/5CSAKvwJ4N+D9QX7kQOlw3Df1UMJT4iI8BRRvkF77L+/1
1y+mxmD7x3+SdmStnXHCBh0yiJqJD76NcKrZMANdTzE9IZS+M7Hwgi2OKyRDKV2d
9+A+WrAvUj+7dLXV02whh0WvMgqtHZrkWziTMMn5ZwYtuIv6alMvca9s3MARjNbF
z32EIFwmqif1JVPpmdjEbxe9zk3NOQfXbJItIJn3x2D/LyCWFZeGvw9AB4CCaE/+
aNNTEMxjaQ22/rQLH0mDoFUK8u5txLZCh5Edzl/+2JVU7X3qJtJ6RGFryrEFZxyg
PL1oBC/Qa020Q2LzaPH4vFhwuiDrFjwA9Tv+jA6cGH9TsVkGaPSZ5bN2hJZaD8XC
11Cw81yrmJZ1DHuFcC3nuT88ObLHQ9bT0mIZkSbwDNVNJdHUVt4ROodfUR4OtsqJ
+HjS4NzTbsu5O7DWyZHaO6ljM/4Z56oLVfe7igx05AuoLxOQkCoFsGdTkgYsRBcO
cahOAAu7TJGMKbQOwMF8xw+AseV+6jAmrJp7A2R/oOQkXoL6GGATs8PkkktclMUx
ho2tSF0ewA9TTylj8S029gvpnn+vyCY5H/60ENMS7ikZ7r9WjiF2IBy2hFle8tqN
1EsO/iumwHJHxqZWYHzRhPtDOzmL3L8FcaRFDWiKnCXdx+M2MOpmIs3SSR3JlYLj
m8wzswudgoVk6I+4FkJipF9EjampZmILCfrcgr1XLyyHXZ+gcv79q8OpjYwoBYlT
dPvjME2bF+01ycOY4AMcS80jE+4kKVYVu/VaVH9cJuNLKIRt5e0VDy7llS6SyXIb
P/3Z5t0gB59DW6xX+Gj5hMOaHF6zbOLvtWUccclHHC9CcLZAVCHlfwmgaAGQcIyu
iIyj8k4wyOJ75ack+gc47d6h/TBubAUXhqO0lyB1nGk5qvJvDZ1PjuTpO864uJ++
eb33VqI2R7Ce5FLJ1G+tZXDU4nxCut1FFawTB9o/XgQG/ru2Lbb2EBnoDtIQZVty
QmjjCs2AL4MaQuGAb/eD52K27MdVnV44+A2M8MRSbaQI7a05CTdU+Demeoc+yw8m
iUVm/K0Hka2Kf9zqFFh8Vb8LGSTmno6XcQ3XtoSiSv7UeoPNvXDYxODMjXm+xZeq
e4yPP7IH5NgUiIWMm2gD3IwXEMgC6er9uq5swGAMEfGkKVD/h/4WjWbl1GA9j8jz
TkyN1TMbD5iboM8JkjBVCoUNwaKFz6wE31kJHRLzX8gKszaTnTIrAd+t96bO364A
mQqSOobBoZYDkvVs7n691owjg5/uK0uVqUvCBzk0vAFqJ833pJW5MmM32TGKsDNw
einmsX8Ql4DKvAKyTvVQ0lcMsMVTQIJQute0ZvHi5ptZGpLrQvBaL5KBYWXiHOEQ
NvgFwlnxZtHsh4RkVg2BHpAzHbgfy4XK7lybonlE8mZ8kA9KPZuejs5NEY45etOy
ZLd/4Q5ddwTVoLzqchWUzyrg/cVVWSgsgTh6NHzrIr4pUXYswkboPUtcXr7wIB1c
4jsNbr7QpwGvixHn+9FHSNeaYM+Fq3m8YlXBNBjILlo920xTcfkpKqhs9lSpC6HP
M0/G3SWEvIWt6bx+Pv3aEFc6fY/Rmggw3oiteEywgMtDykYOs0b7Nsg6YZGIUEbl
XXGYUV1+L9OK9ADidAB32myRjNZNx/yWyhh4V7pkUx9tx3C406Gc/g1D4JT8w314
mqPxexCbzNVu3pw6eQM4Gzj/p43oDSgfzppViUfmp0P8ZisYTfG1VbnflbE1Bsfa
CVXiMOYuXkRke+z6HybCuBN7u+qLxJZoLKpxzjBoq2ZfUaZsIJq17t04q4XughGC
zrDwX+pcrJO+mqsef52sKN8LYWywF+AEaSeVaxuLHTfXMjtdxIJvtN/Nv5w/s1JY
arPua9hMZIJSMGjLTvqm41vlL2rXwyPglPOT8w+SvUvkLjUMqfLF3rDhHvzknqLe
IC1WZRG0X4BmFa/mfc4RU9zUxj5uaceOeCK7EfYe4+kTnv26waZbRijLbtt5IQJk
07DPFX5y7XH+fzMvvG/W0nJ4Mt4QLKjaqKhUSDgydnYIgkdZJRhLghTyKOa3jPaf
M9dVSsy4PTVqOLgtRNQkZsAJyoTgLoChCa8iejlhfCOL0Wh3kbDpif3mN55FwSFQ
wJO8HE4/xGj98CdxlUuHDswMC+5pIsq8Ebyc+95UQfYlrRI8lbdvaenzeR3F0dss
/xXT51c6bmMJ+MHCfFEoiWURXCx9GiV102KpYI5b3PFT2roZy/oL3RM9JwlqQBuT
dDG6q/1CFFKw4JuHlu1zHAZZf1OAiQNyug2vouSEEC/bsMoiAfJyAWWj+0QXomxk
yuimhFUpcdWiC4LFhfJu4+v1IHuynw2n9/stgphggCQ72Ae/UfqJWlbFGV7Swu2n
p9pIFV9pZq2+SA5pnGaJ+LdIYfpVP1yzfGvppKE9lLmou/V/L9XA3xnuIDU4g5BQ
GkZdFqC6MK4YmbpxvQD/sL/4eXUYc3F4Tlkinh3Xr1Aiu6pdNVNDzwj90Jn1H/3B
T7OQWllSRXDY4jG9XdctvMdy9pSckMWbrrBI8hvX2j+GD02M47i+yIzWD475n52b
3uAfZ/F22koOMemZIBjtqK2Fjo4tlLYAnHTJuXpOI1deyv15+qr+qmWV7ZnmYWDL
6TdtsVHGNqx/tIkGelRkxkntVimeUUSupm0CSUS8SYBari0RA8OJkEsz9I/Qqk1N
vTi2yx+EGpBIKKKCRvEX5cVgmeaq/g8apL4T9rCqjyV28wZ9pKG4Ab+UyrhIUUwD
8L1yDm3lSoqy8nyvoL0m6V2v7woHFhgpA990WK5AyjlDyVtq26IWk9f9MRexvmTs
T547qVzM7zU9BjpcKv1I1iko7ZSpFEwrsDv4TOmDNXXZdCM1Ppw+Yb65kvzUMjY+
TZk6Fo9/IVP1Bn+G6AJpp6p6NABGRZsXVJIhEAUzIcHP6xSaBkEKjthXLHC4V39t
FWprW1ksLTWtXnpEwyZAuOv1rI9sfPOwxyDhzBfEMFbWuPHI5vcRZLhcRaB1MKgH
5IC8vFf6P/5WNTrANwGkQfpaLGLCFnyoTJlHWGkPkH7JqdzrRKR6dEFQeET9YdVv
sm377h61J3QBOQQiPMfLNu7TydfE7YXNLP3AsF72V9MyNNII2+0H5c1rutTusg99
2PHXfw9WP1aNzkjXHJWD3tiwVYB9y08A+q1h1ptx3EC+DzGuYj3WLVWSLbx0Idgr
h7WIJ1+oxYVzCbUqM5TvTmtNT1GAa6F3VlAadKFKc9xQt+o04VXwPJXT5RnvYap6
jOi0+fS+17kyz8bGussHO2wZrSdMQookdivBHKTPc0UOw55xDuN7bqtQ1X6k0qHi
uNArwa690v0fzfh6lnb31lzALiWJGrnh0zlvDOY6e+MJLBN89rgoOs+qMXNqddHM
ujp/s6OBGAWq14OGDsiewu7vkg5lzC1Xe7nFuVJENbXiAjUjyMz91DkTVobztNGG
5SncVpcnGVFA1yNJUXpzKF229+LmneIP0ZdLW6gsfS4K/OFbuUP2BDJZvup9BBLb
/W+DFNfq5r0nmtCCSc93ncx4PVcUy9jr7cipDRm9DhcK1ObBpcVLOpJZWy1cFw5H
2lrv+VyjEtGBWqjBgkFp2CXMSPY4PUmNBegy5uN82PTYQLlNUm4TwTipMv/sZ8OV
uBydoj6mdJd4UrTBQAN29Lvg+FFkBSTPDFQQceKHbjfAcdkaYDsADcej4BY+FkUF
p2qdDzgZhb9nG6wGUYhySBoEUkUBNTPMPslOdQh99HGY89oUqucyYeoulwuEwww5
9uPk/HpaJZLc5UevBgxaUdFxTGS+uv4ORJCRgvX2sKHdpzfItDbJSqUcp/LEfSMd
kEkUYQ9eg7MqhIULSdckZYPd6y6rakop5kLhkisSa4PWUenZZIgB66cxMAA3pyJm
H5YBZGUjTcIqahHF2ijW6VFfBfQKfDAENQWDNaYj4v6x2HQDTGsYfCIg712hURml
0t8n4SPqim0gP+EEN44x5SQxULo+axMO4iMHCCVy89YYw8tRo7CvQqqsJ+cq8xBj
M4fG/lG+16Bs23JVcrLY3Pv44wW9BOXI2DetPf1z/w3dHUYciMnsRuBg5d49OJvm
ryZp032SoZWnUlbGVUYglUQVTMQ+Gy30eSFw1Ezoh3qIaAYLzYIWJ2gC0naihtWd
2IxeX3651Q8D3c8ghc/bqWVUQ1vfM+GN14AR98TlJodGHN5pakY8gKbixRNlGbu0
YMkBrTz+iLs9ywK0nT2ADRLAPSVtFRaP86XNMrVjG1k7zYOCTESiLyow49Jd+CKO
LnaatSS2Ub3ujWdpOF5SmT5NwBRHQMOG2uFjyeM4On3ukFBdxJy4DKRh7461jcZX
YefU3ynVXQEdGi19T6/yvWJ0NS1AAIQ6ymwhEkQBDsNKfzlFbDex/Mv6WIEqH0tt
X7x3Yr4OEW2TRHZ3LareVhYU5yvQmgvt5QxsOjUDCw1SYkSF6ttQ2SaLe3WxYvSI
qltPHaCDqqjzxca9thAmCxPv+oUefwcdzcQVUnAAGFQUpYCGwHFE8i6ZfpbhpL1b
9i0Uf4ijgaO0HkjKEj+nXoX33mCATMnoToAHSlHZH0YQqgN37NSkPFWlK6RCnqBY
xiZyiwk302o7obtPvRoHcVY6QjAUOS4fH1D3Xs/y34qWzTXp5kPe4YUwZM/dOvfz
rJwAMeVkXGjO21T/GuK2Or6p1wPoEcLD1P9p2H2j60wex3tiGnt8EvtuBOQt93rb
uyBVQBOUPJ+eH9Iy+e1XdvdFicViIt9NJa4RTfIQOq5xd2ruTACx09fwj3tE5tpO
AjVbudhXy7ESmQZz9N632dqUFDBbBzn/nVAmroj8ikZ94HzvrUj5Q/pFJse9PyhI
w/UXQEQir3Nt2m0xZnFrpq+QxbGsITd/hDauMG8djvZz7PPSGCABuPF1EPh6j2tv
ToZj628RqFAtOoDyOxGBqpEbqq0Si5Tx20QbV5ptzVQFGjJbOUqUeMaHhLTmiG6R
o6aMbefbXTWWyiOUsKKBKjVlz+0Bd04hOHOfK9DfnrpQji6h/TPOHhlpoGY4uM87
UI7hiEJ7PVHYYPkVW+ED6rPNoUKEpxgdVXm6M7Ol7BnuJbrw+WHRjPkNPD4c/QP2
xtge3339kyWgwr6Pwvqu47KyuNjQGGuR50KB8X8OWFURTVfXWbqG9QvYiGu9MjpR
ldrf4lfilOIRXfLsH2CH+zEwpsXRm6nDzc25IgMbhRhLKCIZgCmffRzM5TBIhCXb
2nkE25aktENZjnpDBEtgvrfox5g/KyoRwZGSAUi7AcOM+O7h6Socu/vbnruR8WPb
fLUqJ3IXFd1vvAgv6KInhezEn2zFj8qCsHgZkx4jQDrvdDVkpRM4jWCoYM7MJ2t/
fAMVRrHsl7YgQel5rqnqVyI/EB/EbgQ98kMAYa2k9Tp0lKOu0P620Zyb1pqwJiOn
01i0yIlN2oQ2TG23344XIOkURLsmAcKnVn7RQt12CHMvBK7Qqfglbz+FYAzT98RU
oJMARdl35TecnKPicrfk2wS1mTlnUzaQAja75gphqVgcoZ6l2zEQ9hp2YgYjFnmk
QvWSB3dA/ozVpmnOgzWwVYeFZ/iDUbgJAxTTfJmfQprbVkrE0ozp1+O4MpQWQfVA
0ZpESC1Hh30jSpaAGWp4DpIfzMwIoHA8AG5DshxQghBDMSf6BVV0lTHM266j5aoD
7Pcr1edrhoaRMWoHztn//T4WuD48pPV0LBxU6oRzbuFrsASupcidBRry/a8IkHVU
XhPNXcqbRL0ESbyk4wqi1yuKhlDRFahpSHgINbGeViY7YYlcDS6e9Oj0RKxKEvQH
jtWSifVxIzZfNbGtNkjZW1Le+GOst0GZRx0RgsU5HygGmEYZtZFTtrvmQ+fy8sgn
tpQH4CoSaEhWiAalDW2nzWp3jge534X3Cg9AfXHONDDXCsOZKEIOTbEh/RIqSsk9
18BL6CHIoeJNjTBfbGIEtHyckybShGnku9ml9bZk22/W5rx7P+k9mVRqN5LzzgU3
r79yCIg438mv1ZvY1qYqKDb+BVE/Y7spsQoaea8Y5dY2TDKT7+3CsM5gccORneTC
AyL5YeK1qXABbntQvhYK7kaIw1vlJLgOv9Kl232TgP272bT32BMBlDpux7JEegSJ
Qh/rQc8PJKSIZR3N3K/dEqxPOlQ7SByDdviU3wdMaeoFe3L4QNkm1H2ctosoyuTI
vAbM3E7o84FidlSCvpp6MfBrlyL+NvZldd0jK67HXWMBUOYrQ+Mg1cqSxC/ioISt
oE1fN6HQyv53fXwtPRyjlLdsKcbdMHeYK6blYUPB+37qb9oii6QAzFUxAfhMQrkh
tXTZkMdwjHq63sCH2vvtp955vsp5YOo4kdboHtBHqm2R2ZdtmIrdwfZj0EsAEiGo
JuflsqCXTb8KQIhX5ulCHY5olHhk8hcM0XWu3LEXRH18ZcJQwsxdpF0EuGsTnfEq
/81t5SDKUo1j0xdDhIFVsKAf+wxkDe3qp6i1hGwMdeMoOc1yPLMqgIApz1sxRunC
TZzqIhQedyspksu8Y34+v8mXv6RnB4Qjh6H9kNGqaYbyLcFyzLWxd1MicgRUAVyS
iLyKkLCzXBubK4D9FyUmkc7jixb4dwOeJzTZOPdINb3we+ICUJyjwIsdbWutZ+hr
5tWgnCDNQt/v68tAy/VVMa1pAdS3BgMcq4PgXVAn9SYxywrJ0IxORjl0QdrAywRo
qOwugO2n1rbRLaRgCsolphBhmXZ17buN5qFsZWwp852X2AFQ16IS8jMefOn9kltJ
kEQ8kHUPgdWuzOI7OEz71zwJyZUpfxQXKN0/PWKJwyJDsceMwprZuUhz7y0JevfP
n6xS268kxwwKIDO2G/e4HSYLThOhTIQ/nS09/UozTpHc70WQmAyPRMjgNhuNSJmm
fb7+iQVue5XKrCVf8Yjz3ZQptZYqr5rxhtNe7PGdBQ2/Ne9T2pcFvQejr+oOag3N
d8qwmrGXoDf6dphXjidX8TFlvUErgakmZJh6IcTDtwY6v76x+9Np4VUhTv8lf6fk
SqLi7F6OS/aXuiKRwnxCpQe+YSNCejtXn+/nsQx7OV6SFtelPrhSQhP6eDA4lmRR
Or8t9B5vj429CUJDWy+mt03Af5wd8l/TEjgij2ialJ3ZzJMh1adVoihM5TeKUlvD
F6eFTiY74b9bnT9SoIiuVVJQJ/FhUBLR2+ggaycT266gTYtzxRU1WyA3Kmzf1yMj
RJsb5MeGUfp9FZEOhzS13QEbTnVS06uz5nB/dDWH6SkuvfV8vxhlRoUYUsKtQ54Q
D1WjD+JucDbqwPi5M2VXC6VCX+8Vep4G5JcEb7jKm9jxUeUmpij/fJk8aGgLhMbM
w2TDJ3dch81I34x1kDJuThM5kaJX7IRVm1xZOhC0u2L5zOD3HEqlOmjLxblydy8W
r7XBaXQCeEguD54vGQdX4dPj83xRqnPMYQUkRnAAirNc4A94gtc4yy5fGwlKv3fd
AP25+j15ayMeiDC4y9dEE95aqxTh2bOSEM4RyouTXqWXJxk3tUzrYRr9dcmr8v9f
iG2t7mXdlRvlYEcT8s5iER4MqwWbGNMbWTDhbOW706i9ztrG6i8nwZRHrJWvJXRA
f31MTxO1svtrpyxAUykBHEQCsNIPoIAn93LVSoGuZWeoIVA4XNS9Id4ita6cpcal
Rvb1lP7RRpPI7A0YOII55R1mRjxz8VAfIrcOmkeatXFLLsCJZimkfilXbEoQnVc2
YXm+e0nbBqtJKQJZhGzdsNz1AVfrTQCdrl1F4llfJGhMncKm2fosjUb+77ua2EZh
n9YVZpcuDRkdG1sTuhN60EYqOyoFXLsiiXO7/RORpj0WcJd9XUVAohJe7uiebiZg
SB2BB7/Yc8YU6cn8qFD6MWEu6VVOd7E5cmh4Swp8BQa2NFg67eohkLCk/XPkl1SS
2vn3eiJxYbNn5n4SxLQ8fhOHsWYRbjRal0Fksod24CblZX/XYumMZfqR6Fp2L5Rx
kBeGeU2aPnJGicnIXRBlxoaC+aGcoCd4vy6qH2S6xn6wojYQwnDltYK6If5rAtzW
Y8yKdE1Vwq8DxYHZsPWArujxdFuUDimLg0xpPF5G9X6dD6N8nYe0UltA4KxEXgba
LLituMPj8XuvSjg5udiOxDrsGtQ1hnvaNKURelKqBsceNgklIZ85BOeQApbqD3dT
7lNLeR/H/g3PL3/mqrDg7tO8X3Hu+hQxGdTBSDBfScjdPoIBk+6w6p5HciUd5DAH
+PvQcmX6eKPu1f+9MKaWU6DhZz/ooNl/ype1EG1NhQhRuahF4j2pzZSn2EBNeDVx
JEvDR/uWtsqJJhiIfL3BxtzSfQ6370S/U/w1ZjTghKfYnqrHxUVnM8lXI3Y3nRWQ
3TEzcWeeFxh6Cn8EJK+aqrPfOsVBK/LQMK65W6ZoSfDaXai4PXWA0zi4T5b6HgP9
eiAqk8lSQcnWXNyB9HL2BsP/oa7Nrxm0wfWcUa6ogMFnBPSM9Yz48kJea29THbt6
bqWwUvH7+WidG1PmojTyOE1UGobv4AelggH+3EH6vBvKLJzcP/IJ7UO9JNEirO3P
LR5jufu1KSriLqU2dskaRnU3eiBpDnANtrEQgwBl9J9i32mxZvS5KApav5BnZweo
+2CVew3eiEopbL/XTW1PDb+SrW1tJal6Px3KOztJij90cSmbxBs5qQNgSXBek7NG
DGoJVftmd4e3MZKSjhmLtOcBJZybBWEPmtzU/kcN5ZRYHR1AAqOs51kh5/HfHnpP
WfZ2cAGZvIYD5+tlTlf6eUTAdVr4I58Tm2Mtd2Sbfe2pX2gGexHR3sZtNZgu3PVX
gDEOEdt1sDZCJ7SssSpbTzcRsF5lKWAIULUNPs2m4LVNvIQXWVkzdlppUh09mnUm
n96U102CsdJ2QaB87f4O8TmqzBX/P2WasCi26V/NLGoC4nS9ZzhPp8iYG69Id1mK
TPfpIn7FBqsbad6p5r5uoRCdEYK8VFt8ryNvAoZ5FESwASwjsqnIv7a6wToxaqg4
4n7TsxTkVHwVt1pGvw7FBii+AwHDlGCTf9Z9UfcUY64kYMyVZEnl2jy/eFmjGec/
GgjGxEVR17TGCgIJ+34FD1tbX7YaCBYEM4xtyvwLyeni3U8XAxu1kgPq+Xivbv8i
WNCs0zHxJ8ASNyH7lozbPsE+jmgoUsNFobaY7161M769wokQg0++I0v5V1Ywt7Uj
A/6za/NUpbnzPTdI5OZddROrkPiJsQIBboC0v7HTlk4UU1bLkKP6mNDRVURs2r/N
8vscxrzdeJFiU+i/12vVVeX9HBrZPaQh3fHlofmkzjfpF9ex7qsOQ33POeaK9Etf
GidFEi2cn//dV454f/Jar+ixzFpSllW73dZklaIDy+GSQpAQAo1NrhEXKKlf1XAr
72j+SPMeVFAIIwojnJinG87p1oVZliv6Q2zd018Hv2dR6Gu0QWx1qONCfvWX2tiy
7Nu0A+f1MSU1vfWvrov3Fjby+AcKmPSTJ6e+QkWUgf5u9CdScA7PCniPqeHbr0+E
IsGESEeDOSbTuDp4iyT1Lw4gi41P5pyGqom5N5ccf5M0K2qvW/Q3v1sg7EeHXOJi
KM/BwPB62XAwqjUzI7wrMPVWWws3Ouphi5GSMv3o3jWUzrrpdU/znJiRk11SmIca
sk9JqbQzq+hNGunN3B4RY8tPoeL66hd2guhUn1ylzUugS/hmQHgI0pUYkcz6kbnG
BSc1BqNATabPmRrh3CgXBLc2Zg76JUj9eJO7cPP2S875rvQukdjOpMNshDP6vq1G
c84KsUlCVTHoloPs83H3QV3QGdRGM/4B/oUYeeOyEB4FlPC4dw19jh7WFV7/JsIz
Z6kkglVMda6yJ90z9lBe5PqmMjuOTZbiDv9FMlEC+O8X0qV1T6I1qy13PaEcaJfx
4cWBjjbeOamo+FF/wTa6fGfJgTqwD46p3SVLvjGhkdcn24dxzA/eJfTaqkHggjJX
uWxVm4xuCQDPZLbp0Wqjp9g+5sq8ilQMYSPlM/6WXVaPLXRI+q5I+bYg8rqAEHwT
TRWnREYWSgECV86OVmqt4wXY5u7wad0XyzwdNtnBWYRZN2iDRbMwCK3QcVh3KPaf
ESgCTEtAJOO5xb4VqBg78IGH0YwTqwY7INxngcOv0EUTlYLJ6M0XsiPPBorfRWxH
WjR8556Zq7Sh1W4e53KWcCA4ZnvOe1nlysc+sESQGRloPQxcriOLNT/xCD9+eeSZ
iSpflKJKmrSBV36pzLAwcBKP5kSzTKB+KlHMkn1JW87/scOuJWb/8+Tv4DjwzufY
EWV3nEk9hu3ReeWeeJ40j0yCdmujPLOXDOX/7Uh530iIUHh4wTMUlc7OMPh8H5vE
hab2gTWnQj4TWLo92FhRmDxKhk9PXuomx6nTNDCajmIq0DVNggeWsO42JosXF2HV
5Nhj5ds3+eFYgU5nPhRICv9GQ1oJJR4BfzSC3i8Td7PEPO/rWFjOUXhkoGsJqExK
u1wAjaP7G+GuYEv2eG2hqMZkHLnRzW7U4pT0m3m4tLu+CJ4qlVvmO7ZXd3lOV4+S
29MyVon24Gi4SCJXkf8boqp53ha3bJdu6xeB1Rz/4gGiI4IwanMSmED+YlG9FmNe
1tTikIJdStr5fFd2Qlfx8YypPkslilWmfuPH+n3LHJ7uzxcIq2OZW5b7QS7Y0lLK
7YsP+c0O5oKrgwiyIu/j4WAasanYwdDqzoOHMzdq8LXYlejCbf1Wf9EvU0RMYNu8
x9y7IMDHtZGF60le1lfktksSEFrYunIi8QVgxjSaTBjL3Ty8ceNN3fPNuFXEnM09
3FXUxhQcOwtNmlhdAiZ57+kpnRk8D1ieDIKXLxIZQo1AnyHUPjKxRAw7FYqOZY+3
AwO76piyL2yf07F5iBrvmB1Pn16rrAXZMyDn3LXlQ7zkD7K6OPjxQnD4M2+whUlJ
I+RAGgyjD0gvsNk4o1m8Si98gOZP0EhuzgN4yPRuNsXtTEiMUCTCwWz00Vo10kIA
hdwCjbgGOZpy1mjK/wRf7IQKdh8P1cTlBOwqbMD/xPNZRzz8nig58s1OchKGr7St
ZWpilmYFc1yGAnJKsFXVRmCKYJepLItHhsTiBFa3Enr5X3H6IhSNJqoA/RmZ9HAo
WGA+8CkxEF9ACBrZmTGiPkANm7o+sJqBeJO2aCH0KgAQPM9wsXflHPKIjkgFwq8L
5f0Lou8KpPMVGfvud11jClL0p+aBt14ws0qdxaTtXg43yylTUxCwAxCnpWjJHiRm
vYfeNidGP5y3nhcEsyFvWavvc87jSg8rOntUG02xa0J+2YSWUscriE67wym93DnN
/ohQi2jgkc7z3JCM6dxfYjIlhakpExSXV5Dk9R5y6PWIN6nXblJr9BcTIGoTYefS
CSjoRcJ+CP/elCILWltfX5g4G2YR7DYld7pVlyDPgJ8Con3ABFreU2DFFql7WpEl
R+aMUWOGc29wpc3gKdVbys2PodqZ7r4EjJtp4iWjquoVi1wyxpSiM8xlQ7CRLZjI
HjRW3SAbD/vMTulWCMsLcElJgAQzTU6uZjR1ZtkQOypRJhYWDTdt3z9tBDeabj4j
bir+NzvxI15624qIoxHw531wJOFpeefPQfLU2rO2U7s9snkLsW7o+w7vn8SnB1/T
HHeqZK2/Rg9KdyiJCn84hGBcI1tUUOkkB6vjwH1OsIQXtNMekOdRhG/4EV+6p6DB
cTGw0BVPA65RohyIulG4s8M2q6mvhd0PlJI6D4WMNFuQbCPbhHC0Rb5zKK8RFHcK
+gc84NMCBYjqVTmZO77esxr9bY58UgjvFP8MOuO6Uqo8VHLZ/tjPG2cXItQg4xcu
DYHMiDNk1QQ2qD8jyiZCpXmS/34qvHoQM9xcT7CkDiZEgHFzKS7V2OKlNCT3svLO
67HXm5weV+s3LPptbCcFdODQMTbiR4/H0mHGSA3z4EmiCJ553Hn10WfuEiMnHtCg
oYBIEeoWg9/fKqmne+X/BD0DjKH0QqqRvvBG6e81QCqi7pdfPOgi48j+d308YBLv
KnmYyukrYYUv8o8+1xWn/w3tMWUKf4KG+edOeu5LUMgrZyC9/MzmbeBW5ZAlu09z
rIIpS0uNw57E7rP71nOGOSPi0TASggQK6uP+XF0XBP4jsaangTlushEkzgSzyY46
n5aIKeCbb68RVXlvCjBAEMePLx8KXtYOEu6cWuJR2XsPQKD1asUEl6LtdD8iKKfl
iqh7lVyiswHnlxoN5j5sSprWEJbS+ViUymv7ejBTqRUPgS7MfCa3ajHtx2b6rzT7
mFCTDqt/WpsoOxHHfowMaHasDIlF9oG3QuKYM6/EhpqDvB3GoUDg8gmeD/kzdf7a
7Mq0ZepwHb3a3Muvv/QNHNN3Z88ofoFmh4BZzisUGvGgPtmCWfimxs30anPB3Wzd
52/mnKoOc3gjodW9vtAJqr7jGCeiy0tA+BjXPL0qMxx7057iO38QPKxZLb/VUBEY
gtlxBjZzASwU7ocSOyvoSxQWWRtba6Dk9/hLdSO8B2IhYc49cpXIQ8491F4D/CbO
YuGFBqis7lvjeerJYXg1tLwyKqln6xL5ab10tv7h7ol4cz00mTEI2FdHnhchs7Uf
zp+3QUf0c0+L5uaCWZHxz9sGJBusy+PzY9i7LJLikoT6S7Dzt/VQPVA6aIOV4JsZ
Q0i1q5mfiiJi1/vy5QTkZ9LnWDYWk1gGaFlvOi4H/aoaF0pvh16aqfVyv0OkaJkJ
5CIT58o4gP6U1Nm4OmseqXHW0A2wTdM12jvz+PTtZcMgKfXQKl5llnA4p05aHpFk
yM7CcwcFdAUKKIcOKGr34VZXff+Hqk0sB1sksN6PGpH1PD4Z1WwKRxIIGFtCru5l
wlYeMHuXE2Hbdm1fx6Y4cCDfPDOr7ErpRH0dEugHc+hZNjEE6O3OvhFtfnP79cjn
j8tTrDEvcTMW+Ceq+iVhsdsDYTdndjNL0KmZmqnzMBN6mWApA9nBqw6FqeZOqJp1
A5Bq9QicV/eLN8B5C6FOTjKtvdBd7dA/otBwI0n0I5XCzbabI7yxK3ljZYIPGRvV
Vu4LsNu965mcyZ8UYHAaPW19B7uusVwlp3P2qLNEPNWY5WPPqdDiACLXZgyWp5MJ
Lk3Qw5bAqS1r74uPaWIlamIHkYPXyiX1XdYk9eRVZvnLdPSU0OBFd1luhMHaWoUo
CyDVZlPh9+r2ADrVo3WHy+oClJS5BHq9X/qV8HruRB4AHWpo/Mq4h+DS3dLv2YXb
UuIuNmY8PzjXolAp8kS6/SzcrbUmjf07AzA/iKnpJinOzHfbfofW5MEEYXN2qABT
9azZ4eDygpWakm59ESsxmX7brVMrneK2/4aSeXL99D/cbVbEXOrp8qB06WQ2CPEy
6I+NLK7Gx1z85c9vlxo+HCw5W9xssj+FHPUeAhFL4Tq6lf5mZKebpP5GSk5vFBDL
kyaaLzjAWCacsd3UWvjNdP3V7Q1wf2xFggOZgPptiNrGCWfMl/daBKQ2h86Mk58G
Y5pw78l9ds9mSmunkpSe2rDd+vRQgbuPuDkavQAPc0mB7huWuLAGqA09Gi9OQXFB
rMdwNYBqzVN8ISpe9sRgN1htIiwmhdJbmr72HrRT5NCaFZeo+e1+ujSbiBO13AbS
78RV6shuC+hFbYF0UQta4zn10yGP/oUv5N5a5OxBHJfZ9vgXiUHycV23hTqMOsOS
STBFbW0w0NVur6fmfbSRqnBG+AmfdQZ0Q45UwHhnXlOfly91szGeB+hdyt15sXaU
G3mAmTksKCDvI11gWCuTxo1PkWWWutSu0HhjyeAxhXibvlStaWeysKj5EIuubiHe
cYRNVxaPtkiQkwFoZL3YitZlOjmUWeNtn02AnXvyq4j1ne4tIz/R3kdBj2z8mu1T
gl+mO0MCV3AU8ZiyL1Wr7WAQgxoRBqaosCbv+wTgr2P+LlLPgAgkyF/adquHEMu1
KrzMUQYFATWCo/eFPK96m2Kv5tbOx1CYgYbHu4+6HTCc7YMjaEy5E3TXsMqfIXbX
wA2JNqF2LOVHdkp8RHqOuYPjTDe/LIetIMyMFFKuL1fe+5mr6Mennkus5C+XZfb2
sTgesdpfx1u9W+ovjP6sBtCmq7DVpbhLzzUDu8bs5EL9S/rv6HUc3+mSlGb1/trz
QM8pEM4gDUzH/V+JaVSaThevzSd0Zc+9xqdvW5UNqRuSBVnFbRltWORev/Dax6NA
JPzAC26BOU/f/Kz4qr568qArkS6OjNQdPmKDOfpnbyoMWn2Q1ZDR8xKpabyje9CU
L53CYW1j2zM2WUl/lVxnX+QFUzRjE+rg+hjeQmxFfYfsC12NFKkBdo8ZNo4gOcRg
afZvv9rsddvcqrIJDpIlp1O4fhpE5sYxfxPDrH978vCjO5c7trEDrh/LwkADUQcn
Mjr5N/xpLu6mNdaswl8DguMEqJUYgZoITzgT4PXKItDr6OSoH0K9n9aGWaHD6JiS
AhGRvlOVK2XflAEpLgPifExPzR0hN8V5WhbkSVFyI4D2jvhWhWUW14q27SSkfC6u
wZ5VK/W8Ud7dcXSBOzLIukOQ7idqfYUZ3D35Wd4y8S7I+e9mm8Ddw55U5U5+DG+l
G9AG+4QALUYAmUrFdiGdyFP7kEXWm3XjnS78VLeOF4LTCwoFmuVEzHF6vuXKXIYG
HPctBZSZYDgSzCywFHnDo700IF3a7RNmPS5aztCprr0zD1eyzGp3/7QCwqZ6Y9M0
n0NlEeGywWh0t6jbEbuVURXQUmbPKWIYy833nkub1ji77qYoe6RCQ60ryhTnLn/M
6PLLi8MyhPtYVK3PJDX9+g4M+XBEjB4hpxVBDa2+5fkI328FjsDOAv4eAEqrxSZK
ul5/kLqlCf5ad5RISV783TNNn+HZ6TNHR1LfcxcVg3IV07lgAsBWsoEGMiZisApX
RFRWoeMfiED2rHCeYAVAKFSxSNTS7ZNx3X7yl0b9OPQ1tev+/mUg9dwZPxjpX0xv
VfcS9hpD19OvrOlYc5jSLkZhIpT5ZhBnUiZATYS3Z9zqIUvu3pNccwoZ+o59m7FS
gMLjMI4T532IEFCtHTC4/VSR/Iwdp3/p+0ve9S/pPDRvga4zuO0tKO/p1bhmSqMn
crpKiW7LwF+M+a3XOYXGMi0sd9FT68Zt8rcPteW0gX/MFLG4wbD05PZIKUTb/qe5
GF2tbGStiiGcA2iKA1OrbAXF88L7ZCcP4PTQwKRNytjVvNKwnCEK0KXVYWwSvybN
0n4ANJY9ucjnuymSgCKHZo05tTGf6Bb9RioejnbfLgSwxuhwIN5cXL3w6gRUsT9h
79KoJeqdsThCCOBy3KC3UyDb9lkqUhmaM3D2VBeTWdM8Q3qJVFrDT35Ud2+SUbY/
sS5y/CMut9xOh1d/loJuTiTzE+vIrSNUcXLzKjioHiGdv6RJ7rI0d31e/Xq0mXqY
8mWNnIG9JbuJEcXyU6no6bMl5Wre3mFGWXb5WX99cMmMSjg25sANqh5jvA9Wyufp
Pu42PT4SA1nwXEh6/bR0dnbp8gZzZk0c7SStXRWbIcwbxyCNrOb+wYsDZB+CxbGX
DHQlzCYrqbGbRZSdOSTFAzLjrsIcVeqSEhe+ch4dT1RronaEyusXSH/f3OQkO8U1
5Kr72dX1T1gD0Cy9BqBXa6b1V0U/SYLXCSilhwZV66vXjU7Whzmytou4EOpdDj73
5lA125bciOpHN7kBWjIOZiwzmW0UdgmPNZWBLDdHs9ZolnpKJov9HEHr+3nrfZgk
XDdy4wY/PauXmrJf58RKvJHKQFIB1FXgUdnnjur+L4kCFGFGG8UYT393t6FXvBqr
aSMnnGN5MRLEWZBDgUksZsLkb6qSFZRol1z5AysNfGpklV0O25vIlXCkPH2ZpqQi
5oYYobS1jXYtCP3fWdwSB2CxG49Bw1TR+xjS7Yny8kWCwOPVWFfzeECr7Pl4tiQw
zV3CTHEXKs4TO19yqkNrnhvQ0KoxVV8kK0hBheS8AsrDwY6o0FmhgMOCFsp9qJ5F
g01Cjvpr54hYYWSJ++ckSIX4CVZ94872BYkVTkMpvzPEkzTtQHYlTCr89z5rgvKU
Leumo58nL1p0oUDDCyE4oLQEbyipwzp8zqeOepEAfFuHz7pBmuUUS5Jez3Hc2VmQ
ox5V2MIvLwKW1lBzCywvsI3Z4xazBV50W7hH4LUJ4d2Vvk0mgSP7s4LVQJsnbHy6
EVBfd7Nb6RZmMXvqb2/q5+JrwFrorvMepJREti7FftUkLSDQ6QeSmMrVQuhDFwvf
m29CKTEeB+ejxIgZfmZrmgehMtdGbYIV/2mZbwSJXyfRmIENSU4pY+bPsDwBdp/j
+CBX3+Qfc9nb75IxyI4hPwEQSSynpYZMgH/HXVW1k2JfhIaoreX5Ko6DeP8/HfJ6
LpoIKSCtu81viYn2DHdQ4wd9O/p+kXsQM+biCspCRwphd4xn/MZm625A4LXS8VCk
cjk3fBLtVYX9W41I0Vitpl5T5F183FcmWDePaAU1QlnA+nNQ3S0406VdrmT1xl0Y
WZTqBOOXXsU/opego9uFim7batsSUoy3a4PhJ6erFi+sgz4zKWoG+k6HT4yomoW6
rU2V4siuwNXil/jE/kFZDfSyCOjDNNX22Yat1zfObeMzAAbV9X3VeIaQciYZLoXv
77Fevl2FJfe9a9bUzfgZwr95vrNVrZuC9+Qqdai07MwohphDVobKaZnepV3D8JH/
9X70h8kPWQHCacY73PwTY6FUY56/WMpKK/M1ZGuLZJXiSM/yL2P4bLyoD3H5V2Fp
JpFeIPukbvUnkF3FHKPx+n7tpXognl8pW0Yu8dntZtNNwFvOXHeeDeRnsmLhqFOy
5ltesG1eOicahMVzCUeMpeCmISMC9GlOpShgk2XsHjkG2Jj+X34/ks3lUHnQyZO+
LoXVBMh668U4fL8t0bzEBQZNDgCRGC7XAZlnX8MzDueBDemqsiBZUubqCU9lEoT6
OLlO671Fx5oWBwH9v/U0zIKQCZ+BcmqSKRZfyriNyHF72mfhjjjtFpOuUH0vsHb/
Rg6M8IusN6elZrnR0neCogjFNAnl7I8gOLOW1+iEYD7krVi/mSnuz8q3YDvxyj0o
QuKUMU8opuR6SitqoIPs4GVyrd01Jn9jVvEfKvT/QVapdr+IQXmtnbVLu8/oaQLL
FRHB1Qf5cVmV5g2sdzM9UVUmM26SXpuLR14dbL8EzjrI06LNWq+/JfawqGcPNW7O
9yvIOm9gHxYeMNBjj+kJWaPXwumGF8/fEAb+I/KUs82CDvVIZmRHvo8TKuH133oC
HkqcaSPWHRtQQ7FNOJ73VibX77x1QIg+SgLsyhakYeIGYVUBqSvR9Bnea+ggoE2/
lNCAL3Fbh5YJw+ih06Bvaik+xjMcOEQ0ejh2UOWFya8HtaLJyd6u2iJk9JAReLG/
AhPgbQHdGC7/cbWucmwHi2lT0TOXu0JnW+30xjLthGtscWuHoSpAMElCWg8kc249
YmmzfGCiuiAGbYNlFIh/lWb5SUAU39r1L6npcluZ7MWPPjkIVUHUfasyBJ3ZaAWQ
9nP/j61SD1Z0lyUnDmliiUHGeFkJ2TrTWEO0ZyBqeaZx0dxL4cpeM0se3HEEwhII
ErPokzKFrzXwdLRY1lYOSvX7/Kq4yv5O7JchfRyo3afwAri1KVCcd2SB7i+qjPPm
jIE2snfQzmOBxHQbe4RtE1bKNNd73z+hvgRAlOiy1DS9sxWRXX6uLVDK9x2J/b6v
ChdivVjPFwKtYh+JC1bw+/iQdHzzAD9AbSMMu8qopUwCU5oh2aP50ACJf3PY0c3s
SdMNiIbyPlSHFy8Zq4ChjsK8bkGkDr9S+jX+0VkNX2MMWyRrHdJSVbGYLePi8QWa
3kCddHIcZSvW46fVlkk3wvhAJbA1VnDpKNm1fkHTyOq/m92Jx7RIcfZYsBTO0Dsl
jalLUsUhCqQ2HjHK+SOzRtJlNEidZvwInLUmBJdrXISs3RgkiKOjzbXWCBGLO+Zq
nTsDOu5iUjWsJ8SpuxoQjd3JzrUZ59GyZx/KGIHQz1390PLAgRwKme76+KRjMa3+
cIxkxQbhqwJZ5YPjqgLIlQYwhftWVF3g79xM9OoirkigW+uxztf8haviFEJ6SXXw
m7W7d85PCPVilDtamnc4aNptcRUHSjVJj/Hoqwi1uTuQveU8tgci94hOK7Ujbamb
h9vNlx1trdzJxYYyHjrLXUNnzHf6+sVvjMg8oqUoqYeXKpZFPqcyOAb6qHgDEUcO
UiGQUhSpVqiQeYxwTmW8DKPKFq2zH6racZutS8AL9FeClwiPEaAK1wjpWTSyub9k
7Y+a9nEffZju+ALPlZh0nJswEPkB+uZGxOyjyPIruaGzo90IssZ0ygJUMLF5pc3Z
GBjrXR9clwCmGuG+ipXOuvBtkO+OPeJO26Vh7QtRh1JfDcaw9buYFhJXbj48eTxE
A8g3LHcaBSJNPZ7rimbW8ESncRJj99Epa5pPa/6BfS0uG1rE9gcy0HqR6MaDWiiw
B6A4NBzpVev4FIzA2y9IGXgrwLHXPWj6H3lAZGfGivcw7gCxJ7/Y0ZFpM7bWcoqx
sexgD/r4FIgb0goH5BNw3hdS7w0V8ASvJ4LYrlTf9tnBJkyVUc2RDmcvbowlK/6L
iZWoOx+QkFrloNlUSTOdGwV5dqN6zhJtLmoM8qOumqX8QSSlblbJaKsRCKRYIyml
ny8tiBMM1VhdDJv/xC8I/QX9RvhoiHodacZ+FfPx6xq/oxvAWjveCJKjsH6KEqSC
g9+F3VCUV2DukKhvogFL4bLogsR02MJVJy1AYIfwu39gs7iy0rZirwl6nd8e1eBf
iUN4Fn80rWBc0J9cY77tDBCj5sSGc42b1OpqpseYjGy9Ga9iULrNfsB894l7RVd+
Z7n+n+w0OS6i9A1sGKrvaJzN090i3UKIJHZPhjc7gXJr3YB8+PClNkedNxB/M7J/
73lg9oReWWlAt0Ib0AsJqBadl+dE+HvjfM0RjmL8VJWCmflRFPbRuXhw+NAV9sG+
oYZBu/I6oxpTiR1BJvdm89QbLgLArSyRIZpPadQ6ePp2pFqNI7s5fPbwn/Mlv/Xq
zH6DMXH2SNvI3YmG27psXlsb3/oM8hkQvoeKIRqDuN0QwNSc9wBVkxs+Bfltz9D5
z2vuXWgIbkwjRqJtSKjtAm7mjuoHa4N1/1QQNdfRJpJg6m0Gge265Ey3HMZuyTAi
91qnTjx6Zq1RP5SxNjDeJ+t09uYl8GVLjOgWRJbTJiOSdqn6HzA1I2fZRAOqodf5
AX6om1iMSKeFTN6vwjUXmVhNan4VAJtYHBNN4LWH60GBrYqiAQKIVHyk8lOibI5I
6OmuaN7dxwPPSEMcFh6O8uJKtXDl5AaNgVdsrDtuUi5SJXXxYvbOruToWZED8E8S
yoJ6TQnFPJQugHUTMIJSguTYygLA8QwPbsZoegFAODAEU7pyuqKK/vl1LWtYbxSs
iPqigWom6Zt1lW5l2ZKeKh8VXDEUUnraaUNGZaVzxVVEv6NuULgGaziwZmvEks1N
2cOv05Ar3v8ANygLBhzlkL+p18HfKc7tKUBZaGNBQ1TbZhfAhPX17LYEdYrm62+b
WM7PAXddh/U4Bb7OY+8qAPEUHnKvXccyxVQbVpWia8O/3UWVKRvcJJjFzkdOiU3O
zB4ffI+gmfBHoE/U4JPCwBIjMJ/YufZuYYKqdZAo6ipUvbJofhcs+ozM+GLlHvSw
DA1iA3cKTJigexl8nlolfOjt+hRwBNCV8Gr9p43ItczKQni0gq6kwx14MZCawTwv
BKBUoaJGIIaNz/teXOYqpGYDH+hVaxLjVvoDq4lJ1lMqMn5KIkWKgxvATdpMdVeF
obnHdbetXYpq1wDbPVi7dkjZEndd/zNsihs2llTzKzBFTyz1WDx0qih72vPm2r1S
n2gjhkeppiJ8gsyPDXP5jllSbX8b7FOS14fe3nb+F3lrxpKiWKS7HSKmrhTAK3BC
QoKV1IDjyhWdbGeDjkshQgq02hGPsM7+0CBJqxPJKA8AJNiA9xf3qzhf7ypYlS6C
ls0FlArAAnTYR9SRod/xw5ULcFKdmU8wPElDMWBg5n3PoHNFxmeJavBsTi1yNlV+
qQg/6LM0YW7sjuoDESh+pKaaPWI/kq0ov8VSeXxzvgJQVi22ELmECfnAOVg1+yov
YwCBnbBiPBRuu10YYqN6zNACfCSNbVBHYeRoMpl/ock6+QtxsOK0bEb2cYrx9Xek
3sOSvBIcuzS4f8pSk8sDs/iZZnLJTgIKo9PFdpQEa7Liuhxgk2BjeY1MPkYyZV3U
9brL71PPNjq0Fg4EzF3NEo/G47aWUZ2iGmV8+WTfL/TV+JgS8tSQ3K1yz/RS4E49
p/6X95w/Xebrw1Jn0siOm036Od9mTGQTpWqC1BTB9slug+H41Gq3oayaOB7kTYS4
w06WGILIVCilroU8f9onWSQ2kws6swTFHBY4z7kwaUuaFWUuiJDTOdUTmTgwk6DJ
XBU1AMd4UsTHt+DkPGHEKUb199W1OCHN4o60IUTNsxagnAxmf0/czTvfrzYjDsYx
QOoKN8OGRKYXzy4RPbnCFRG38Bcyi/tXGIGVbErYI2uItszxcK4GNRmsCXiUhqfu
K6cOb+LfW8AzLe1HvCUKfOGAQK75mTmJLZ52eSK3nlK3MmF76FQExD/QzqrZxybq
UUNbENfbM0LCQfixv6SP4sv1Q39HoO6NSYNBpLCbalPGlZZTKRCazGw8kyZBSQMe
RtDh2X7Q8Tv2K1rouyEqZqLwYX763Y1L7dFM3UFmL3sHIg0SCZzc9EmlYnmAorDz
pGImmalwSoO9HYF+hF2qdSFRr9TAFNgi7rOk2NeKcKuHq6hC06m+3cCJf2s1bd2a
s3ncmM1/OFko7AjXgfwzJNlqZFEj9rh3on9n8pzM5vQW+1ey8uL0kSwiTAxB1LAt
1fnVnG5BIuRt2aKwMRSy5nbFwTk4rVYUhPJOYg/cgNcLbzYEHgYcXH6Oq3BsqyD5
zB3K6+WnrtxuF6fcTSE1o1gnS7AY3BX6NaHw67FSRwms/n6e2EoYDp2IKx7ArQP4
QW9bHJHEMQSslxjpi8CTCeYJaWvlHX1UENVDgZceqDrDJyJKqb5uymJaL0hAKfFj
PVtquHMIGEzt+kOscur3cB1OxnpmCotaWThWGXEO1StAs4VYwe+6sthmei3KRlbg
ju+9qPsyc22LhwluNixQxJ4gxTS07ZbzhFpnhM2QFJbEgh3Pu1MfANC/NpP8zp6X
KM7Gr4zQwrwA4QD68zZnlVTi6ZeLpKl6j5IUFUXchyndCENAfGzyAVCUzvvpoJU6
1txyXz/xgfI/5oV8rjGTAgUn/Eo7Nk8mNa4q3ARl7GMfrRkK48y4cjcq+j2YghyW
tsgdvCjYQvjGvbzv79rqYsygyJPFiKu4gvUePtlc5zjkZVyVIC3jMpVBWjL4h+ZJ
K7isW27kVE8J6pDlfHAozRhvB47RRA3uvgTpff8TD5CsZe5SjS2bl06uLXnjMbgE
BR8HedPF6KGRgWCR2ZRQbkcxiQXqp0KUfFujRfyfE6d3VAOQaj3l/FWbFGG30Bca
RR2DI8q8kITDeE0DJD69CaL9VImMSr+Q2XKRgQmZfp8eA7bTj7J3OSNvgPICvxfv
5dwd7zCNnv+5VbpJRSHokCnS8OoTJkNYGgV8dyiv7vDyJwLPHWvXIuRemt4iF2U1
SoScsvByUT7JohNOAKGt+R9IKgQjaSD+8dnm7d4Q/0zTdZrTOakHwP1i9vDELkrk
p032f+ZeE3zzXyTsKZApZylygAVxU/25L6BfAhTxKD0kIEeJP+xnMuMgvISps04h
MXBi0LNvWYPefWXRXlr6KjnRSz83n657vXyAi5tAW+j4nrBLwgC5aKsLDsRHQ90y
qZBn14jNU9s4ObwUIA5CnLazq/zQRscde8L4dX7PHjfWEcpUaFKECwycOsOyAjd8
yKFgx725WM1rIoPf5JHg6fADTmFV0pJ7Ca/4SXZpjYfMYOe1AogPX7F5NpTpoSt4
KLtvKoKUH17hLWKl6AVnzgrM1BCiTBkrKYwNteq9NsSf2IAAVoW6Sro+zFPjqFFW
/4ftW/QOGQOn/Tw8V8AimruPVjVxMrrJ6WxftWhJAiDGokbL8wuAOVa7OXWKpygF
6u+8sW/HXgG+zoxuCCfkNU+srqigKpyjrLeibFg74RssZa0bXfAN5yW2bzukd1JT
QjkrqUTHB+6FxxHI/6tXpBJ3+tB2btHMXZ6h2Z8G4fsTVAKxPcguNJXPoORwfJUz
o47ku3nvBazX15NtAtu7abC7gv83w1a1kJv240jBGqMgvKT6ejPc1PqNNNkZhgVI
P29iNzU18kySFx9ld7iWBc5Qjpjcme4WCF6mb+fpDhk7Z37dB5/ZvqUo4ID3URyN
c7a4r/kMkNRnTlkXhwhSz49LHKRRY+XO2UdNki6LZBlFFi0obb0x64LwgiPn2rmn
ewneBiWcyCNe24ZkQgpHla40/FB4xzCxw30MrtfP2oyZxWAlce6kkpl76JowJ72y
Gq9NPB6/PvFG3dy4ZDe0Ol30mfSrhPBzuvMpr/96BkmTmC1T7+nziHa94YPwjnH1
B46ugIGlpFc4sYxZDQJ72UWElTUu+50h0SGA3mnSsbhs23yDK58KWYGf+PaN22k4
qzSBvvz+PS7aTLeBg8NItZpCp/F4yT4crmPlm3MxGgms+5qhAfEeeKFPvBl3Kgnh
tfNSokbQ2uELmp7odtsC3G5K7aY2aiKDIXZT8bWdd4oJggRa32G2Pr8BRs2ez4OP
x6oqqLr1R/otTz7ilENtDZdE4BRCruyPRwc1uAypHi6GsIkLZCMljxjYGl98MnB8
z941cp4fweJQh6Y67ntIHpt8oFB4Er7J6flwwsK/uSq9nvDec/4bFMSzFk0mg9DS
pbLSJYlvrVUUVSOC5uMJj8+00JJO4cWayj1tujZge6oxhZHQ6iF0aUF03hAAorzk
17HRghjQSVRe1wBYn00QFH4W6iQ/PqFWGFgjs/KhA8boVXUdVWYyfwadTSfQad2E
hnAt2KTl1vXNQjKRCz+lIPpB1gg8Vvpj3u+kW/YP23Ob3Hp28uzNeCxHyap5/2D7
+dbhrrxTa3BVHvyosp+rn13IyP/fVClar7GDnOzADgokU6ACi9ecrYZx6QJAcjYO
oc7E8T7EihEPL1RmNjYmQsWChu+wrGHNhEGf1LpquSW0M0JpKZiH6BwTDTxtUOLN
Ex8TrtK7FeVi8f3aPg12hDhzL+F4RPisj5g7izFEvX7nVDkIuVZMJD/PnKmaWZul
OUNiUSvmeADh9qtH6AvGjV+feqz8KAqx5CazmqAZbw5BuTwRUZ7LSTb94zNGKLWt
YRByJKwnLl88Owd73mSFRjkCqiR8wpk/c/iPD54Wtaz8flsUCkI+4fhc0zw8IrKH
AE7jC3mcfUeaqW719CATvstm/oG4KEd8koqVBGGtVlJVrwYQEgvCjCR5ZnyiZNyN
ZDYxeIF46Lf2+zsoMCwRDRqDkDTeSAF4xOdcjnx1JNYFFFluFaGT6VSKUZV97Egh
1FIq63GKuPv2easzOwRn/XKhpqL2QTpjBRS5ATnRxvQLQJtQin8uI/rWFL7wng1+
Dt/zvRpU8XmuCnDETEDM+kWkKGnDT4RK6//khSAg92nJ2aboObJhI0x8gMNNw2Mz
lon1T9hxZ2rRJ9pAQlRR1ENef+BwIwTOi/G16lOJdVGP8oZGHR8hy+lk+YK/fUuo
vETNzeM8vFTX+5Wn1a/r4KcSBS9Fzuethz/mVREdWz7u1MVxWImINaQ8nqDuqdOu
Od30J+B9kiQfW4q+Lyrxqp10EEM0kUWiseBHQcj3DLT1plM6nWQsC7ZxP9vMGLd1
bg7X5f9cc00Hl6p13zJfnk/VQ7ERg0+6w4dgKEa8TmD4MNKzt1DgHDO1Aw0+SOp/
1n8oMfDDWLhcXnLoU1t40HywYdlWPLMLhRWwteFMqxGnLIe6WW5JsnSMC+PwGuuD
adZ/DGzUyL/3BvSLscKus14APznamXRROIwtCR1j4iOyq2XYicMEcWPyst3xDmbF
QuREKpu36Tl96QqzYdEZKEawVHH63fglTPFUkEieysChpPe8U75o1WRAvcL1Sye3
d5ysDo9P4E6WCRuIENk4fRFfXYbiSGL0gV9KOhn1naKiUklt7ICf/5HLiqgCg6+K
cZklZE8IdAJeo/REwRm7IHlYp7TEy/s86xhlyb8Zij4koIafKM2AabgHIyWTKd6v
7j1HUv/C/9N3e2rNYbMVbxAS0tuSmxhHPqPg8kiJOnPXSKOV0CZPGM9bEX076HVc
I3rZEOkkZEiStex2lyQ0AfQSugfR41n2yK/Ml5jhaEne7nCWCr2dvUttW3ZBITeV
T2dvo9zBwiQacOFpPnwwRW5LKVFhOVVO0GkxdKFffLwpydUOoe8Sb0QHf1ia1lJN
QgoNhLDYcICm+BeQRxTt1hMxkU28csGGYK2dD+2m/QX1ctNm/I5HPyOaUWCITK/P
O7+FwapeMpZKhhOtTXfyN84/tX++c6T6WDP1RbyIr67wAXWxvUO7UH4gEesetKNX
WnyM7yBKICt0RyqZ9HOYf+yl/TndTD6H/cI/RPJg/3c4n38O3XptdovXvz/bIKCT
eTurNV5DBGyQ+p4vrs6n0Z+/GFngvWmh3eFpJJxRSu0e0MGo4xgHSaCg1HtbCVi/
a6rHbET781FIAtqGD3LAUz6+hpmospB67+GaxwKNmF8pPAQwd8aKowR5LPoai234
TfWktIXi6fRiS5eFDAbDLJICaFk9z4LfHEZlxlF5vPDeieF4qTkytEaCJ/8A4g0c
Fdwlq3fnkRhJCqIfokxYEnrAMT56UdjaBkCs/5P2GaWKcnmiq18s31ZjdAec4EIT
F+Csr+tkM6hCXGfXnwnLfu2fE0239C7TM7imqkWutb3dD1IeMpN8N3v/aS+WFpw2
6j/kziv4Kh67UHlUTsCCry9qTAk55JLuBm3s8Oy9VSRNu65WabFGugPJtB139VsS
c2fiVmNPbIRrqmGsYGU/YSbBKb/yHMDYRxLsdYHHR6SWpVsATZFrnWBjOKGpp7kf
u3l97S3I1oWwkmXZIyb+pPRg8l+ef+hieFBk+a5UdN3zJpP6byQ919kqF5WV84Q0
CyH6kzcNNCUFSoeUlDdJlgDXuMUPbqKP5IJ0WgPSxgd8VSjLwtOikMSRi/n58rn/
0d6EBqTdWui9BjsbZymhyntFN+33P0/6Yw0eq63ZgA59Wgvj0Awbe+qxvu2+duSK
95tC6julStDIBGT7USSlol8y0itGJ9ygPKRCXrP3Aozq0xwObe/l0z+cXlfoHXN3
jU3pgpyJ7QErelW4jyx50G6ZwNkRq0kHR/ne22+Z2ms4FLYpYJcgQkZt05weeLDF
Hg6+EvVNWZAatn7JooxWJVz6z/rn/E5doa/eW2aaAzPUXoJ9cZIEl4s/y7URNtYT
HownnP/Oo8LMoVFmMjFOT661uSbZLFR6NofHoj+H7l4apufPADFXJGqDNGnur1wu
Imtuf6in9oZCGrN5PBBb2SoWvJOaO2HBND1vLEAcF3oeQmcnvcZXo3d117wmXu/g
O/egdD5gRr6TZRE0j1yUrwL+/NQwtkgReNuoCz/uDhf44urZg0z7DoNwU7ag8cgA
G5QQGUxRV12soc4qeMzGW9gfJ6PbpwEd7IZLdHAHGTGFq3AUu5ND49TD7RVBxvdU
KX3c/dEWNOkH/SZ6BZjGIxrS/nDM7RVuf9bP9IDcCJAKfy40J70NB9mgqUXAC7bV
mJiV6kD9W/6oxHBOXyj4BUNHo+Eu0zENqEJx2V38g2teXY2vpegvLcpdpUmc3v2I
EeWFKGZAbI5o0F8xjvpVU0vEdrabvKB4r5EkPRnBA+C95m3BARwdJBYYD4D/iYtq
38fwqgJ2S9knMI7DDwS//RPww0qtHLihiFB952IJ6yNwplVf9uHvQQG9wnjHvBZV
x89csCWN1guIeCjULYhbxWsWHOl4ZaJ+O4XszriMo5KBDdegknReTUjP4NIlyo49
z+47Nw9hz5YoCTjujyR1km4x0OtxiewsQgRzJA8kzBP0XDON8kBlMiHOVYSs6Oqb
YIaKzBvoEVE4EgYTzqeeZWm8BiGzxhexiFFyr6KAqvtWVhcNrW8JAf+mdcGXyORR
DZdijTqrs6AJf7GZ3gctnV1MhKUTaTa5o3WKpqQ1MY7OUdjSuTGTGhU5OJM0ucqE
LLRlZE1HTICG6e6S91DwJ/7wivVEk9NDYqayVGEUdraayvGIx3i548aCsiri4YbB
x06FzXgu4P9hVS1bNoOzMNk95h4ptt8w6eAYariM3unQvI41HYkn5VL9eMu+2rkC
voDqOuOk+g4iwFia+Jx66wYj3ReYsIyA4omYdvHfMxQB613hCUTMhPRvvKTDuyqT
wGkZAsVCr9YB8hqqxrdFIBIidgWf8AMG6NbheHWUmjoMXs7vM8C4dj7scE+KHS0F
u53vHz626R1RUbkeertujwfCWzOouN7r2hxfWkbY6ysIOsBigSWlP3G07krM13EY
MtOWb4G1o1ndkZzOPoy8iHb+O9iFyy2Ode0s+qxluAIwXRJI5Geywr6e5bVNPUan
quahjRz6wpObhEZLglG06FXHD5GLZQkKTRkQ+PWsSU+MS74TDFvslkZvbsMiFt7J
wZRlGDKpTppLCao6F5PKL8P6gC9lLILoGiDLCi1n3sLkWZxxAh15GslKg9BaebHw
ial7yIS/fng7p/3hvQTvSPtn/PGgOoOs5JyOtc2LF4gwEzzVxQee9DUCF5ybkbuj
ZjaYLEaFc8aRjw7tFPspG6feJGRpUyvkVw5rbkuHqjIOEHnknqDyh+TrVwg4r3tm
hbsbgqeO7YrMNM6NfO3TVAHoO1QPL3a8EG2KnTER8NihlQsPPreV5XHMKBE6Nww/
jLyxzfZGSCS6GVMqwoMA8HZ8POJ66FkOJu4P1rJYzYElPAM1dIj2YZb8cKe+UNCN
bTF/q24yoXtwaEv4+aq4qR+uiyHqvXz/Xnyw9PsrNwI+RyWKA9Tilg5LZaS8DK5I
eV4bRFE6bs/KRmppQj5qopmrWzN7CvxJC8nI8BanlonO/iK27R84G77RxQy7c+Vp
vxG9/PuV6qDAHC6oG2wWTkl0CXUvDJNw9kErECWSFJkff6zWW2U/pHWvjGEHcd0a
KQoaI16lKrF8SgD/wDDIphZWcgw8xXAqzC0ymygFq00UbaFgCEFg5cdn83+r4fUs
UbnYNBs6xgVIeRQ8JexAPWW4HxOj8VugF1GYaZ+pRJj/kqTE2OgPNZbh5nRURtpL
19Iwi6Fxd2hlrj5RfhvawkNEBy6P/NpjoorGnfToh5Pv/J/Li87ggEokS25gIba8
0MZ2pyhAnzlfOTUT9nJ/D/i4OL2tb4rH40l1Y2Go0eIzKgNZWv7Dpy6+hQKMJggx
oPn8Tpj5kyYOGAlI/jU1M6BgDfbt4ZcctiOFqUAy12SHncd+AWfoqXz8xTPwfbmI
KAzJqiKG25yu/aoqgnh7T20QISutZVtEEMxKFpiqMwg0Aikf0nNlctjb8jTATFDz
27/L4yjDgCqEFxmovfjlyLYzgO3lh6oMxivFesRlLOggZdiVHZEGosLXylcMy7iv
hT9R3oo2fAbwWHR6n71UP4KSoaQCcODshxv/545suKt7Rx8QyWGIpwj5tWOq9bm1
vhMd5AKLwjqVI7js27DjDxM3GAsYLXaDP68hrov384zei4KYAiXclfaj6OWx8w9V
Vwy/zcaNlHJuNtgXQd18Z54YZSCeMdcXVVGoU8zQlDx0EVFsibPKN7RN5W91inLa
YBbNkE5PtKvYtwpzUS/Ief9084LLQ3Av+/JrsYXNfwyAvKmdPNCOnkIYUBFF2/E8
JdVm5X5S5p32D7+fO6P+OPJC+jgcVSS0uz9tgl684gEtB3j3bLjPrMuuTILxFdhg
TRah7TGT6TFru+21la7nBu/0mS88VR/KN5cT0VwbdGsEgBI5xN15ICqpyFeAu3GV
paX+XwYE0y2BGtKAQnilkCmbkbMAbKrv0INRno5zt6S4raO/tRNyocQOMBgnoOzg
SkJ1ucIupt7DDGE3v/wTyxbvynPqA1EvuilUgoc/HO0m6U2n33VpC0xfSIiCbU5h
d39jRcWb3ILPowuKv2bIGDvXHBLWCegSD/vvZCJddKcwA7jNbL1lhuXCt/nL4Xqy
ND77IhwZzln6G/PhTDHz3NPZobldnyrnFhbP0sz+HY28+2ZDAWwNxga64UVqDzmM
fHpmvAte13VVux4WejUQs5pcg37+E5s7BbMb4BxvQoxdvhK0ymnRqpsIrZMQHMan
s64HVeVKYLRR0dqPd75yrQCMcDJWwEtHp5vtKAqT39isGot9meOqm6ut/U9zIsmA
/1ikpAxBr3OAv9hInfzDjLuyaq1OGK+o8XtaS8G0itP2Ub96vjNryotR1H5jXKZI
/j5jUfahg/9VWDd3rAcuDGTHlNlxyxv+XdfU67hjKgW4SQtGJpw4ehzoUuydJgn5
qBRbP7cyi6RCCXf80R4MyOtinmwpUlOeJEl6JH6kVIjt8ZWspDQX35PmWCu+1y7x
CElZe6Rwbr32/WL/S0JeoK3lwpAZOw08v5+eFC6Kpv1sWBoQ3aSnJkP2P9/+vs9H
PBRUg6IC+S0IPueKb65xE6qn52p/oOC/CTtFPn+4iK7ng0Ef2SFP7ymO/7+rHYwP
D+ZnZ4G572u3m1/F8/uAzPqb0ti5zsRBjKEOnCQXp/MFeyGtNMIyAuJPdnekWkc9
Pz+CQVH2PpzH82wvlrQ9HQAYFuWVfqsXwGbmnazQl6wuRuNMlByxKyf86UidLpIt
0PQPeB59d4HaHSdaoQZ7nApTdlzG6Vkm2tilK5sLm7qb3MSmkgYRrx8hjLPQA8LM
wArQ69uMEy/U2HtUpYrjkdbfjsitK1DYHK5X+BJZPoyZfzp6dKAKvFKoWy6sLrQ/
FAl/d2EC8gzcEFyHaOuqaoXtk+4oeU3wnQXB4HW16GLyyW0sHtVnc0jja7NfYoh6
FLFL7VyxhdS+yrgZLS4c+7hTDsijZsUUN7oK6htfaLX0f56LP4/XN7aFPfSFsbnm
Gt/PFFKXZgaoc/+qdv+mYSUnyJXfXiqpHllXUjgipcAwut4VeV9AaPKTkSfCSYSz
9SYEekNzeDMoO1mjbWhVzbPkVaehrLIIJuUPRNLf24p33FCQSjEQYzzKrBVpkZJk
Q2COAvc5q/VA0Yk2ndPlfaEEptYi4S208Nrpq59g8RwzDNTU8oJK/wJvtle/Kgyv
p5jDUrzDWEg5HDGZtTRgxwubNNOwgWaVkQJeAUqnzRtJhWn3oWkJu5XRqfygUrP3
4ruk6OKCaK8VgnIwAaLz0CglaP366elZtR2uzxYFWIK4Hlxff72S5aR0qm0gXG3e
Fe7W2wkVaOojieLEjhcDjhZ25PWvP+5mflYO40+a6KWBtvRfqoPjdysugNf56XtR
OQM2qmbYphydjPO24dpKO+Z9De23w1+BymzN8ZJBHiYL3ZMPQpU3TcjgdzOCv834
DhM7QtwJ1tbWr5vqxbpVUMBjccrjhrWIPqcVvlUAC4JkSsn5/F0ngsQve/UeyzJc
H2t5dKkVtvmg++ARe+6SOOewCH6DhFPq57KZw+VV+E0A304vp/wHPjqH7Bc0oaef
DYCY6exc80vuSaZlvIz2YO5EBIdUz8g8ptKHtPr4XSjjC2TZ8mXEzeH3y/XTIgwt
TunD5nPmbfBoLjqoZDBFHF5AdhbuZRe9nhFk6MXSCJ4dYQhzwFhVZv2+JhkaH1bF
ajC1VPPajT8nEKvCF83XapWSTd4ltUSuKUC3tNcYfFaLRSvKRYbHLFEu1PZpZGZv
3P64v9R8eN41Zh25T3yt/W7F0D9TidjOZvX67ro4r6r19p51zneiB4m1wXJPKOSp
aAmASXKPDxeNB45yeLmNdC4ys9Au+BybDeqFHvcNzWsYHmy1zSLXRa+LLpGOfmOV
JVC4XUnhZxGNpDx6ufk+0Fpytnd+baxfXy2xCo2vPfw6MjpKr8PrOI3co+l9MSqU
sHwKniowba++zi5BCSPUV4F7/ZwL/ndGgw5g6NFU6dOfErABnwjyzrea+5Mxz9fi
uPb3z63fVu5yH01dXImIP58Vrjxncs9YkIPgv5CIUOjXdSjmYw0LGZpPpGOtreaZ
2chftI9K6QwsKOsR9GHYNRGAsdxKOqp+Rcl5n1dSjb0gYgw9GCnVOFwna1W8yu6y
7MqbYwqL39HOtsvWADRtSRPvVclMHJJJ8jAjypsH/8gMEvTZwOCkEiGxZsurwo2D
/A0a/mHRGNoB/UOkIQ/VkNm4y/9cTxhNSxrMPdZSPbBt5VGwOVas0dQt2i/LWUVi
s62PlITASqh4vOhb4nUKdSiCe1Ze4Mb8peOj1cJkSWul3+drDxgt/ymWWyYXwQGg
NvUFHIsB5FuZKzl+RGiMB87afb91lE4ayLpAjhIJg9LakEcMacUx8eHpegNCVUAK
S3Ux5cZu78bZQ6oOTQaCocbnYNyFKCT3+OlEafqnc2gwLXfyjuQMhO6Y1n/fWW4O
PF0tTbiaFoumEx14wLAf/837kBzvul1oFKZFULjoU0kmg+8HfMj84Ck3eyQGJkrO
ozPQ7Dyt8AlNW22JJYDhESNN0iBJ1d2rE4hGgFJjRH2CVUPgTm8XjyRvR7yeesZr
/N9l9UXwyZ7b4hKyBqdC1lST5BK50m1p8ctVyl2IYeMlh1JOks1TE6fz2tzpj7kC
1UAYEtSZ3+q30y1VVWdDWQWWlovEMXvPRbfHCg6lKU540wuYNDGmMQMbf85m/30z
FncPD74atbkTZIbUYQ7GYQ67WxN1YnDdJASiRhY9/Z7S1/pQKTmwvO8qI3qejp/R
6p929zqXnd452ImaJmoXra7sLHcS+yGjwQ273TXGidwoLNC1luhw096yfAuZn0hE
m4CCYFBgCBtr8vKT63Te/6pOq3vyJ4HYeOvVmiKghkeAu42AqC7aIlAURK7O2HPF
qwFd5gotWxe9TslWknp8erM6NZ3/G6CvewsLiFftN4jj+l9rGVJAOF+D8ZWkg9oT
KECNQzrkO/sXz4POxuEWNBk8+5D6Y+0r+SMQiEOtYuEqDuHRilAUzZ+KEXN7Odsx
KgxCxLtkBwcIwH1Bsrb/ujm6g6Ptcn+7/MrewOrmVKunOAi96mFwEMvUJayPK7yl
tilyKUzvdBmSZY2jcYPickaWIjSPLDmFgzAoFMzFOFGmu7VlXNVZCGNgsyTciln/
Mw1QDyGawNQ8oHcbTP6sOnw5N8unzawjvOGwgpZjF/w6U+sGYgjI5576oODD3ZQ9
jnYIDbUdAPPhQlhiKlTTZGbVivE7d1+1HJfsHSv3GPC/Y/EnsVCIus+lnAuiuOtQ
yispaas0ZisOZRLQC7KDcQnDCSUpMhuhCTT3DEqed5w6FsQHk66Hyxwt3A6YPKwq
5hvlSFf4gRZeDgkWLIXmU4TbozHSBtQEEUE1ttw2bHDq6DJd4NDy8J+Vm+Xgr516
qu3Jjq4mnoV5/v6Kd4tLiSV+6+fSSYPDPctnN1c9GzvIaXYynUAMZ9bcJujlH+ov
oSkC8OJFDB/opgBreLWho5hBIXF+ng32YbGDTsElznypfijktn2XHurdPm1QopDE
knqnUQ09T448ExnsYibmcVWy5ppkYWBlPFZEQhQMnqHdCg0wl36ejtDHrIx/6ckq
zZ5UK3S1x5rYZZY4RoasmbXrDyjzF4Pv4s+5rj1ncsVXz0/TIl0GhUzYoi9Uid+1
9Rd9P0ISlu2zQOhR+J2Z3VUWmLU+nX7nlV1ZUO/95nA1xJeN3vxkBO2PFMB2It1q
TewSsqN+UzxguTZH/ZYQXpkQB1nzSKtqYHcs6BwFl9wIljh8knXzp3MdMKwuQrJz
4sGofYck+ys5kr0W8jEXBU7VDZ2KADHHDLeRiTuLTo3WWEc9ZK4ksXruoNg7qfpA
wTfuNTexR7hOVaD/8Fyj1ybbxdHUTeHJ3gw4bj+4LQHs0JLqz+9G9D1bINPmMVhs
CbUfdMqBDa0//6u7TOUcVTSP9JS2dhnadz2Btt0k6nEVFizg7UsEzLxPoneZKXTL
KuQOVcuVu2IdV/ztXhXhzU/73tLwE/8S3dJupTM1MmuVofZrdg1CLadSyRDK14Rp
RoSwvhwtFfG+1CMwC24yLym7vthlB/O05jPSrYRrOegaWyWYhS/23stQa3vy53io
HcRTesaxPaMJC3LmsNPX9f4KR3nr5uO6SmBJhtFgkpDFI4dHDQ5sPmaz9aT2QVPz
OBCUcEMsk53T3uteRbIvsFeFvBBtLqnG9v64tWpwczXQs/7C3pHpHZ7/uMPMXQKH
UZ5215f5mO2zxnzRhBOI3ccp+w0v2FA7txalK3HqLsqBefBV9BoWKwzjfPDJ+cuk
U2G6QVS1JYxnxxb2sg3O2YhemM5FCTMmPYaIWiwrqWvMRFwzpyGDxkhrXi4JDByd
UarlpUP0FGOEe5HrmPZpY1tlAoMFtKJ1FW4RI2ghKSCMNn1TLDtAXT9WT82fpWIl
R3AcqTiFJy5Wk1WRd8N++Fao5QKIj4Me3GUmWj94SkXvH8wKNvwxXG+WNXIUi3uc
PtHaPJJglXg5A8o5QjaXJVcd73vpRc4PQq38yLfENVLZclKQKVCMm9E9R0HsA1zd
INH3bzqaOlaJUMXp/KwbRrNcW54oGU8XtJVeroshV+vGK50a6lfqdDO+5PP7+RD0
TtLtCPs7v8jBzdwO3bu6dahFiaUH6pD96jisurgxkhGyrh/lI+Zq3Go4DzCUxr15
SjcThl2LLBH/z5yEiG76XpTLzZnK4q2DUNDHBpS6Uu6o9hBfqzDe8odLcVgdxf79
mzTtgje1rBRnNDnGPjC8oz6XZ98qI52yZNoBBYNWBlpCaM1BEsT43w07OKChDlg2
b1VBt/qpYW5jVdCQsnQXwqjgO+Z/P/OgnVOrpqRmcTsXSGo/FLB/+TzmDicYKYYw
Xal2HwWxgSVN42rdOl4INgq6UyDwdzskowJ3udM/27eZObf6pMCm2tMxxnUjBMoc
PPus+9M1LeCCYFLMNmiowyyDpKU2/C58dyUSypcz1BqZ3Ku4Dx2iH9HdW0R5hjyg
tNxtl5zGTz0ujowO+ia9/9QXcG5Ph/6lirTG88we085g+Xnb+FuANrG6AdyRdLET
qWJk6/38nOcCsbPW8UqbK/6VCQuxu/SGpknHax7pMqPuBQp15RtqZqH09GfG7yGn
6KQvNpLxQbQygcWkFgr9QuY+/8mkB4TfI2DnEjriNHcxbOU9vh3CIri291gYxqQ+
lIPeh0NKkLkypNyG7z7E1u/Pue5DCvae3lVsu3PB2XJZV7UiRGPU6u4/IThPuc2q
d4O+fNicvlTojGFg9qLD7W4LJv9QvVtX2ZjJYZ783UiziIoQkRe1DOD78KWsqTHi
IIMTNDARBhuiBwhlK34ee0SjT0CkL2X0eg/MBw4CCNPN9lO1zEnkcN4tjA8+gKhy
mZo3aBK2xp525pGAcyzHtkHRmOk7Jlxfg5oo6TxBm+KTlMMNIRSdFroweY/dwun4
bCFPEY9BLMqcKMcobwZojtM+eU06A9+tFCcgUT0G5WLWCFhcjaB2VBeUp0hWpy/3
UA3S+h40AG82CRokoaeZK6eUZJVNMjQJvalCpCVHsdzmSXPOrhUgeKXwIE7UU3jZ
OBkRtrrkKsvStSKdTm5egvZp2RBvML8sNOzbzcwD61p6AMoXxOI0UccYBuBKPD66
DX7iwZbYCzd+4fFV8vH/8rOk3LFouxTeNQjyJq9gGjuvtrB7usIVdzJITF8Y92w4
EK6B9Z3UJHwQFuLIAhI6OMi7X6t67lkpG1n4JI9PA7KoRKSqwaEyVW6rtG2zHqSb
GnjLJBjuVKLglOMTUuM4kpO0k/dA2fOpGanapMV/xpK/YML60irTGrX3B0iif3lW
Ebb+x36IxmdY7qmcsQl902nMWhLDuv6VYKWNoiYBqG8swrBFF97m64OtxyVzaTXN
6202mRwygu+tH+LFmnQMh5pI2mgUEGCK+LGW2PxSUlWWsm2iq8UBWA671bv1ldqG
9GofAc23kxTd09coc4MlcxOUamHZcO+ZgcF1F0whowgbgKAwtuIIdlT7IAD8jS0U
RFtTP+xARyyTIielIR5fOJ+lWsshF0Farc9O7UXyWhe1JcKUyF2tnaY1uvL5zETO
iNhpe1K4YnxNeQVpsmIu+UiXm9zj/85TZURxuzdNvRvA0zvDpCwXf/clagUfl6D7
gNC2k3ytpvYZuL/PMcwNFoajtz2R02Vd1VcLBuCN4FdqD/w0cyXMFPjsEfYYYW1E
Jp5mMTpMwSj8YjUZT8BY/Fis9aIiar29+lczCbmxjJa/ZCnul2rk7iirVuuo3e04
PUqfES+gkbBpZXgRf1yqunhi7lr1LVBTORuGUSAEMBvEIwao82M9HaLpx5Z2EC3d
GGUFfhZvOzhxHSgfK3zH2w1TwobLgRj7dqI5T4598b4gpWp91bQb+bb50fxeDV4Z
PfTVUY9wR9PUyhgCXdgnuny+Jui1DZhPf5iRwHqqq2ec/qiLSDJ1MZGSQ5FS4OV1
jWIWancg2rqd+/0t2IBUWc5ObZEmdLMJj1N8BPlajox+7LiihQsNrw/+dGPt7WjZ
ZBjxhM994wBfsC6ov+Z4tWTOkvIvTfUAk2m9pLTWV1Dtn3sA+lO3vta3wAM7v19a
nC4Sr1Fpsaor8NDe3MdFqH6QErdZr3Wg/V6UV/w8E+haavZOaObCC4eyigJeOGK0
JTZKAQr2BHrTykLcwqVkMleMbwp8e5r06mvwNsPduqG/KkwjzCFyqA3eFbknDdJi
z8nd5++60AvIs/s3E0VoLkdKpHwTCqSV3koaF2TEmQBZ/uxuMEdjzygEE9WQoMG+
LKdNI3fvkVoi8jnqroy0GUpd2B5LxCRevnzSCXyuKpx2vVFCoxl74aFkOYH/7kfv
S/Z20MKqC+ommspz/FAJc//Zjn+zcXE4OLdEwH8Ar1VsE/HxbiW3c6g7fOB1kQqx
NEizRpNUZ2bzGbcJMmfQe+hKKJIWf072yamA2FUjIvMvGwXfnwgwBAmYSOgdGTOO
1rGsAVquZBv8UhZsIr7XW7r0eOMT+eNKG/AhncOB2IN+WIkdTsmVrP14mfKOeWzP
Dt0aO+RWZsbPpX6H78xDIwnFNsGmCCFs3NZV8+B07gfBgkb2QiEGPuxjpZBwbOLT
ryauLlHtUTTz79k9O9ydPgSpJHxSxn+M0BWS/o5eBuqdiG+Ua6J4U3L4ZgVZ5bU8
/TGbZ+Ha6XYsPLVMhACXYMTo+Gp/heH+KRop25SRh9m836sZ9d4F4CPPQgonekgk
rtFUTTL1g5IH7YtxqfSPLCQxDqQUveBCZWGZbIHcDyUGsM9n8OanVnlXg8GmjsRL
s/jARO9yKKJj1GOmazTuKzV6wr72nAl9WwLt/iVZEwcOugkO/vnQQwFZwmdn2WIh
kd9bTwNogsB/n6lvGCQwgAO+ebxLlbiDxXG9ciRurAVPA0XURquD3dG4LS+BrMLI
xUHHpQsHPQIUJksk2nuDXdF/xtJuPdfnput82pJstVMCnkypnI3QHgegy67zP8qR
dGwJHG8l1CwtvSOyB/PzJmhrQbCKDcOD8tyGZl+sspYK+mAGWlABbhGJhYaOhRI+
j5QKYavXPPSzp9ZD3cvTfjQSXGVHXffk2EefNkmVXYZVlfc8asEnpwDerW229Si2
upXbF52RX6vxCic7kr1FxwvyR8eLCewH1sfWCEvHS4C95riTSmYMUnSUqoCrz8Ix
av9n8j/xteo0fsEDkZ8tbv/S93NCAu7W2t838boud6EIGNN5X6DEzAs0EJTVvubZ
NVBvtyb3MixE+6tDb06o/pMyLU07vj2awHNdTHCjxmEQ1V1G/HECvPwxwhP0IVFN
VLkIwloTagUJmk1z3ze3LkpVmh/E03OrIL1YK86OKtO8ysdNk70PFf+7OMreDQqy
8+bXJHGcck43mD+u79AbFCOysONY4Te+p4g0fXYcU1JtB3fXqt6cftalJIt/o01v
w7ozH0VBTRkvTHY88GmwjdLfZz3ZgscBh6GpHdnKc92kgv7hzi9C/PvTqlyg+NmG
MANd8J6eB0Dh6InOvamgwngW/sWR3A0vAQ6kTobebeH3YE8z0Qts9RFg4fIsE7EK
4499/eaqbz1mnu8fFcGuweM8iIs3uS3csYCC2mb3SOXOGsXtLQxhebyqTAKr1dZp
daABd/4al2PsI9JgV5BftccOkc9XOXG9XGaZy/nGyzJUtz4H/gmeePt6HyXzV5fd
SusYi/QEF2tr1D9uStHpQqX5aUvVMtYa2aaHwTf34oR7OX/bdGFRzW2nMeS7J0dU
Dt5dLCLhH5ZaouhFoIgTB2KAsM+lIaO0yoBhyEIErQyp0z5A1sfygO5b3PqDBU1S
G4nBLMPFnVLLZQh+vmHs4wFg1nv5+D6xkgITzR4Uy4zwLn5H/IUOcN/6TheyjboX
YcMDvOQmKvyrEmaM8Xb8blMwneJ5BMDwv7fL6YYFd8s37dM3GAM/jIGaVedLtW2k
LsJDJPGH/RlbvPPFOfwt7+k9kdcMMZnBYTfei7sj/K+kvQmYqBRkHfOiuk1/J7Sv
/ENGyXNQl1uI+/HLo2whoF74botHDw96FKTU7EqgRWHA3s4OowFA2B438XsUahSv
PwYa23+JS/GTq4QsR3YlWMyDRXNJZce0tpKAVbQaoDNRMGvDh6nfv2TCeAPqRvBp
ATR9pg5hvCY8ol0Kw6fSVFBCCoax0xvJJgwFoNcccg3Z3B8sHGB4bRanuznD9MHv
Ko90W96B8eljP3nM2CPAOpc497g7Openo0Es+x2Msm2XLG4f9oXT57yzQAja1nw+
ZCQIQMznbFIJwkJLBYtAF8TY1cBfGRopZQ8NrOTNt3fZYWz+nO7Nm/VEhljwafEB
/70weh85Zr8tH1P3p4GoUEoTGRxCHmlTpybQrHMDsw2czvJmZVF23zgNPE9KRuWQ
n2qnm6UzEVfuMFrhN1Z0kEPX2TY/Rrofla5IKyZEMWq8748rtlhxmoc7jPVQ9Pit
NzQTCC5iwwDy6Bal5nUCwCnVORTUt191ezymGBkvf5ET6fNiOTjfPpUK9XztgwRW
1vV/SZLRCVN8iiXHTw5s4U18fluSAE9rAF6BfQoqBc1KyE6LRsy3LBP9tySJvIW2
xhWu12IV5OhC8Wxu/Pc/2oppAfSQREGWktU/W2Q/89JYDe2NwAtPQACVwW7HrO27
p8AafQrC/4BivgnIFYsgT1x+5HO4dROUIdhLXq9MVds6LJEvEw+bZ0k+V2OEvyVO
aw31jdP1jYxsEAwbvvbOxGo+Xc87ZlIoj1GEPzyUbhHzr7FU5jAeeOXaTj2smTBJ
HN79b6sPdJF5+X3/vKkmi/ov3aLW5CiW0HT4A4a/EH4kl7wz+triKOrqZOOqDGbf
aBRJ+aAvLehdan9IYlvzqVGctNpUxED4ncYua1BZ4MWC+3HtfTNGqFSyafaS+kVn
LObsQhwVSZmZo5UU/xNAp2HmUPJ+t39yuPyzWgdVTm5pKIo885lKRu4vifp5y0uy
C8JHP92BWJHJrYC76Z67CE5QE7sXOxCtUtzAxfuXPkEIjeCdkioUrTJjO3YEtoIN
CoCutmad4CSzUjl+55ydnhOVqNuSyXEd0hQ8+HNZ/s6cFY0Q1+1KSMPiRLZPeSKg
TqBWtV5Rd8MLyjz5bcjOw9tyYABYQ1EbnGBp4drNCvNvblAYTt493vQlQ8EOyu1U
ce8vIc4UqwJ4/khaaHv9FbG89D7oOj3qUOk2JRYCldjhbF4QbRKkKUDfnE1jQG4I
cRnht6kM6FVW4vX2TR6clrxP96QQhjKC7WlRkV8gpsdWmhXKrcsEoqEkGirr44hg
RXzlXzRi4NEH3NtN57v27TnV0Sf12ALft/DR8ovtDui5D4oX/cP2ya7O1VQqos/L
3Dak0q0ZNlH7uI097sKgpPpMU4qM5nK7Q1MC8oqaUP1hUJ3/reI8PzLwYAS7K0zd
qXr+eK1+iaBfIm9xeninTQ0mVgVtU/ifsV4eK1+ukuRNIj7DqPbZPAxh2TUhzD7c
yqRCez2wKvLeqvXXeUFA6SyJS2Hn5dyrnT4yWge3irGKcWK2yzd8GFo6lAvv23/G
Co541DZ9hI5gK4vwkoF/GIIwgnzPzdOXpyTT5S9/0psXfrbTjhvypgi58MzVDBDX
+6O/o/ckA+nzxrW4wF2HRF9HQIxsez2MeGg2cY+TEUS618E4KJQ+v1f9lNxxKuwa
/aWjmuVwz5RDk+Ycygl5B6f3kAhOlR0bcMW64mtJ8RHJR73hRVue5+XTU41VVQKg
jJu+pWh5HlOJnPwfdyCzF4tSfBeOA037LN/aLipgavjSNl7KHOvQLoXAQHGoIrVz
qi98Ag476SMZRoGPLJGqUB21m5Otpb4vRFZ5a7aF6A6ct7IQRxIZcyD525CecUx2
hcfAKYuthZ2u/voMUAnSRbdIVdzTEVC3K5A1lVim7DlxCI5d4xLlZIeWTdIGrK7G
5PJLAF9u1HAtaLkoh40CH7SBQvgIHUM3vrZArMFJbpSLyguztlsmf0m1JUDRYL3v
PVZSa3hx9qig7rzqI0YEG3p9aDcCx8hNNLyUv6Y8SnRfEWoz11/q9vfl1X17pbYp
JVXjcHd9zaY3ljJEySQa69u3XHmZextEv9LRfY8mpCCJCCYxP2reMYlfJjVoxcGF
LISP+WkTPL/ibncxqxAGi/Gq/nxWZA1riIFT9HvCu19EVLrQIpVmtB7WBtwtRYOj
Q/w39QT81lh4IqAs+yGtQ0GCjuM9ufBVbmB444y5hlYjNYymcoI+7IDt0NaJId7K
o5nwaQ4UaQidIdefK/uA6DJ7ZWqky5Qb1DluJqlu7HAXECXZiGocR90hdVggDSWt
wouKQAB/XBZ6Jj1CJR73kHO6ozk/OQVxbo454zuliWbpmFSPf+Z6lkEQMRXw+2fR
4rjl1tsSR5BTvKmZ3h40yweiDUGPFYjvggzR0L/3/Eq4MI0XNv1wQZjR4udIVupZ
bceBVvq0FZo6gzc9N9Qh3WOTZ8/jhpHfHImifQGt2KFFAT+PjlUnRRoz0B0Xwt3f
8UO8TTV/ZQd+lCwiIpZTDV8mOdEY5Si8DtY5nbsq3Bjc8/TXu8rQSFXZbdM6Hxw4
1+/WR/yFr2AutjCel/Chlm6cCqXrVt2qAIZ2aMMHI52aNoQ0HeZQwer4VK0NAGlE
twwkiO3V4LftuML5gqbDe3gtySY0y/YpCJ0rv9wz9w+FwCgVlk8dhmUS8/eW6wbH
3huSd3xHBJQzN3OZeKe2B0Wsphsw1mck11j+bW+odRI4VegbJ+LFn73sHQ4S+nPh
+BgjNaV0DDRdx2IAOfTUUlAoOTt5+KGdnesHtvH6+U0epq3DM3ga1ZuLhBZT9z8l
XuQckiTjtXzXq+Ub4AXUbeJCRrXoC5Fz4sfJDza5Us6Wqb7T0L6lq8xYZXVESI2I
LE3UZF72xWjVrQckXT75jZVE1GPRrl/ZpQvojq0OYYnqW8Hc5mznYBChC/fAlNkw
WLVzZ+L1JQOiYIwGsTaCd4yiuKM2QhoAurNya4q16Myku2XnhfCGzNPKAyswJjD6
qg0ZOFGTMwqC2WXerjscJcZO2472vEENEkW692h1TBpm3cV5H2BoV3NVx717S1d7
wHhxzp8Gy7LBxRanGlRH0cKW8Bl1n3ES/ttWEsfI7i6qfkq07eW45eSq/bM8vgva
8CUPmbHGtlxryScOgWHEDZALMMm4fu26z8nTkWU0vf06HYr7Q+MyVNfKGvO0aShO
/oqLyllK3ooYLPxmdPoHTsheig8UVr8RQ8MWf0UazpZeEWLFi2evONl0UhTGWHhO
Kdb+wnjCy/HbeyuG3L7YYlmXkOnrgFJr1szV3sS5KJ2Vl/TNTTViyCR3kGx/j9dJ
DOd+Sb/YgWBba4iMrKxe9apsziijkEdhyKb1xCSAfiaX/W6+CB25LcZqM34deZGQ
J4eRdzUsE1t5J/pr5qrF/YXompv9eBRlC6+2kRsbw41quxTuEkpucnYDacc4//Xi
xVvZCwxTxwrkz8X8LxYDvyY8mRF+6S6x/AKoCO1+qzPCwGryzAxR3jiJFgKkXPzw
1PCyi0jr9LmIcsBmz2Dj/wBTRPgeI1jOWyhGEgd/Znd+JV4O5GEuIpPo6wn7Bl4B
erIM4ZTsJ1Ho5rwqsjb4RY8+JTwJ/VdydcscYflCd1xvqbC+7oGaeIGrPcF2Nrmz
YMrv2tsraVRH5yZ1E7Wyp8qXNbfq0bKUEQunAM5m9KG4M3uEvdtnAqFrL4YeiUMt
KC3To/7sLkGUh97++TPPxQBWBiT6n07eSgH5V3Ii/OskVydHWModuUUU4Ys9YrqD
jFPPLhiv9u76HYiBf3tTaGrS9ujof8xxSJoEdBfqEt1n8KYXAs2lNNEqAhGF4MBU
MyJe6raMgaYTHEYgbjF5y7EZjWOCdUBxtpgPawNzGRwAEPr2C/8dLiovdFBfg+cq
KzeZ6v36+tn0F/F3TwcewDw9mtyDRvPNMLoALPrRh17s7hQQbQzLf6DyXy3NobsH
n81qYQBl4c+wyESgsDnJPO6L202lusitoualYB5TGP4nVstH0H0+yM1q5HhCc2z/
5HuaZE+pfiknjSo5fX1RN9o7QFC6Yi5/IuQhCoPXkcOdLVhsUx15ZNTrkc6AymKk
74YWCqvXDkIVQgjKQEyZfWLEkG71ua0542E3nMTJMR7nXeOHbrzbvmlVR9geJ/qJ
xKwVOUEnd3D9UvW1IVr4onvdGKhmcV6tTDcl/Pk4xZ9I1K6mZYhCWTFD+V6yR1qK
TjSuO+R+iIvU5ENsHEYUAp8+qBQgQjVip7SDN1nZmgP4DCqrwRzTZVWzoUVijuSL
mc5oKQJuEx4nkQMoZrc/fbV6+TT/5WfGGQJ8L8Vb3mZSi4iXkL546UwQLeRZIZ5D
xOgguPIZV/QD7/G0qUxTa1zsCpr1nFY2ENLZna7TZk8LxoggyCVAjPvsf7VURgqH
Lp+h4LaNKqFD6auX/CoLu9Yv9raerMex1Sa1Za4bZ59iZcnzxjHlPY13JAJXZtWU
WX++vmX+121hDfTpfyB4J/1nLE70q8T/McMsWNqdt8+e+sm3asv8ABdZIDeSkWOF
12RF2ns+52RYHI4wG/j7LrHO7f9f/g8b8jyVCA8lB7dax/Mx5HPmouH80YgvlgSj
bPIoMdkywrLDPR8jVpdj5FaQ6Cuo+a7Jx+f3i8gWWq9jozKbNT2q7SKH/2y41y1+
FjbhixmGSBCVx6Toyl03R+JKErcc8Bn3EuiIC4sf4SFnEi3Pq9VMKD/a+YjJzkX7
PakFFYFu4aA2yr7AJCVN1UJPYzSAdU/0XxCKaxabbr5tFBUgqGcvMJwk5j2r2Xoc
dN6+qJDFlLiUcRbVE7ZwmIlou/ahB9sqGsd/XCp3+W8TwP9HIsuyVZ24RfIeiabK
XW/ecQ83w3QKoWEmFT77HCP8Gs1HMfTWxGgQWpPclMPMmKBZ/oO3tnlGfsG54BWR
ziPkkaxAFkgrvi7uoKaGGznclSvN4d1GYB0EVwcMxcipkpv+S8wCA90SN8ZCPyNU
PWOi/2gpw7j3IRtmORlLf22Q1DPzzL8eqoo6uTOn/wBqoNXFxBlC7gEaYprgq37e
BB7rku/Kd7bBJ3I2EEoVfIUWXALRONGeMD4vnXtTZmgnxbwArQYMozps/OFQ/igy
8v8IWK6nyVqsF+a7LKPFNEt7b3aPlfz3nRpxkeKH0+Y5YIYKZPTMxIkOgJdT/zAe
f4JqsBv0+XNONtO1Vy9fEgwQmsFaYD8Vn0OU3Sc8InY3LdoyScNZ1KtmJVVKb4w1
C3qfq5Bf7JdW9XID5aIQag09hNN7dkRiURlzf+apkyBimEhWeUMfneOt8qRHxMbu
n5TJImGGkecToZRIxx6VoIGvWwWIiw8lhMDpvQ+/BqvVHmt+kO8j4s697i3uc3IE
+hrkUIxUy+WUwuQFKi3BVFeYSCNclVnG2Cp/s43pL5By6YG3mdeOAteMC3wwoaWZ
XnT/e+US7GOa0b4ea6Le/4wJX1dvpZQJj8xwKGDPerM7W2OMzALcLT079W6qIN1E
JWeywTiYoWaQzwIgJp0uAqeXTZk0uG4W28tkpjafy3/TwEdHkmGgUhhJNs6kUp4g
Ov/KeHy2LuN+9F0juO+EYApsHvmxk9FEw5UH3nqzRw/xJANzwRjVjo+pv6x96W4x
uplHR4OZaA+dg3pTJ2uBZFD+r/MnBLUJfFR/TZMFoKs0wdG23o0eEdiLw9aXEJhR
+tGRMD0RO/HlZz65LP3EER+COXvr2kFSBtGQxlfbnZ8bB5PDasiZ+yPvSYBPlIMP
4x1/StxSZzdWc6zxmTNZQlIl4pMi4YXBx7cNJnB6+rTbx3wKhjOLhwRftZjBhi6V
jQh2q/1n89dAGBqsMtPZ8yr8qxmW3gG+ILuPFH3mgrZXk7wHzoz/S8fx0YIb2fxv
nRbVVoFzlPY0lbWhva4a/INPIhZmDn9d/GM8y+LwFovL6yBUmYe1rPEu7xONHII1
c0nTSdlYMgP68wiyfsgRDW/cTiLPZ42iuff0WNjcV4pN0CThr3zS7Y8eGsFGIcti
HeiUlAPA0M+7uavlSZfpgNjI1x+Jhd+gBsyroDKzdOVDrYQr+CO5gPSJLnx0JmRE
rDpWeegL2dUNOyTPaXdyORKZBGau5x2iQFCamXSPhQnumg+aT7T5d0PUiWJLfnxT
Abbr6YWQwX9Wz3/JPK0tnrLYhE2Xw33n/vpAfmmolETwL8VeqivP9E1XLP4XApAU
JL2m+t2ZapPAj70hMqxUPwEbXpSxTEjhoFKckrH/QLjFpC23fL+yLGS+A5l+SDK/
VcS9zHgxg5ay71u672AMLTGNP8Oqtf0IK5hlXGDnQiN+dOwTFeEWkrD+T1RHbv9B
/QhEZ6ysAShz9+3OxZqgGdbzHN1gPawRpatjvu4O9J9uoq9GATPYdeFn6YRCmdyP
zP7X5aGiCgYyQufSSS/UBewjXdgo4OUDlEFTbe8+6WFqd18vogO9kbhzxYRVpbBe
u/Y49j747v43QY0GZZ800i4lcpbKrHLE1DikpmC6KNWviz23DzEkQoO0C1lMI6iX
QDYqT2STO6hztRLpoNbxI1jO8UkqRz6s79BI2ohwgXcNEgfoO8rxzjXMvOcWDb5J
LA+0sAyCkfDsWQ50tkc2GiWfYQfYvj6+1O6Rzge5SAXQpSAgKIBeEaldPgkomX7v
4qdxKcM2g3344nGLGyB0YXvGJ3GEQPdw7ARwDLS+KbT3Mw2Zelda1Vnh9XMRC2s9
iTkoRopCXfKzJGYOeOwnMwoIQge4U7dGn4zM7Kwnpsy8pL6Yta8X14S7nYSoPMg4
SrHZlr1BNAFGuVs8CG7xcW1KsVcC7CWvLW3S1MxWTbuQYGi7xA95TIf9QnYVRR32
jK7d+XQnR5j3dR4DcZDT9MEKjPn4NzOyyXqc3OMhcRguujZ2Q8pPZHoL2oS4oamp
db/m0VqOPsdZnVhlBza9v8R5PGVOQljWeWYG4l5l3qNdEfOFoFNCceWzKa63Y79i
vamyKGFEtCEkSA73Snxof7jS4zTu1QyfNXt77komd6FIXJFvV++s3+de4/s55Nda
v6alXlQ9MsR25yq05d9iTxT21UmgpAthOF/bW44/W/VLkqo7t34rCKucZnhdeEWM
tg1gBW6cfRIejqjf14swowCn1t4tUnn17QG0uqAN2NSdgeG8VXBmGWmlyclYIoed
hgiOvPw9VLCshYpc1Pn9EjNQZocxFOlNiCQFNpfSt9ysj3pJcssKAsU8E++34jfX
ty7m5Zlj3ODXIBEO9X4l5/avTlIkEkEWyN2DkDYbow4bxZaQESa0kM7TuyKHCtEc
+sTlNP8ejv/50wOBYRLRT5xtUXVjXdEtcaDWovMio9T0rOU6AeBkyvHEPiqW1Y1C
d7c6wyaanaV9CBkvE2zPlO0ZmfokKqo2fmWVJQHyFy/0vTCI+e8e3pYM5FeonoGb
qKeILHB2FA2FRia8TJdINYrhZo5cBk2980hxq9ZxvN1iMza7HrmnoARpfD3y9ni5
xn4+1Mkn/eGEgZURTEKfyIK5VfHCRD4I2rXyvvG0aH7CqvjM33rrujshC/0wnH/q
1GCEM/g3xw9ii6I5LEzh5jvLU8pvNxk3AdnnQ5rGRnyV5O4eu8irg6u8QRhRgAt9
K8rKIZ9k4HhgqLVJVuVVLaY/33KUKhhnDPM3ao1tDlC4LLvNrtk9ifRFgZHEbbCr
uVzFhq5Zrdgk03TVBgKmH6MxqB6Bhtn0oVzd6ti2CPfXTnt9WaAAKpYw7145TusO
H1Q2AMlQ0wnZjpfdU4dlILv1DwCxKm26NwupYtjUHqklb/5HbP9h6K5rqB4pbpV4
QXzwQQHJGhTwt0zuLSDBisiROsROIKn+agc9StvQY/u5oHQsYAbqCfululZMVDJR
PwGfB4m7HnDue8C28YIZunlab6R2nZwZ3qk0OzidOmd3oHxiWfPW9GXOsdvKHTY4
3u6JVt9va2MAO1p83djlSPt+EgP4yoGC+HryYpIkDaScdiyFIBKPCn21/jDOjX1H
tncQ4TdFuoxZ9RsCBRvJQD716DWKqvwwaECD/rTrHwRSCFsWCyzHJCRaoH5axtH5
syeGEyqd5VFFhs0BXTuSGS88ebhsCQLroxcnx2bJqafwXoQ03MVhr5rDo+EcIiSS
HI6O0jVEtEX7CmXCQmr7HLXMX6MpxmNj2JLdrlTIqgwlJcaB3aDywgJuHyZWgOkG
cs2Wm7UaYQ68JvIGYDAIQSHXVG6XorKAZVNOB495U6zKkDf44Miuxj/uQQbdPFOd
X7NINv4uZiVu0T0OMjgh06oP8rEto/KxmRtWGLyhZVD+RGUXrwDBDN9j6aIMX9e1
I89KnVomZRzvVYrny4riWNugxtKt/15g/w/91ldpS7wu7CBzR9f48MjCG242IvcE
YDDcnPHZhwrTupeKbL988kscCNgdYyxSL02Q2RboueofhFbURgpk1oPEfGc2DaeW
RBA/Hgt65xFXF9F77/CUgVLd5wA7KPrUxSyS48nKAe9xqn5pxey1TwVfOEyST3Gy
oGOuK/ZN5YYRB+bjqZFplOMODUAr+8GAdrNrrWog1BSq4tFxd7JEO3lbmQuKGNDE
tC67hjsEEQCn/DCY/9jdZFMcLy4pI8b+GtfkW+DAfARyajVAiS2s8+Y4emU4EWc8
AZLstXhy2tv6Ls2C6Bsl0Vb2cnqLZ0wnpCFwNm7ihQCR3L+rnYrDQ3hWxs/idNEN
RjTyyKQRvozrCDyn8lvj9zbEZFbGomq/+5rgPLwBFb80R5hAQ3zhLDxlftlpDEkv
4IVyh2foZr95sb+5iazU0vgUzUgXGLQulZaat0Pon3o1VKoAKIDGB/0BcFB4aYJl
N2eCeAgb3eo07RXhR4bwHugnoxDjJkWtD7ITnwkgMoYpSGm5dtyXVTkI0Oup/f4u
rzgYx4FYxxjTZAW6To/PVR2rFZPQBob8uVoXIbMcZdKGCs7WKvXM38dm28GuUetM
bZOhrxuKGeVamRv285ahgZzC7Ccd6pGooKnSVilUe/jKyS4JgS1Wn/XTgZzzlWzr
mvxaoZkGaYPtlvwNJT+sew+fbZdgsc8WfhMHUYW5CLHGnV9/OyuFrlQstp+noLT4
Ko1T6it8h7sXorfmtOGwjf2xx42E/xlM0a2axjpORBQCE3kRZqy2iVv3CFTowZDd
aWP0cT1qcAHIkBjNIQwoP+1yZ7wgvhATwXHEKTtKFYa+8K4Pc4iLkrjcPQhhcIEN
d83Vax8C0rlLYCKMRim38+9DYJ2pR9cGUgUBCnOP2gqWqna7JkMY/Tq4m3rYAjTM
D4VyjgVaKwvw7Z0fL/p+ZbzcDwvEsd3wQtgB7sMXeck9++rIV8O8iFdDN6EL1DwF
Eoi4Fo/mlb8pPtK67YBx3nR7vK6CpxG7Kti34jCdXyyLfkDxfAA8hschGk0x7+VY
M39WAWQkW5HAaVl/a+BklG7DlzUzUOgnCcJxZIgFGxUq6xZzLjJYgxu7JLCF/cxG
SYhoEY/CS0BBPkNLpZhuZinZ9w0F7AHoH24nJB4i6i2L0Y/R3HaqHObuBULy8SDR
AFicoOP1Nso06lz4tlY/z17kJYFjmEltdSnJysOwl6MZu4+Vjp+Kx8vewIREj4er
t76d/Fl87ILBqbCgqyxQ0zb7t+mGG7kc2dFIAKsjZj4F9seEvpLNCgV3GGiThMWp
E0birWvoRcXF988PQMstNx2NAs+0u/UqJ6hw0kc5fDjjXg7uKvR3O6CvCYEkQluo
XqgNoWJc3zTzLBe65IirJLYhP5mspZ81cPGFZxBId1AuPaccDoYoPTjDL2zwef5w
YkEGTxoHtaIB0RmNHNOUWP4OP2zxjyjQwlx7OZB4tjq6OAz0FGxnSOKXQcQsivp1
RaEjz8wJrd+wNNNEY3vMRUWzMjYXGfsUrw0eUVZ9yFvshIJsDJTQKlUIKoDZbf0t
MNvfY+aE81QerPp8KeHh9opDtGWQOCmXAuWt+vZ2x5swg4n8ALwigT4qui7wg2hK
qImfQMb8uQf/SpTUuV1hKCVFHvQro1HamFG/3P72bXC0jyQU8mfmaPH0pX5Yh0og
Wj1Jr1P+8Oyw/lEBLNoYZWLlnq28CFFQo3ylstgudCLXSA6BvBuZbDxToZyreFC4
4krp5PRA4ETPByrfMYozyWYGr5PDc4PknmokX7NdKENY8f/PACG2t4GXjLEv3gZ8
/evOK9v9/4xUKVUeFIZgjJj2/9npRkz2neaR0cQIqaMkInHwIWyjJzSiWCWhpHbm
QbfRyfn6DJo/Zpm632q62GwuQDGjJsvGAQXIxyJV/5sGqLX0Kk9FZNEKSk+Bdxlr
OhvE+UzLVWBPrQkdw6e8mK312Gzu8bBiNt+G60+ZM/NHiO2H8QvReHi7L+zQrOcR
yEJl3YJSBeDkaYZghHSqLpvz0y3J8yQ7qh16/EMG/VCfTsIoD6cG5C5x1IF8U77q
XulX4ov7YfQPJR0IoZJfXbftBGe+uGHQk5QMeRqGyHodPOK2ibWWlMDMOnGHsTnK
3z7W//Na6rrotMeKKRUnbeY3UdvwwzRqiLD8s9RUKtBFMRHKJ9gmY9hkaBxocsSb
gpOpTiBp80IS5PM7nfnhMbZ0Cz6BpfKev9Xowgm5g2wxgosNFt07cBLZsENKtSKQ
U4UA8kvdi2YnOS26qrLZSVde7x8yUOxQ7ISKIqHoiXx3GYGsIpebBYJcoeF5nZwx
wiJ4QFlc5ejvhs2VkNygj7TmB+x4xqYIzdihzKAHX4SLU8P7aD3IYuYKnhSNiIRR
Jl1kWWCT51D3GKPh2Jz9pG7SAmrTQ7qHHwsi5ewtP70vvF/lZBlItrfjRyALZNVy
O1WBJ4T2gebrN8saMKY2pgvQnMgM19HRzJJLneHKO5KkLgtPnxGp8rYGYk3sd3T4
hC8Ovafsgm6jVstQLB2Ink0ADUceDYvjs3eA0rrLuzK+1vbX8/FfXlBdO5EMm/ma
L6bTEWNbE9648YOery2+310fuGN7Zx4URglT0r9vJltG8Ts/04kwS5cGn/GCyoYO
kolRSubl66kn3Rd6gBitV6TBR6PrJqNd/EqZ8mOaiTuKSlHxUZu+ZxoJd6FEFcFw
nHlNG3RgpPhdk/jUpVnezTm8z29JahQeUE5hoEv+DH5+KZ+mlmSJiVSD0j4eqF0p
Vyh60C58eQkr7l/k7UA9feH1vNLcVGSsL93QIkm8AlDW8VK5nwUL7y4BYj+3fYrR
AwAUjT99TMuZD7TbhJWDHDHlzBQ8qfIf5lXHXPaLGAhXPeJqs/NEcLY2MyHGW4HR
mQGK5tXmrdUp+j+8AdFdaU49Z7m0tTQE/2VlH4hi2DXuCLg7LzkuiHW0Nd5T4Pge
JsYL2HBY17HnUcUm5PVQO/o7eibpZbTtco1Z3IwV8BgO9KNKMBye4STCwv6ZqO5d
zRYGyPohSPiJKgUGK39x9yikVogaZ8pBGVZVVjkmAv+LVKDNgD8WUrsNCrnvCGL/
57NoQckUMuaCf2QXhV0ipJfXJWJ177FNdjmKxkopQ139LH2efIkS89AWdJEFeggZ
lRCqcDV9/2ekaw3sucR7Gakr4GTr+V51SZWDdHTjmZu8E5yBccDEN53vZ1XYN89w
3QGKAxOge+LeJP6wXPauTexAU9NMurBlmeG3hJyKU0IAplPOfILuVvBSO31M5VOv
K3K8FY7rNqEPE6zC8Ybvo4d4rqZZ21J3O66MLC6cga1git+Iyglvs2aLRoM1J5Cf
kbtmB6yVcP1w4wv8mUIrZe8Z6aXKBV6tPMhp3e9DKTZIAQrXwfHcps61hWESmc/I
yAQ8OGB8m2uVCumCebZeffvuv1J94wMvvabf4oSlvfb9ESJVRK0mlF2Fp1quHAQJ
FKlKbTNHaYQqf//K9sM/pVS/JPZRBg6F6Fle9pOZ2VNIv4HnTTSf9ihbPmRHIv8F
1IDZE4JZz8E+Kg26Mt8Ddb7OlyCEwg9//Vgab+2ZRSF0sw1vDTcd6rnyvUxcidRJ
NiGvK7c1u8G+joX1ceYnf96cLh/eHTheMwPIVom8Cz/OC2blXJHy8HbQ7QkUl5hh
CCP6eppmuAxOMTN0YcFJXmbZPMqNQFHdXAjIkJhvD+nvoZwcTeafTQDXbjMy6jrL
eOLbPbGCES9bQq3YlZilvaKtZL6QVy9CRdwQNlDv+1hY6kHZ5hEnkEgyhRu4pXno
cuWwiuXHJGkSyNgTQEQRoJKEmTdx8qNyRCy2OTs9CcEP1DTAZxsDfCoIM0+umobW
DRlLlBQE/HMyrhoqM9I+BEpk+Qk6wKrVN9+l5CbpldyQYrq/TlZnYdxEokqABFnc
QyUCzL+FaZR1822KkGZRPlDNlA0UhoNeTuODdjfzmwGBIWIPumkPdBkpVogFL0Ge
uvDUv6A+oMzQKER8F3y27yUD8Y5NJgpAvDaecj/LPnUAnXJ0Mutqb14djUcN7Z26
a+EoyW0BaVqTTruU3nqgZ9Fi5vMXKNbbknvS+lk0667MwQdiCEdPJq4FPY+RH7p2
V5rY+VDUIOx8V0ek9fzS3rsniSvsXxmt52xlCgHSLliMcKf6xcDt4wu8XG1ZyFJV
7iUQQg8+Zi8qFvC3RPRETPr5r8CvCMYymIA42c9EzRSgtcS7owaP1wzWtuYDXUMB
mtno7CNJeL5O0tnN+nZtdm3aXYeZVNZqgpcpHBjOdLYsc1z29LJ9Wj/T3EAr0eyI
Cg8mQNTD2tbdAz8eWOaGn5ODIdS30eaKTYi6Y15LT/DpgLqJe9YAA3mVA+7OON41
xqTWDh/x4+XcZ00BDgFQ20302sJwWrO5+n4IAsD+/Odp4sQTJSZQEkFEhHzBDIpE
xbkJexFPOA/RLYJaX4gUylMBz7DtM2a7wq0HLQNb73IqJW3y77lIS4sutfaYVc7c
v6r5um++7ckNjcYO+en+rUgzYQoXuSGg3bzSk4u5QzF9y2T8GPeDx38OaKSZQsN2
lJVY5pdCz7oVa9Xz/DyKcAym3WcRLezAkLaPUVn+V/uAN+QmMG/Qa2B7mVG2g+Be
D2fdkJdx6ameS5YimUf54yAgWuWkzo+3REKYrLH7c4oPrxaVTSo1RXL0yb96iwJe
dxy6vIqlBD/46RlX7zEhkqlogOeQ+dDPq5TerJqlShsRRC8+PCESD1K9sGebVW4R
c+Uq5ZzO4z8507YAs5wuLQpJZWMb14XMzpfWozZyvZJ6O2mAlnDtJeIMmAdg8jyc
Ltle05rX0P1ecueu4k+pLURhCN6Ps6nEa4qYvfVxpl5mN+kjOxZ3q5lqD0Pwrole
Ui+HJcArIBAOGFYb9eGUe/aKJnu+yk3txvhGJQBSyctLFlBdwOUXJHDdmRQsThCC
5rvkctkn+AVg9QJXjqh4baz2tpXpm9hz1TLwKlxlHcojIZX+o4W1jQqPMGYuQ+Uf
E6CQE4veAz3KrS8CLcuPgy+z1P19E/t0LUe03q8NIRkLVqY/o9y8MddU5er1aHfL
emShjl3Zpm6vEAe+dxoArBa4rrg8XTmKYAubewNMj68xUhgw0bj77bO9UI5U/jlk
mkZ5PSEoqoXNKjRUKCCxRThS/XpT1Y5Lg4DRV545fRdHejScurYT+YleyqiNad6/
1a5Fxs2sRqWiOww3OvgS/ny6TA2nXYQklxjeocQJpekuOynaJFk9s8wQYY02JWTX
B4yIFL28Tz96COLWtPRKFkC3SgGtvxmHJIuDeNYzhbS0t+yz8SQfZNQNxdxgD6GO
3/udD6GFpmGWXzsPpY1ghlUK9sBCewGvc6T2pZWkBPmWTZg0nt5NYHXabuz9DqkP
9cmT1JfdnaRhoNPq4VIgLRQq641j+lK9PB1F1QEyn4nqTF4lesskdnrF6JEmqdL5
5ChWu1X/iLzwXSVZ2eZAQZzC9UaHYJAjaj9wIZ4QLzW6Tc81YZwweKGMgFNqdnGo
wOrk74QAAsWfnfHSNRNKPwvsBywmuRyV3MEohqCyx39SHNt015QyG2GFLhdFyc07
fS49UkM4gwEv5VxtcuN4fT1dMNSSo2zAR+gF3C1JYneHe/EZ4ODKvImT+bAjZz9J
ULJdBr9fuC/BKLpAE9iif5qvf9CaetiysiIBnkTqeT0Eh+zgsB01Eo8eps1HHWe2
9itJtJgysoB5dCtHlJlJSkSLszRrD9xu8l6SiqLxcVgfCeBxn9rSAja9V3/7C1W7
u8OmKfZcztkHRmNPgqSZBKwFv54hwLGBcISXMfhJdE0yXcOJ8z6iDEVNMRGOHYUE
Rpj5SpbYfdIkmDZj1hQ0Urn8xTPxXSLZl63ldefu+LkOFrFQKVmZRHU9mG1HjoM0
iMWwmx/UoKygJHxEwBTKBfDpVkdsZ4cllZ3EBZji8Usb2IeHP2QlI0TJVWCBgumk
3yleX/K9+Uf1tMtw10qlVnHRMVxRtFAGwIUbixdUABz+7YGGzEPLfZWDAbXuNMhk
dIfukSFnMRrnVUUXOA3m2ctjyATsb/c3yFjSrR3gMyNu/BmqS6yx8XU1ooRuGFpM
jFdC4Q1c1rj1aziPdRpQO+iQAZyt7//s3Irr+Ay0KwiS5E1MM1+f5iG2/5GpnZbk
JvNvJ1vPgfXY8m35FhsmTRiWawSZxEDJ5TaB5ddI33xmGEDWQJsHh57PXysaseb0
qWspSeQ9PgRtTJhOZZySlNtd6QybKtW+mG5ohhGUxAMAaeYzMdXvpNyHqRvWuL7l
sMRlhxF1S/pLhfQ/JHuZfutAFkSuZRVfVEUA8bCkYoXH+tWOPWZ3qvhyCGN4sNN3
/Ba/beNIbRcd3C6jCI629wQFfMAAh/S95fZMMZR9DlSyBBQRWk3Op6HtZjuRJAO2
CyHi7eMqeJ4haDNYBG1y2oyV1j0MeF5ydTCUU6xbIwp74SigfalDp3yXBWGj1Aeu
qsvOskjveVYWfKjY7uiR6IyjmTjcGAh1wGvD18l3JI30vJv8OlX0pAfKcBp1+8lc
LNGBsqIOjp+LgLtnjF9Zpq+g0B32/JfQHj6gndDCuxh4IlRWZTXRPfB5yILORLCf
1t547dahgQbjPSnFzXLDnebiHXJqoHXFwG5usSbYfIHYmsFQNT+h3hF1EHlTDKcC
fNa+dcsJcZq8g4+j+qqcXRsQFzThOyAxaGKEXr+kixAssvLFklYC+ph/YAemURGW
apQ3IpD6ejwxdBK6Cw0aXo4GXbWneMLi5eD58P49WJT31T7mmFThujNolEfBqr8Z
QzOMs6IWIoyjqU/EOOBE7Od05Wk6b8A+T+2Huz1mzaZGQPzVTB4ZUgArSph1zM7/
1VQZnj4sfjcagMEIhcSCABxA0QDj07rS4D1/7av4D+bGz7wIlInIiG2K1LqgSGBP
1MYQUbstuqzjjbOTB/TAlxOCN53cjJAEcFyJHkpa5FLiECdq9h5Vdru+m71igGjj
kIAZyki8bxOeFi9UoNY8uHXv3bRK9/jYO7PVv57cdlFefUeh0Pjb0qH7itdC0Ygw
Lc0CbD7F8dW/JZV1zqtWqxWWJY/KCZNbJIdBHh2ZmbIV2pdqyVu6nYIyrMYcA1v7
5uIglP6JticvNh/7G9aKh191P/+m5buPflLt2MEtLbJ3G+WKgx6RQQiTbO3WZwTg
GLszCT5IeS8a/J7MWu8VaILuzH+YB4OmavHgzA6HPhLZ79dvewtwSRliuNM1HGjR
gGXqyd5v6PtKTAAEhLXZCXTiI35Zle7T4kNTEIMewzIObFK6b0+DDw/ZyI19wWgv
g7djiUMIPCG0wna0kBxP9YxWgWNb7HsOXb6e+JHI/j9QR1ssL3ULIQyDBi9urW81
ObrnCtz54Tln+8E1sxf2dEDZm6X1CnUV+wiiE+dCH0VcK9RxxrCD9HXnYkuVtrcF
/Zb1Aw/r3l+DMh3EvTxjuCQyLH3S3fZCmi+VvfwiNWrH7SAtKCmZj0L1XKWwGA7o
6OXNVmRjrwo3C2sACHGucmEVceVomL5taKCg+KqQoqoBkX+2qTj51UJBE3X/kuo1
6VmWJDEfwsxk5kqwfqfbCUAq/y0ehSC9GCrNwYG0zQd5zyBpCcsQD8t1ACxEceQ2
aW3CuPv5G0UhMEXsA1gTne7OYyeUeCXEtvkF8CnzZg06YJ2PBPQXr6cDQqTF86H0
IngzSBQCTOgZxRmDQC1Ql6h0xEkeL57Zcngn2kDQo0HWwdfhhSnpIIFWk+bPfNMp
lAvatwMrbxWJEd+/vXf0LbjWieqpdnCjQpeDsBCqnr8Xlgg8dGIrizRKZZEBzev3
NiCJScDlwVBT9u/3H6lChG/rDfhlxOxGkOeYWVrGN4w/ilW/sujcH0jfJOmmnb1O
cm3fp2GijJcn+Lxb5MhsNMN+wBUx39O4ybxKH027LSpwZt65d+Ovl3TIH7JgJlGz
fppov8d7r0lSetV8rLttg6y0ByyRCdIOmPXpsiL7CdnLcVskMPvxDmvAzSqvOHbY
rLiwldx1egIAua+bHxuSGcoJoFFsnDyOGUfdVIqBerbPryFEGrjlUlV18Ln8JvaD
PmaC/LnNggPyT9WVvZOB8flwWR8oj9HYLWU7TlrtEb65b0QnkWyHSNN/uW3m/wLK
VvUgyM+0n8BJoOrFQa6WoHNVV1kPlrTCVZLG46KPFaCT8VHuBa70kn3Yq8qaHLAi
7wgFf1wjzaItVyWvQK7OOYrAYtviQSrZhcm92Xzyo6sYjYzDMA/jPAr2T/dQ4r5Q
wkSp4TpjU8x2RIC2wiiFtdhZTUKYzan5SeUUcl0jAtL9arOfTxy9iNvC09i3gTfq
gz53wPKgTnB+L6iZlvL+4F+fMRaw5hFjVJi2mik5PvBqm2EEl0Y91gkGjq0TE9MH
ifg970mdOa+SlNuUNPhY/fdzW5eaOAB8u6qw6tbVWxR0T0il6RvmySG22Fz1E7sY
4NF/+o6WiOgCA+dRF+fXE42r/7OknqlUF4Ki1Wu01XaNV9qarIa1908j7VVRTHso
MK0kn4XH2rRZYbpsSUmfLSiM1UCXxy+qw08DMDj3aogrTDjf2JNZHl3SBHSBzGIW
/W5ZW8IQbyjw/cAoM8/q2fEOBWQvAn0rlpgJrrEqqwtukX0Xe3u6qzfqnQWmq7Y9
eaMiRxb5Q4NM0JUhsNlEbLsUgQKBxJWeSIMn5JVTleNgZ5XhPe7m2qDIIvtQm3tc
NdX/3gncQnXGyDzIeFJ5ILYOHIZGwLXw9kLVM4SFY+mpFw9Wuf69lZkp/wjfSLVY
Dgv6a3e22sHmlVB9sDX3mBtVz4sztUf+NnQr/qcKNRUrHFAb5fqe7Y4aTz0AqOyb
bS9FUlcpZ73X12Rjmd2L6X7LDhIgNp+ZUVDut5w3nnGsDbj5WBMQfBqZRunwZXvd
PwMUd+USA/Y6gVHC2welw1x62MJN2bl+3hIKDDbA/Sw6lQz7TZNuL6iJHWjWQwH0
x/uxaIj8D1TTLZRhatxUBEJMfb9Lp8q4uJUTR4qnNO2vEXOOnb2kg/FZ7SsSSfOz
z6Eeas7ccsSrg+Zv/cnF1bH9NQcJhNvT90RoG6ZtahBGoXLw36DIoWyGlntWO1DC
iDz+ZgmInoVCzacEBLk/bHsKNVlzib8+7XdHjA0wwMouA/tn+GnIpRp/oEEi1MOo
7NC7AiRStlzsqZF+lvU0ap0T8rj6b7/oTTE/tA11cdvBOHndRoVaYO+6Nru9rnmp
ojCuGW4biS8Y347xSnq7pL7z0H8zdXUe1x9g4hIdogaS9lQtuH9RQ9hdTIfJZkZn
JnKCRMzYzX/XNI2PI+E0RjjQiczRsMrWNiUei7Czrlf9BycnnD5ZvFhqigXnj7F5
TjayyY6WOO8qXAxWhstqetMjuwSLVc2UEvqyFKW5hJdbtzZikMERTcdcQRaZmxi9
smjaX5e9Kj+Y4utLgh/GIfFlrjOB6YZI9AvqBBbpmmmlfPOlPr2e0Wn6oB6BoNYP
2F+h7T0eSqWv9R3mhQRFTLUAoWAwuxZKcHp93x1+4QKRbx0C7bFGZXwU60HIEcYB
u3MvEjwuiNOwNP1x9Cvx2JHIg0wseVbMFotbrd2Csu8wJzYxRDodmIv56vls68/v
H+fYrv/uu5Gj5AyaZT4YT3KLgSuY8DEmsRJdeHKrikUawJfM1q6X31oLbPYsEFpU
4f/TE0k59sab5qWN7WnyNZ3AP7DY2kd6p4aR0hx9Dbzev9FUp7anhYbkAcSiMV7p
qRNKsWTqXHBBC3dqqUqej4XLglmcIRf71CRhj3Wpv6bSHuCw7xtYsn/1Aip3C7/c
C794/Bd6BcJHImBqYubuSJCE1igFy9VMyG0aKG1d/mxg8nLQXOhhFzJU01OGxKn7
skLTU+zU3b3MO7S5aAtDsDvSexeukfUtPQ2OOlwmr7wcYwG/YNipuLMdY9EEY1+Y
aOJwbnb7WliSAmKONhbkhPJlsLpYbvQRuWGI07SI7jmV8ALRSNrKwtmT94b63EvL
iceaZ0GYRH8k6CKclO+me+AurgGy+uq0zgONoKZf/HoUrP8B1JONDdbtHoVzxxhZ
KkIBSGp8NYr/EKbESi7GwJhhlcCg3F1c3gLxLtvh1Qfp4NA/cAw2TtjR1U6C4nS7
t84P99qFbAXBpTvoAS3UV2izEUW7q1OGIbDH4RVBfEssTzTA3iWeXGHEJSUo3NkP
O6zFrQMdVml9nWsxXtVl90HE5DdH7o9qlepZxIhvXJlsLnrPjRgkOpiWQouLO9zz
tIuTo9YvW/zKk7069tx3LaGZB6vY8KwX45x9rsTXghEHNRLGIPBIvhIFYCpAeBSB
3nzsFKibNu5KDxw16v1uTEaH2Knt4XdDUwT+UEYKlSzCb6yvqlW41hHk4+UENv4Z
oIPIM4GqQyNgNpIc595Bromfb6a6Bvo7P1cLU6TrM4YPWSEELvv3mFMDqBKmFOhR
S2qGzefEqgjw7Ph6Lqy+R1oPXdPaLLilsQwmfTsaBfzWkL8HbuzakRgWDtC7Q7Bp
bQoeN5Jz9ZAdwGy31UVyrkeu2J8jMfS6/aEVGtWGTqlBYhZ5qC9e/teicRRh8qFf
unM6wXbo1LcJIRihCe8wsT9Hb5+L0Ke3W3pypAol8bxOGbyTjP5awx0cA5aPGjlt
4CPxRe1RJb2/QFIVZtwcx/DxB4tCdsrRr97Ja7yjbkTR2Fn9VeCr925uIJzmo6DQ
iKWpYv2xoSUFpvMxbuBE80tV8qgU1uAk35pVQUdFELNHCtiVFugWrI7S/qDkRS2a
aT0uJEM/LJhCULUCci7L9pT+3wjSMy09KpnpAWNHAzIXPTiwK7YyYYpjYB39oyKx
9AZcr+mVWIe/yRJppwwfuv5nh4hN/Ot608Ecqgf3JgDHS8XB1v5jkTK7urXbbldI
ltghghvCdyUGw20YwgNKl43o1Ut/TDK6mWslqZTs48UcrpJ6OQF0iYBCxPg219/V
tRUKZ+sP9Jnj2+GxjgNvlGJ+C0Ns3okwztxHxipp1jOatOlm5nqKYMzoQddiGNVl
qo69rkm1PTO96Rrj742hTx2yHldFzpXie3fWBQPJGES0gMXM7wwhXg1FwvfMbhHa
kRhc8DiooXf/JFvMdgXinYAQq0suwEgHSpt3DDLDqPzQGhTNrTaJtQfsKvdk/CsA
3k2NcgtpnkQwWu+mxC3aSpzyMAtVu3vWIugei6iRGDUvBGJAyoKvc+fDFPAZxJ52
/iym8FgEhGii164ZG9Rje3GcJALpKiLza6ciWYidgx0O0f0GbxoCX5+LsgZkICRL
nwXtdqMCutw5vO9Kp2bw3dQofFwrYRZzhBm5xZXU8xyLkL2AkAIJyygue7pA++Hq
mCHoxxqM+AaY8/756CvArEaz6IJan6cPURYy87+jleU8dXh7Xncn57l8YqeGizPc
PTFEdIGcAz1b5Zbdn8rwdSJN+CutHPQCGXxjBxPAKcRkTgTry4nazp1+AwQdOnAU
L4+eh+ko9+WvJfNJBAcEKqi4p/S7j75Ska0i7wKLDiBjgkBbgd5jec8Uno8goE7g
VGUO2HqLD860VGAuTFNct1y1g3PTFfBLPzzNP55JQM0pEMf68luwpYNNCURH+bDN
L4laxNztzyKSUdeFXMbh2VdYm9RxNEIp34xuFzZz+QPudz5rse9RIzsWvPmyrwQm
543hzM2NWDEFQVeY18/xjIiJ5W19WDp0naDiyQGVW6jusr5eTAZd92t5DB//9rKb
jSsixqsMEZ1gT71Crk/n+NBpG/wMhIn6fHJHfQeMovPTwF3uxOZkOKijtJ9KLzHE
6I+re4RPJk68Pye7gsz4SrmUJJef+jWwvN7fQ0TKUa1MYBsY3N239XlnUMK/2q9a
U6VW5hIKnc7yh2bdoD8a6Bttvs8kXGyQztNxoC/hfIxq0vYRMhFOrByn0Oc0dt33
zosAd8SYQ27I82dRSwDG+NlPzH0rd1iizDeie+g06N4ipk/3ESuZImxA5wTb/EtK
C1xM4SaESYj8Ej3z3ZEx5n0+7XAiS9MGD9vHFQl/ysmQQxSqWboysxxhN6rvoAsI
w3YPUmVhVCrwqW11Sb3icJ/qsb71wbPznIZmPeeXtW5qkStPr6G1QuE7xJgGCVDU
NVl9k98eniu7eTY0ye8F9v3MM+UjWpAojUv/kOxtpbxZCm9aMEMLoVAxaMnbJ0mc
kuZVpphai0czpWevcDfz/xw2O4d3Ld6WnXl97ruvnWhRaVd9XZFhHjL0lYb/x8Az
XkddIOgqtdFIcWNtiOtm8rQIeh9Ac7euHfWkfQKk93tg3mWTiVE5DusYFREktLVf
gBKKLtE8iRzVKQXQW0AjFviJ0rGSaiV3PmM6z7SJHLBvFviRnhdx5Gp9t25EO393
XDlKYr5npgLZoy7aLmwbobWFRmbDlkNz1ou3+9JUtzsOurj54i13aMzqNUQzHZjp
HvDNai7bUcoHEBAswFWIgHeHSbIb60pROXxFB8VRXi4FAPJInaYnD5c5zr3JDpOn
mBm7lDOta44RR/na0oB2Jg13066kM4hSPqP+jtO0yG+SznGa8DQVFEkACxD+kASN
s22gxK1jpOXiO9RFPXfMPjd7cAffUKtr97MNxZQne+Oz+7M8X9DJyaTRB6XdAeQZ
8zyi97Du4MjBdlZAkmr+Mzfey9n1zUevnj/APcdT18OhZXALdvPtVV0TH/IGqy6o
lO9R5dbDKXQORaEGJiob3ROQpSsdv5FnrfbhRUxGpwOG3ZuLR37YZU7wMEwyJkWf
5sCs4tJP9UveCiNOObXSXa2i9jFYhs65aeETzPMljRFuP3Ea+XsSDnGXymzm56i0
2obxSj9bKE5o4xEvJ9D7UTXmIzk6M8g6qR7IQKJtI7gBt+AGpAs0Yi8PLda9zTkP
I8FQBXMrPvzp632lPpFGFEEwIbsdJKBWzjC5EmJc0m7Gw6vgT7yl3FQF+iEqA5nu
EzBfAqqRQq+MQ1ADwkCXnWcQOLbuPo9ZCX+4VKc0hNfbqkZM6lzU5T0hxyGzA1DF
Lh58XYf7A8TDGIaMy3/fYcmv9XC8GV+he+pX8MJrUuKtF+1DhvOFOz1z97QuDy1c
LXJXkk7MD7DgI8M/9Q26fHuz+4L6Sr/Mzg0jhcnnC0OVvlfjldqUXndKUJH6A2QS
YExrT/HZggUtgmfpCJLGSFy57oGlIdUCwpxW2r9wgRiho0NOlPFP/Yj9RLIyXC5J
yqHMCOieasPKuW09maYDqzHGu0sI0w6wgOVwSkvGB0VG4rnwSMoOzBfge5Ew0HxX
5uqPhS42UA8uih15pClZL/5Mv6hLgIrYFUJU7y6PUgShbQRQa2IRuz95Cu43swqy
xnyX635B82d1U0yEsemiybw1ZqIjRLtIjchpm1XHJOtfUtBPz/V1ar3/u1Qs5AFw
eijyZt3GJnNaCvkowZ4czU7iBH5pPlXh8u/m3MsHGE8dypJvexip4wTZsSqgitlm
4Ulht/Vf8q0ZR33uPDAF1ROSQ2nX/aIPgRxty52hGz3ttHoabv+r8dheUrftOQ9k
FcOVRBY2O3Ebm893CWYX8f7UQN4T0ob3nJ2q8bBsJaAgTfut62z26XjHsIAySSXy
jqyU4NXqoywVPFcXfreydpkbsEW4bzqHkpo6axmlSkdxBVSf87pJE9OUcMGeR1Qe
pSv7VQR8oDKsBsERNyYGAAxglQ7db0t4GAiOOODR2qpZTp9Mp1puD0Z20ifFcUNU
p5LfZr5TJJky/w5E4SNwHSAqmorwMYFTKwjMgu+PAj1bWc5lLIv/HH1IAXcT0JZ9
z31bUIrKo8BZd/wAAjsVQZDClFEpNoEHrmjsMVGiXhKee83Hlxi5KF/+TfENShZY
xGwUa4tDG5oVZr6g3FIM+/eQ8N3tm2vbCB6o8d3lqv0KNoo81sBvlJeRYB9lRLJ7
4T9r0mwIA3V1VPDa0UF+0M785XQvBGA/INnLtwg6KNcry69XYoSkHh5fZtvqSu92
UrZBEq01yM0/J4/5Pz2cOH9DxweX556PdEBHKV6xEn16sfuOzOpDRy0MbvggJIf0
cNsKFU5F3Bot6enFMoNJGZuPHivYm1hF3NYjseNiQrBfIoe90gpE7VOWy6hBkKFT
HtwUwffJFMwO65UMPiP613jLc9GZKwIPPZb25XmuuXHc4+0hEI5ekNi1Vfd5nbMS
16A7P/+0jcekhZs5aSYyHnXmkUsn/dJi/pxujhibj7PIT0lRGueS37WxcAn1ykeQ
krAWnSqROrtdN2B9+NyRfRu0DrODXEtd+Pg6U9aJh1PjYAfSWnbalAkf3AOn/fC+
wZImPTQ3AH5s9iZhRKl/pxyG3xnc+H3BD9IPIZ5H0aOkpbavKHaeQbxGra9Cctqn
woiTACSQR32SuaFClp4+Iuj3uLhFJ9gUArufmBFJxKl/AERRq9oWL2AQuJ5RHfC1
ObvFRF60yIJK8Ch8YvWTtzqLdqlrKGzctSEw+bysFTroxEIimNuCtDHpzTqBph8k
3Lb9IIwQbaD+RIwJYBylFXyapIvCY/YUnbTxvSdzzeIjBFf2Sn6VndhlDCyV3YuX
B1vN3ImN9hCb/mtjS1ZY2sVJ3YWHWf8wUPvEUX7W9mOMm6xUKLIJ+HBX2BGa4jVA
nJ2elq7anasYQyHcFH4GygnKVRbA/qxPyIhcqPIoPoVTWkrtGwetYjoACqxnktcL
y2HRqki7Clrz+Ee91MxeCrKXncK35Spfhu+ciqweuH6zO6p9q6lzdfE6dbJtECFI
qC5Rt91sjqvdYGcL0mFwnGEgG4xF0GQLdipfdVLQBr2UWlAFlZDLGbubmf1L3Xg6
ZsiKwbAKZxXULB3cY4P++BVm1Czp1QJX5QXMdSyho2u2ZtT1vUHmCRAa7dyLptvk
VUpqXqc/u8gug+p/ITm0e1dYTUyg65x2W+s+E3iEil5kvvwYsLvL1oZB4l5mSJNw
DtZWCVCnx8f0GB+6M/tSAHBAsAIJoFZgCZJRH5sOlAYiRWh5FtanClLcdyVBC5xx
bvkQO3M9jKV/rFC21uPCifT6wctJLxqMav8d/oCmUpgXdpgxSXcU0eh6II8SseqY
McaZ7rvLFdxCVTz+BZEHETgS02C14KHdFR5VOuepBaLr4MUfEWHpez3dt9LSihcs
KEB37eobRFH6uLTO6T2ydtnnQH2nVTRYinbUIbNE8PjDbuWWf4Z3689PFRaqrkuX
n5foxfTZWboicNg5yFn0wKDSteRQB3mYICzTvLQQOiNpFhMrSnh31U3yV+3Efy0f
fX0a9atRHutDFLKvdYR7EWHBbCw85n1g7KlYaRPK2ZrG9D0+98O+pu40uQxTYbHO
4R8sEMpW5dexV+urOzmwvk48pzGcAA7tGKQqxSRUKx/+t1G9DFfqUcVx3piZR+/b
w+qy1ZcoomqYA3A+wP9knDYKC4zozxvBo7uSIr9cDeSmi3R85aQPhhUk6rSq9ZS5
MQm1fEzBFXzVjgAspTHzU1xwjBYvqBnpzcMHkfEX3iIrdmbHxg82WbWfAx1UG5Jk
I6lFcoWwFAcC8tnontKTkf3yfmLa5GK6hYFi+82DWWPrvDKuGg3E8cwgunYhzYak
3wlvoExyZBgA6i8CXFk5k6Bhf2ywBK8MNxiOiteMl9c7dOIXBUG8J0ezd0hXctp8
DoFk79+NcP6pMB3N+ymQxThnGZMkq6vBljoMadygdmJt5FM1u7V5PqaPtlbxV6XN
FpDohSompinVHBQo/xxLePmEmHy0CHoS9rKt5Rf7A0z+c8UgIF57JmyhWdCrrY4N
U5Ecjn6S/n80eZdxR3M9OpzEoBkZ9tHj4K/vtsJBUQWia+VAEXVHtZ0Xc4lI5ZZq
+dFXdCkbZOmFBTQSclO13OzhTKTFw1S4g/e88aAqb6k+67FqITKtb3jCfPVha+O4
fpKeg0bmKAdsUMbRAkrwgjqsHFs+htL04l8BvyikmeRRZzV1KXzek+BVC1K4BkXg
u3IlVKdRuuJcJAVFosYQjAW2wd2WzYdO5FrOeq3meTGa4XJNj1TZWB9TONhgMKSj
5Dn8K8wvxnSqVpJQRF163+5JjXF6dpB3r9WbAJNfR7sEIu8oR8nP96Rdx3zsMkyN
MPSDSvbmHRETgA7ue3RgO4DG9XUhn/HjcGICnUdezyygNm7tVigLYv/sb4ExP52Z
ijWY0xHjkvFIL9eKINgtoHMAYCaBVfe4p7OeNbSPWSR/oQXyVkxTivjES+OC8Yn8
d4m3KfJbWNCZ8NhOrJY5IDWgTMRM8IzLg/6qo6IQc2l5eAwZlhg3xCwIv3bclMqt
njmPvgMiKYtV/ucfM6zpAAIooZ6Cy2lxxULCqNN9NhskWegVcFUTmypRbwMxUeC0
lLxEfaC6coYCNTBjnLVG8zKIS9eL2lNdHYcIYaY/c49AJLunA+YS20WdTdujEw6W
y0CVuGsicK0ptedAWg21dwLe0Xe00q0KAHmqdl8Tmy2hPWkLnt/KojKky1sgIUeR
Y2Trm6zNQ9roPUiRIj3Apk8yZfHvehI9LIw1dzkM3CFoFevbEZMRhvoQVfUtjOn8
DOmrMu5/ZXU2VpDtydjxm73ky37T5TqDDxIsOlvzvFojwaTDgzmFfJgfjorE+kV5
LI5g0yD5Qqv1Bbh935ybJSMbhjJcgx0WoUwN0eIqMiOnnftfUX0TlL29U/Q8toTF
DyJo852tEEt1/mLKWJ0XSPZKqsjqwmYe+6m+oNn57Y1XXyrpbd4QgvasrJCB67Gb
J8gkCbR5Lf0tDIkyNKKtWf6LtFPpeANSbtzRvIfr/F0aRIxq6+67U0Udm7Xao+Br
/TEwk9X2GesW/v/xOZRLg602ICl9pCtHr1aXPO9lUwLU/F/4dU3ua+aP8EcB2LtS
BDPhTCUF9I80MXhibtHwgY8bNM13V6HbGt531tM0Ec/CwmkFWFpXDSbmZ+0ZjtPB
I6BxOBzYKjmy8Skgnoh8VHxjAQ92oGw4v2NC+G81yWANRhHpVx62y7qmlpLmPCEh
dfrjivUdqYsNgmyE60iUrJoPKCDJaqT8pV7RSACXrMSyM3aLo7VWMV5VERItk1lp
XjCoDeBniubFiLaA79Jl7iFuUri7UYXjtBpp4CDOiNmeDpsPkh2s0F+duRGcK2td
cISUAdpuYWRbez07yRx7mLk3O4GwbuoTeCLVXH0+I4UO/zm/uLNOF7BjngBHPtY/
7WXtDsknjAog9JGJgFEeSJPlQyEdAJQIZ6eqNfE1ubUikY1kPpwiRdfUoRUQpUu/
Ql7YPEN5p/BLGkPqJ1AGr94K7IUUGeOAA/7La4dnLMOYE04ODm5Q/bPvLZCBv2Sr
QXsvJYqllNxN0C7Abmm39rCv/Wd/bI2Uo/XOu3H55PLmQiqYvXK/r3ZuLouhujUa
YVxqQ8u19IIpoP/PM6Z8s8v84/gKnhJap0Gg2sI3rm9fmliJDOSIWPcSbQvvg7sQ
kNEzKtkyFizikoPzn6r6QsmVRETi9e7rNyOyxDmoVDmOBPkIMbSiRHQS1jo/Rheo
DhSplYOhtgBltqJiInP7JnVjrf70NEChHM1yDZSTj6mpszbXAyI4L0s0lq2RmUSj
GlF7Ts50mhIGVRKk8Aar5jo43pdiYTIx4bmdN1uIqwkKRUYhmMoHCqfJnCEvlFIQ
H40w6O/VIFmghmMkzD/eu9yMIE3dL4GPPKMYrIMKRDtZWMBkrzZQu2SCrZ8B0M6L
I2LNZXN3JI8Sb964y1band+XlkswQEV31EnNcPqI6Z6m0X0yUlJeOgpiWkk5y5Wm
fACDUM66b6ITYH+NJ5MpO1uDE8ieH3A77WpElab0TLhfsEmshoLzOmPBgjrOOOVj
WoaeSmuN58adoWxAcqbXj8oZlRaX+9hvXsiM9B+vVrtjY2hnnU88siHj0J86Lx/u
LMP/y0KitA0h0/bQczmTyyNHgSqKg1DlltChVyW4QcJU4mYij/QYo6AfrY5TNhH3
CeWRZFxkejVqE9X2Y2Xax9cXgnvtYRqgguOgHcNSGHLn/FXIsPFJBRrxnHTJBSIA
X/KG4g3wWswusZRxU7RVjJRvPcfe2dXQanwuLNPaqXJBXFfQxF96OzTtRYaT2CsY
mjtHuRMCDWn/o9VDm+tK6l2WFCTvjQIPRJcKPjnpYgh/CrLamkRKICBhAmSjO8Fh
VhNafajd25oZWYQrEHcD5f1skYUOL5C8t1ysa1z3xSOc7mc8wk+lPTqqUrc5k1D4
eo4E7Wkh019qqD/i7F4x9pKtHk7Cx1o5i/qnbdZimosliZHv+fMZ/CqET9tzMbAm
9zpRnzfWUqgMO3HFZ+StbfwmsEegJiYMe6oicHYJOw62Ug45rcyJeI196xdsPfy1
t7zc+zPA8MtOxoYNJhnoCK4Bp07gOBZo7N0k9xK5pB7uXD3b5vg1OtntoU4cfvgW
PTDV2CyJ0gmcGKpGAEb7RMuZq4aPWuAcCkoGAGdzZq/FQrYeZ4icQ+19wFdL/XxY
zsnZZqSh22u7U1nXKUQLeHLqz3f2Di6LwMNKvVKN3IXsvpcnLz4lc2iUzlUNu9IT
qzu5GOpo331Fmk+HVczG/TwR9O0AjyGw82vtLVaPK4wzE1ub/clKGxdSCyNTx1+X
3InYkhn7jpu2Q4Zu99zv2JYeJFxOM6wXeWqMVzwmabWs7VNH48gjKyNRLKpYHO/l
5fkG+IQQMBwCZ3S3bM/cB+w/1zCJ5DldjucImzyY7xnqjQOxW4qAGFYAyKGqop87
9WGL3zAtEbG4+FDXktU2Fv6Zi9dyPrGrIEiHx90SZaOv9HBWUqAiZfyASJ8AlWic
bSuEz4Ifns2XWCKV8wuyzYgTM8yhb0/TPlClqO8ozTdx1Waj03uwGDjqOybv0cU1
2GX0PU+oglVFo4jM833ibCxzZjF5ZF5oHREoSTd8ee6P3cIGSFCcSyfYvB+GOLoW
uAQp5/C29Sp3kky3cAqFueuJNIlCWEe96JzPoM36h3c/O4pzIj7IVzVLBBHn81/r
2VtzMXL3BevTTecle5JdI8EAlnVSM4wlbrhdkBo8yzDcQXga5AED57LDmObBuxZ3
JTnV4Du91RacLB70gakVmGDVZ/w8tsdJU6KhIwPS/0dXM9PqEOUYTDcOLeOEG5nu
wQ1+B72A10NHW8PwDljikkjbXqehfYemijUQSRebw2GzuXe0f/vvJDvrbMpfcGzN
O+Za7KD9kyBIFYzOAd/kU94OR1Y/XDhuT4DcClSSHztcYmmlREW0h6pWpyri6k1t
yZD8RdTHJHM1vY2ZZq4s8vrKu2GwkHoRw1dw2bdmB/o4pbpt4TimnhAFd6VBaC17
xRs/ErAXXO8uIlnWY4NWtC+K2ZQvrxaLUzZDf/6ofeo5XrNCnsKkQPnA0F2D1xw5
OEzWn1JRqPvFjPbZUVHPOB4YDJCjjogXywFWdqPsoMYUhuSs4wEVufp4Xfd+ncEr
vDXLd974OwUp6yEcX92T/miTCN/JDcvWQp9oqah+V0aXy1RaUo2yTHsiCfCcj3vB
MM+FwsUzN3y/6j8EqURCEHQw/NuEWgfNeF46pmmcvNV+tkTaufNhkNhaXewIuv3q
ZusXEmPI04gH3L75HHxA/Q+FCKZdfUiHo7T30hBM26gqx9lVimxV5em4yTKwITqo
eKzIHdxD2vg2gsQj158JsovTL/N4W7S+HKCcd/FmktmWqyUZBtKVwA+QR20tmsst
7L9JNRdOVngKydKrXOXrBBappzFgHxUitWccpYa6vcMOiUDN0wvmnh92gkuWB/ZR
FVQVixTiQ/6bt5WUsQNka9DsLd5IfpqRIC2q8kg16MtrJx2t4jyDv4zP3Fnifqur
qhkJii6sPFI8l3Pxiql9nM/kJBIBqvVvBO2a5d6HaCobdzieFgp/dYvWqIEhe1jn
XQHfF4HkjPwUgB6hBIg6BrN13erw/ed26mcdix6LGrJ97Qzf3Iaqm/kFV+Vcc+tu
ObZcqCWtTJTysk9LEiYpbMqS+IuMMQddU5dzL35fIjiksKbGLhkShZzx/rulI7V8
FOX+wyJBReqXIcbhuqResj8YMVsEeCvovDrTq6Whwx8ZUENT9hVgNvxcXho073Jo
U1PwP4iNIFVk/RLiwCIaH+wmHMUu1OgTr1SvQjU9r2grtEFlEB1a+1gEez41VQeH
vu+mNtwnsRP1dXuUsMuaHOuJyJuEO4MoWfbxM4gC3aX8vjX6Qo3Fj8Em7PMuvzEJ
vhae/LvJ2NT7ZTA87HmH0TbGP33KBzyWdDesRIFqlxj+L4ke9BB4RKcx5AIDxZGG
9hDNA0yMkSDkrT9D8Lt44YyLnscwPXejLcmcwse9VTi3Nnzrehwc6CWWLikiLwnL
NAM0iRiQbUWXVPKdkDOEQ1BCiqjGISyKX4smiOdIFsPVUSuEtLKZhKmz3LDnTrZu
PnF+mYXnV4YRaAkqyl6ag5gKPkm9kizHlVF7nJV0uZrSWtUSqGyA+S71a385KSPV
MSyiminSvJMpPskAChBObWpBURF3Mp9HtMg77NuMsfqkAdELd481I/Fv6fUKlYDC
oWlIs2oeCMnYULMQbjv4rl995LzdHu7h8AC3OqqFKxqLrl2RqjbYKzvpWq3AIulq
X7fIiG9dTxtaAPcDuy8r/PyqhJ2/ILsvEMqXEj1kM2hTJJq0zqCgWw6Hz75UtJzo
ie53mWK3+ZQjQv1v2Ri+O1s2QAq+PTnTSnNfsyAVRuRvpBrcDih9jXD5WB3BXifN
hKcsFoNaW3YC+fIlBZxUL1QflQ+d8pLZ/cXBYo8FVOADZF55LuvRG/j5vE4A7YPc
J0jc5xJHXSCVZ1Cb48fQJas0+OolMjTj9T95OPFmRoLxpVoF8orUGP9FSf1WFGK8
oJZ66YMEBGXqPLrNu96uQH3b7U86bmvhVsHo+0kYnjIsgIG6S8aLo2OqXtcE46EK
tKlJqWNdZ0frQPqYldqGVEX7LynOUePqe7MmYaql/VU8SeFo6NzyOIQPCCmoR9HQ
RZUe7kk1oGwQj7nQ1H3Tz1+iccO+SBG0Q5tVWS5EFWco0BEoQdqyMVtK3Wgu7BNF
nKc2pQ1RrFoQ+lYwQivShenfaliW7jHYvFGEqdM08ywMe+vakBbX0dqf9Up3WRCw
PLiHZFUJCBnMgB0d1qXpCEIqKU6qgm4nX1CSzPw1ZeazG0BZGW3gRz7R7NGtNWbm
aZPiToCtnLifm5nVEvuy+IQ3NVpSMDJuAPBAbRMPgWmIbiBHhfdcB9M5XzXwhDRc
NISIuKxAev0Lx+9TowLI73CaIUnWK/CB09Ynw5zwJAiWDKRg5iZhp0T+XlYHwg/n
UU5V/4eaSdInPbVa7VbiFNTSc1wwPefcof7GI6XOx5mDsV2O5pE0klV+gyFEjysJ
x6mSl3L2vcdR2daQpr0gp1rONJEIRiFQypTrlCCEldUMhuRXFazBa63WyNqm1otL
qTPY9967CL2Sbd6ZXW8IGvWCe07yZeA60ioIG774spj6RGMfKprgcjevWW7SRCaL
5zG00mAt0bvJku/JCWS730pJr0URb6p/43r+phA0z40FTxJxZXTFdRQcr3Fqwo/w
qKhVkqkot9X1aDVOy/IXReBzLDUuyBuoudlqTeSU8NZCmpvnXXzCvtMkZw3knAdS
Mzg7BktewYFDRoSGrqZLV7uIHUZ/7O+k85uQwGgvJGuoQNlZy8klKWul83U8tUX7
ceMcyXBQuWe/mQ32HIjVn7wZiyGmo7pxGolsfxAYfB005g2Y2bvorIHwqp+X5Ttr
Wa87KcLT30S4P8XE1+dWECvFokTOE9O9X75oONWBZ4HBOlPT2wOVwY2el7U/CJQQ
eFdRtzG7fWHsSdmBeJ0ClcuibAVvFMu8O+yEPi90RXGTm+2epjB0r9IdSxvj9IOy
N9r8+thzVWHqz+thZK9DACtuu6kxhT2JqPHBj9fP0iZD8fRvbg99NBwm9A0i47fM
P34uTEDJ68TAtXJuFLfOd6dKleAxbDCa6seRvCxLC+nk+pBo0P4oMsRT9VMMDwPy
3aMcIxK90/6dgUVESGxTGQsWIf5hqzv6Dscu5hqyU5ZbpTkpgsjfPbS9LPuAG3uu
Ge0wlafcK4H3y8SHeqRg7oMEXKFkxxPu1PEr+CqYGeKyTw/cBarK1fu6FNtz6OO2
u2zaL96PYGPpeUB9KYsGwjxij1yyR+VBM9eGIRg5J3Vmb3iyC2sTN7JcHp9cIqZS
abCigwFNjQ9WM1aKnRbwrhEC4ihCeAKaIhXSa/8rYnR3HE0q1Ts8NCbcRFxy51Mi
E4tkjfqcFq3c/aZczefct1t7lA72nwdO3D0UDI4wjbP/P3/dkZa6BYMMgZnH8AFb
u+GThSLBa51v1o6Gj/fPjWd5pJAhWM6TYok4pbU8nEGeI3v6t4JmZTYPl5X3quAE
qNjOj6ThoDA+G1GDq4KBsqkoOPvWVpB/DhduHQDKmkVkDKnK99u5G5kkPMUYC7se
L/ijFZqzcBeiA/Nm+OnQ2wBdrtya5oujPB+JVtsO6OYWktU+MST6fnIlIcso3gIl
+0Z3+djhKgwb8prpAY0q4XXqgQGwq7CbAHNfHp4nrDsbVkb99LQYYChQ+X7RFyDR
VojaJbxsPM0bOoee7HOhX6566vOMKdNo1nrCqQDs4W86MV6ead/1Z5pMiBT1ZbkG
aKuE1F0GNgdEtwudtprbmXbI+VQt7Z8lqHl5w9tv2hPFCOZQWEKBGTLWUZhUp56y
fl3WAZjWeNGvKyKmZqKX8j7sgeppbRhRHQww/dckBPLt5QLRjX+2vb79kqBqbq4i
I/3fk1dUEdxFLmS5OXPq5TJBF8H+gT5nLfA57wpLqbgqoI+/gYC7UnCvXZPZkEVB
jnKBRo3CGkBafxxPqW8rgzCfiR1T+078Prp0cgGdqmN2jh5PADUe+57VkFf34wwT
XLiExeLYcx9K0DsFOW6B+LrXgCw+vKuBfPwk7yM4dgYjyn927DK36bBHHUlRXBiO
z9Pf6YuT90PTLKYOaWP/AlpOJUBafuaFDDltqBdHN5juOlliOIORGQ/Q2dyE7Qsc
3iiq4l/zTTmdUjHMBzq2f7sgjoAOpScFiXgdyMC2zua9FL2SEZ8HPF9zhvJ9IGFg
SSI4ImMS6ZxnPcPZPqUsaEg2TnWI2ZiCR0/ZEzXmC/qJodDqrmEAgfAIy2h/+Xdp
n1mrwRomouWMyTurLtiB6EtsKW6d0XVNUZ/sKxR097915tCjow3LzgO0jJbeDYVf
nCqA7hgcoiTQNA3nIP2jlCq+dn2Yz0mCHMrvaChmPLAdjAI/uf48EZ/8b9M6jJZW
aidTDK2GZmYW9kJX69iPRwrQZnCxDgHBUXix+7Zwgs/Lnu6kA9Qb8nk2mO3YbJ8B
+J+YEZLQ3HNTHBGMh7ots8Vdv5WJTiLl8w3PhEstB2hHLVwzzBO/mJNYuOQVQICh
cktqwU6BrjcpkP8H0yo1GRon4K+Ub6pL9IN0W3hzWZ3IHlhdluatkxeSmND2557H
PJVZSpFtO1v870V7NWWAXjY/aN2FQ+nfofT8/C4VOCfldsZ0rmBn6Npuo9EVR6Qj
lqtGZuHW9kUHIvM0IJXf+7B3tRErGIyvmwEZKeDeO/kZqdwQXPT0+I7/i2eixEzh
JJtZhry7r3GHJEVWlScsW6CEPTUBqJtF0E+MuloLJH78/mk39pWZqAkGJcwRV+F4
EfWHLUQQaOmJ9bUAAHWOnD/pTlpMFWV4Zbuec8xSQLwa1GAaoU0LriwwngRO3bth
OjJv64W59XMuB78pp62u3cgqUJdHlDEuh8dHcACPjnU/ga8uWMoJWqpzlV9adfE7
w2mSbsQM/6tBhsZ/SgIZqhSiVt3ulIQ06+ShlD9tqvSepa6uJKbS/hfqo7j204vS
z96WK9Ea0jAmF71GtK+BGvCm2OVTKhGJinGgRHmkYiKjLAXb+/0gcpCDUBZwKhDl
Gd60SsNxRKprhzIL9aLEX3R2cQZUKW0tWVtbokD+p88IhTmiwwkq8LD23Ump3PjB
0bXw2jVr7nkQIrpnWCqnV7qyd4RyAUFSx0rfaFiqJTRkZPpB9/SX2vshSzTGc1cp
4M53ylZKaY1+JdTxkkOKPI4M8dk/oq5FJytIcRH7ZTSRoO/2mGiZw1w+bnZDp4Qe
TBtM3iveh+k1z8zHbt8rduq0KB03cgepxHSssIEycVQlEIckSPAN8MSwdk063/DK
vV8+16AW26ASCbT2M9lAYg25C1nQZYQwGW7SrL0rWZCKt2AvzKX+JOyzcZSrzyNc
W7UtXoT7pvBh5RdjEiVr6T3shoXZWsdHMuUKxsfnWXjV+R2I1OuTbVufUYVpETte
H41xQkOoxevm/kuS3jEHTo4UFc/Cnh8oSP4LFI5vauBdwDodjaNH/Xg0MuT3+o6x
KJYpNIpcZg1UhMXamXqYXgj8kdkIZ/L7aSEA586tSQIycB4TUYPSn5HqVIvxtFyH
JHqsWHzE2dYDwwr1Q1DWe1N5vbolx41j7pMBo/+4vsjtB9IysR4BTqHLVQUREYPW
MgHsHt4aGyNL3++rjtNeXr+5oXOdvvZSBHJ4ibZcbGXFvN/0wFXanSgZ9RKAPA0C
CJupu4LuwhevIOIftxzIHB+o0yr+pxWp6gdpcYhIWX1+H1SdBMrFIhDxIYOWcdTm
Buhz3vqnwiP7uNPoVCVvfDmtVVCO8gUgT9PoznvmldtRW29aQtXPSmOFc2GOjmys
7D5bY/5WcsAoUAkacQ5gkPg1MvaQVV6HRSp7x0IZ1thTRpuOnsoyYpi5i4df2beD
WTtXyqpRQlbkCZnafi73ZphA235rktDJIOxLddLO5YcoJGUoQMTAMzeBKnHn0iAk
7RiXZphUaBqdb0PVUdTvfZrwB4iKMQXXoymzSDowA9heqGs1cqSu7aMkZ2nfjX0k
+hNLl7E4MxndZIMRjeJni7PrOgFe/sWIzHfmf7HftZMP/ndjyEziNE9yEHEqWQ+5
2ry486ZeSVE4E+Cd2zyg3mTdLquOthPFoEPgL4ObrIT8tdvs6y+wsBpaj4zpf+pX
BPrqD9PvuvYdbXFNnPhB7AoBN0kHSkSxy6Qrt7zYGtHtox6sBVuyNlhlj5mCrxB4
+80zxx9fvJdolUWwhWha4ahRqrwodCRjD5Fad4gTaSp2XTU/PGcSMJ+U/9C8YntM
uGwMKrelDhcmNHqxwEBC2RoZ/uLEh2yu3UvAC1Rld44XJqjGmt8BVpPQiwVAmONC
EqXwfXga1DkVOM9NRnVmLGjXYwv5y24RmkQvlI6uZUuAyCboQwCmn65BAGkEEfDg
tX8cMAETqeTZkWFxfJBD3Ts0RUqCP55KY9RD9mgetslX2kdQlnjrMrpX2R0iwuIA
ZfB5cmXWzYiIgiHsf+l3iIZV4Cn8xQXafzFj/0hHLjcFwuHIufTUmPRQlZ4Kex46
3euyXqZDeUpUi+ghz9HCJ5EAtXi1s5sxJ/xM0MEb/23l608sPMMVqOgLs3DhmzJY
Tp/SQlrfYcGO+DFA/CIfdcXRC36RfaLR+dQEc3rhG2TXx/5qWqKvaM7BYwzCNDGL
umFySi1o0S6G8bm9Syl0m7wmD019hZkUHgHZzB9jk/C+T1MaJ3c7hMG66ssUbXPp
VL0R7aqxOENWiNwVNPS6TFB/1o42NAfSmCfBskODNmxZAJqK3k7XLZr2RXgVLjf4
hWNJE8hh6PEOPwaJtzUnsV1qEWFCdtDcLbiW6ACASUN/VKc+bTkgErm9lktkzV7t
up1FNEQlH34yJsqWQlSjqKITJ4gZsQzzxYSPVgPwQ3rCeOlg+wzEokAZSU0jlcdb
wcrE8+0eqRypX4Ld2aUzbLvIKMRUfnzV2YkssMTWY4oXkJQsoZ9Mk/ykCNSAVT0a
vksBRgwPhVFci+9xxnCQCfhuX/aV2qiZlXHLP733lFGO60rNoCvWfJRGW61FICAk
LMgESpCLlP2Blv8XUojattuKAFUMKUApP4Wtaq0iGAPQX2SPHtXHaisk0+DWOdGX
CfAV/kcAbiyyPmIoNcgYwRNPzdtMZJdqhvtMo4WEqQC7hDiekTaA12lj5JScTZGz
NKJb7eGmwYTwxqz9eG3Fu1Ep8NInqhLUaT7gkOfzmHiJhqpMLsG4oj20DaYa6F9s
IKApxzkgrT4lxah2vOdDlxlKJAiUj2AoP+bee4KXdrMDuXETsleOw08Jr3Vh0oqp
IftKSuZp6lvePbuellIQAYipMYwhUZYEjZsUSBtQgnYWGVpkq7nzSRnRrnco/cjs
xeG5jP2XeLtw0zZLMmajkpnfyNQOIoiW4bJ6R8WluMSOCjYKzSrm5nJSee+Avado
mRXU+UhLXIPIiD2bAX/W5iYscKbrSEspkYkdXrooR2VB8RahCAcGpcC6DlQCHwWK
NDPszxgG4AA/eJEInvvnm9VyqCNcU2fUNSWaj3Z/Lx95kH9vLXmHOH5x557o/m1O
GpT8AoUvsbVT0Y8jkGWq0BJKQ+xeqoqp6UUZVZUlNdH6iLLi52zlCxYtye2Po0uu
IUwE2ojxVwdlKyH0wRXZRvY4x0XNp8iB6yEU9SqM3gcRgfNafCNCfnobGDvnCQgs
+qEivfRXFgdsxFCHSDryxUfTeVP1Lv1CduqJoYlE3QgrmPNmeznACK4EZAlWD8af
ZZomar5PD3usI8GW6HROFKVdC+thQo6iBBAsmh4MD1bimM3hZkZXANKx6R7fHqIv
OJ0MxIekKcGP49CQOZKVnf+0tR640uKfDaSdtottRcY2TawqcZhzNNQMJ9kGBNSV
1dscvQoxeDhVI9GgUtbNVMu6gy6o/sCy8G+Zpr7aZJfdmxOwJG2Bj/ieeSxke40w
vQK2g9+8BToD3+w8noswgPh3nMAsYXV7i8PoXvkCLEmyDqUCEvVNeR4AjBJjDQGz
d36VIHIRWfHxWzGRH4Eo059Y6XXrmi50r/sj6rlML2HhH2OAkIT6+oftRn+mvxYT
cO/DBQ3ygaWuo0EKcca2xLKW3DUbh7zhfDqV1rEQEuDcVmbRxyqEjGuC+/4RyS7R
UA2s6kT5kqHFPsyqkmlEGRyo6Z0rZ4U0asw/9dm9ZOzV7IOsooZEop3lb+i4z83o
Ay9h4ucTACLGgrOFrA6XvsXeJViIwyT8yxIA9gNuvU9WTt8FygRu3rlyD596qgrT
ahcxRh+OlffySh1aqrKaa6FewH7JNW0hy+m+FywxKl7GfuzmQM3W8CKAky7a7bJV
mMfts5NuJkZSnCSVwW9DibU/GnTHDoRw3ctv9SOBi6sN8pUDlyFSVMeNNPetiiwE
+eU2jf3ciFu1t6zXjguxVT0LBhNMOtLDU/KlGs5Pe+mNW0ph38m9B5eLnenKUi90
88PwTwC0R2IUelby/8/gCUe3/BAo6X56Ivkfy63Z9zmZF4+9Tb06zNALWWoqrH6N
xYe6FXrEzts8QS4cvTxJUBToxeAZfHdaipkg8cMOZU8QWodIpmsrL31FhL7nM5jm
gbGjo0zuPnkTKcEr6N7MGGplpEn4MVUYQEs71BtEibENCeJQ3zX0FJOXxTAnhtjj
wEgBxU+xdGAlKp/qs8Zja4maPBkaroUzAPHYGHaihbevgyLkT2srlcomuRUH47d3
c5n8SSSf6CDwnB1V3JpaS2VbtwZAQVLv+C04UszCqo3KcJ8GjOC5ZtHpLZX45DFy
58PnQhfKRlMjPvwEe3r4dbfBeQX7ij8sE08O/RiOIrKzm6Whu6oxoCegSqVOcP7W
xIzkqPiCxHxUq7QQO4OA0Qh9pHRXx+31yoG7iUz9q8gSYgCLoF2etD8BQ3NWxbrt
RqNrEQZ+2xZTmU7SbePlO7qN63s81ElNqODZydjBlMQl+t32BMTP8RK5HCpTUMXe
HVctSqe3MBZZPPieCJkLTATunFunr2cT08teD6KpppZRhwi1irgjK1Q4U2mdYGSS
BRQ2Py/BbDwe6iWtcmeW8u3V6Y5/71hSGDSfOsKvJG3xOQgiZc3LWKvBKgUietOw
pd12TYlhY44YWzXlD8v3WQMhIDoZn2SVmcE+4/Q5TPBRaZ2xEzDy84lIugYr1z4q
y2XakPETI8ACInCHjXI0CfCv6xfF6n+LOo1x6qJUVfNpQ2vyCx4PXK/4grDI9tgo
SqwtMBIiSlupTeugoAEi7Ja5F9hnEhV9mv+Wy8VCjwWwdagkr354ONVYjXiw3stP
qpATI8yHyUp39ApB3urx8whLPsfJMV9gs4QU5S1yNJ4O0LiHmT9SbxhMDiPkqDcv
nj4+e2nQzYsn+f2sr5r+GvuokpBIsZldYe4CIPFgeaB6osRBqd2qpq/q5wgVjw7k
amRZD0Vlsc0rlPb4CEhVoZnH3xfVRxI+te9OWXyQ+GrsOPrhxDrQo0besAA3wq2n
GLvKgJ317f/xAs3tMu5qsGTGW1rpCjgl815hYJu5x/iLqmpjUTsKbHsGA/2RIwXB
eOH4eE9RqaGTwP4AEKWQrqTg5RKL5l7Gk35N3hvasH2TZ7sWgvD8Xi/RLle9jGdI
vQconNT6jqyGZDltHH2m42XPLMFQMr+hXd4P4D1ioPZod1RcIsgSePV40gMTx53s
8ejvdUgDKi1jk1s9I3KuElDinIeM1Mo7z65/BAEFVkoO2e5HRGr3p2a4AC9p1nND
ugp5ATDtUNfnp6cUanZDJy1QP6t47URItnY/t9uDKwdWCmYKQYh9qC8aWvVlFwvW
ZoEaIqeGqpoVx8uGN+KdaHmIDW7JUbR0U78mFeLKUGtxO/pTxrLTS7Eh1E6H3Ieq
RUGHaDNJHmYrHwezLQEJpZHyofAsxYmEwlsVOsiwKh+90ShMrO5YzE2jsaWG2aAI
2taifJrQg4kNxtRKNVzG6Ldn6Zr5FOEBKJaZk7O/LZizCjTAyFrnevbjfzG/mOcT
rRNrRIkuKb4Jh7iptzJmnkXjSR8dDdQ/yfLBFARQSXed64oLWkbTcq68zeAX4PrZ
3PDoiCtZWftF+aNrwlpXiHVv2SXbUkNW+Ftf6KVsWgxTLjumryvrptaEir6c5Rq2
2sLyFgNtCTrG24gAeq6B+PMCuRGCIBSZC14wKfvhq64HvsJahRiS1Z9iaJ/bA8cM
j/pjcrXhy8yn4m3rgaywYr3xX5yFmT47mrcpwIZXyJbidKE3HHq66WtMyU4YWfDP
QCBpb2v5J+RwdDHVJ8dzyUekrNlLgv6ypEPekvFg23lzEvG8DTCiCs/kS/XCC/fU
bVFitKmPZeOvF1fmASS9XZU37tNdu9coGp9dGuG3/8px7aq4eCKCohhpi8zgx3RF
5VWcmCbJex+qeE0R50bW23M1ZJsCJcH9DSuTpw1zwKdEWf3dG5kPzOcwm6qkdIYb
KyEbt/ykLk4iy/kIqVErjo+rxrneZyI3Fu0uBjYiD3S7Kw9Th0NujL6YdRPrToDk
h2Or3TYJ+laQma9HyLRv80A3AGFMi80LqvSPtMbcWD+lyGBxxCpr9L4ldb3Wo1Dg
p/vmz7gSXZJpsl8mVAK1io4q99YtH+QrE19TdnLF+00E4nB0QB1U0HhnOIiza5h9
e7gW5KrM5A+BQkAQfwvPGhR5+N9sFdicPUttQ3+y+EDa66XfBLxH5tsC4tMA7MB5
uPzG0SFi+Zy3WDTMt6H+VFmJMvdtKRDh8/KaCyhZdisStdkj+CGlJUv704GnWJ9O
kz885YbHjJG1dkLm3MT+bDrF7LOQIaSZo7UWlwFerN85He6Or5eXytoCLQwbQOr6
UThhYv6mlH5PiVPEbWO++EjAH8NizuZZNe5haq436li9Us+XwFy6AE6+m4nx/nHc
nq+EQJKAmYN3BEwPWOci5LDAdrwGMuEM6E9SrVW/1WzXy3bch8tDYXgQgaygFcKs
8HiVA7qk0qK/KvuIwCGxv5JnV32dBSwBddmcdf+MBist+U2FiXHhj6Xix7W53Iep
qqqFeCh5m9veYGhoYrpx3EvITo4JHTBUnAnwPIVAU3guMeU/BTEkGpg+Rf53bY1L
LeUUoBxFvAgFeYw8j7nqpCPjYb0occIhu1/5xKJQGNkhG1LV3IG4OmSHZ5KponvK
Womq8i2O94p2bZ/EyF4aI3TuAecOyl/g75apt/uMxdxiMpDEGNPfKHnMTH55EnpH
t1p0u/cU3jY4C9i2U+k0dQyL//wD3xtHW35DcRjZe/VPEN5gNL9OCcn9o/I55a2t
x16H67bF4Rd0YDtHp5AUcpHQmlqJHUrp28a0kmhjfH2IzUmFHSz810uPAVqqYB6R
PEHTSdPr1p2PwTGWO4B8CFlO71yTZUJ2h3pGk6kpicZh71tEnXYpJHq4GSzmgy4t
NAf7mr+W5JjOdL5yx3O+8sEgSixxIEy/905dFQYiC4d5y31NI3Pyvr/Cs32+h3T3
Lb6iSc4XCjVtsap7x/uwghIKsZ1IlWkeuws3hdaAwAcHjIPOp9hPTAGSAimwWfcF
Coes/C9pqh2XOnixStvpUchyoC12ApUxWzbxoBSNTTirZW5mNNcvw29VPIEZwJYe
inOOy9qBRXsGwwBWhJKa00XW3Tpq0v0HEoDCh5TUFo6vFtlfSomi8vgB7JtOaHFO
sY7YVbxu3p0YL+Tvxa7lyfz9lqMsww2Cfwod5tkEEP95AxuxR9aYOk8h9SrXriY7
VMXM4C9+HjVxHsODLFGuxca8I2OUWPGAJUiqA5ltdMFsaN903aftfug8b3P4N13D
S2OFCeLxd1/WGEBMZBahSJJ0TWcZg9/Fs++kwcpDgo+RaGtBUCzNm1GWsb95Jwy6
OFutbimPwmuLOKzKdBIKrPdgmNTeYJj12t+V2nKnKx142p7oiWAjnA/1ullgdKJ2
DvKOEb1nVZCcDZ7ArEA3SoOg1OQ4I/wM90pdTIGs+FZUcQUe+dT3irC5vKN08l5O
qqSFYeZZQ2LhyrE0Tz2tG+as/4OVADKgGk9KxqsuEV95O0ljzfJzRXvl5y4TwK8V
a7aT+2DjYF+WQYS4EynbEwfM/akhN0TsYdL+K9Dgh5/SVhx0uN5hWlPXmh+qlg/x
N/KWEX0JyUez61cuPKh5JFl/INRUwqQnk8r9M9zgZMXF90vkhXUce+SoDiebgOj0
GXaStP3bsHPWQONyKFCqzmzHuBK2OVO7YzybZFOVqTemcsdhl51rv2DMzMeFjWwz
Ky4K6DCen1cwycE7gZ39jtzQIt7N7JoNyDxsfZu548rRQbaNXlkzNh+6neyrJO2X
MJE2bKI4/5DH9pKV/6po3oDWADYSjfji5QsdugV6WrZjMUeThqXl/iXtSMY8T+/d
EdCOBvHA0h8sMLCe0N8VBtH8F0ooYbVNb3KUtYRw9HCliY7GzwOkgDPRXl8Oa0nj
F8EQWT0/PRI0mzZYoX8RqepFoB9aHGNCSuEM1w1w4MshHjL/pQZytfjD6aNSrZlI
7gMOqTP4YimSkYA7uowayLS5NOFGwcEOPUz0I9WdBEOwgq+z4kJPYNqVz91xbjDm
+LDjJ3byJfubqVLrWme5nhZ36PC8HtR8Qc69KAdbTi13VsH6w5AapgDhJAktHqrM
0d8Cbkb3wk4FJqoY5Iq1xSSN71Uxv9+aJsUnQpmpuAwMdUce45GVfL7llqMSgU9+
KtpLtNOPBfLJoJhKlftTYzEZFJMAR2dbatVuLAXsNsbYrdKtbK9pcAH5i+e0nCvE
aGEVPiAFaDCUqZ/s7BjNXEhMCWqcIfPZa6afk2jfPVzz8UgcO6NtEXwyi0oEjYg0
6P0yNuSgP+7giD7a9e1jjPLKfMaH/lbiQXRX9nBra4AD7rLnc8x0IlwEaCcHcIib
RX/vjmaQ4nP/1+NHUkqgqSGdqnsRU1oj9VCCGAPYTP+sACS+GOBqaYteYhKNuS6X
ib0ptCPV5EZNsnxl4nSAhjUoffhGoBG1tTejub2ijuItkTMnXf1UWErW7a6ynhK4
xfyePDGQInC+TQcA8DsonwnEnjPAzKLgJReI//U5hb2FLT2xs7xGTlfbS3SGuNP/
nUHLQ+frdr3atsfVUhL3hYGpd+rwdo04ett6lZmg2teIGQHAT9TBDO8DBZZGRK3p
V0I6IWgRyFo8/ONDXz+mELe4jv/tybC7YijvgsW2om9LBoJJ9lvOM9mpK+6QhUFX
aIQ3UsAQmEl3WtrYhldLiURAE5jJHPDrz0FtyllcAz1AnwhywqmkOtfT50QYwENW
+baTdPRYt5kHGwuNEDBUPiJeNeFXE+j+r8qDLwBOqdUgIFD268ircteQFfbONcvB
Szu9XgD+PquI+GiRuuigBumndcAwK9XpShbtRQjqtLdw19fskyWqnYAwwgTO3j5f
unVYH45+bdxswmn9JBYM1fyjDk+OOwBsj8akkG/xWo7xEyqaVErlC49PiVC4Td30
wpjml470cKAHUKfNHlCSwlu1cWyswdrQMMG4Saqc/P9vN8DGrmeeb6OpeFwE6yT6
4d6XLiYAfCbFo8luAVFHf3GEfY8LyVBE2dosFKhGwK6ofar+1DPfMpNveRvXn3+D
oWRNT5q+xU98YJ7bBIHYFuJOqKXe3erC/tP6DpYUjuspsm7G6DjtKEbeFeFU+nDQ
SVFVr9K8YNZed/dYXTIBPZicTK6ijjl9YM2HSnMMad0PzU5T32/4mD99THpIq2xZ
w1BxWb4tEnNoheoavERJwKW3LNI9/1Kg8yQLSN8hxj0H4PJj8rcoM+jA9g5qAp0T
QyaQ0go8A8qw77dT9OVw2mlJQgXzTjuB9bwravzmY4kfb9RPdMUO0+oWq99b1fgm
4lHCM8h3ANBA3qG21020Ppuw8z4jhFI6rncbxtSaqspPF/Nur5TBjvSAEFolw67n
7DgWbexr3QxmsI5/1eCVoXSbPVuRymWA9DU1/30SmfpYl5N/ryc/rKiLfEi9YXku
JOy2tF2SRmV9FaNMPr5n62f400gXZErP9SWseysRbbX040NrEoaH6aZRRxt0orYd
w3KF1+fvzUyeVI4O4w4dVc64pYk+nBhd0sIAprT9ut33yb6/FS1fWuRKxoqs3w5L
HfwxusBCfOYNUKpUjDwposgx4SE6kMBse+GB5t2G2HOJPNAVh7xyZQDa9ItRlc9z
Og09l21JNKjX8WHHshumueUMTji/2sy8NfuNbP5GfB8W5PpdVRyjJdyAuEmdPIvQ
x3C+oLYoMzxd1omLy50PgxaaEfFzR6rLfDGl+Rvlee2oVVc84LnJUw9rKt8AqhQV
D3wcg47JP/vYFrPYJzOfq1tElaRA4bO0/y+4gB/8tvk8dTzlETv3zQeceZodlQVA
m65klXiYJxXxNrLSbvMgvdxVOfJd0Sidz14uNqrJi7IaliZdF7i3iKvKqNjbAQLg
JoXMOvvzHVwS3u2G2yJYRKBUphPv9PmitSmgsAKABS0q3Jto7Lc0/5fw/ETo0yWs
+GCdaYmXQ2oRD61QYDWdjERiHfpBF/U3wzdowGAfQU/U/3Lb0Ta8BQb/FI/Cs6VI
e0MNH2Gxynthq+TwoW5hjrQ61I4OWmwqb3G8J+RVbAh8KZsoC0DO4ZsH10A4NCEi
5pPOp1BR1yIFeBOSg06s3hsJVB1viUXScjpwhDQFbwS2YK8aLM6lNfTWZRUw20Je
AwQZpW9kwjZE0uqbViVnttGxbQn6zP9A1QxEebVv0riT9HKVwgTEYlK6R+eKbOtX
Ua6xmqNfW9oGAvCqnhw1RXpYVabs1CxMishiIB2rgPzMw2xmXldNVpt3ORarVEN6
T+wRik5p/Frzp/TIiazTcluKM57RBEJQXeXwWtzX19fXl/L/NyLc1+BrQP6D0Uw2
vQvDhrVkJFdYNlvqmxpiH0hpJCx7Wwn+ndxpLyD5U4Wxl5fVVyVnhldFmIIakHUM
uG53qh7cA693bzCVgV2zdGhAcRTcu2yke/4JlcR++oi366vlfwPcQfmFt72QVS5Z
CRhWoXeH/Gb59H7eL/lC0TW85Y8VnFrjrjvUH/jjRcgtXbuRHltWBtRzBLdBLzd2
IBa4fjFTtD6O9Kd6/IJkzsykbojm4imWCvaHgB/3YVAZixx/htGhwf01vweZjT7D
OYg+pFWvggJlqDGEKZ0iJXZU77jqjYr3r4+FgRZXgfMAiwWfRwar5i67MDIenwFN
9L3fqro7zqKhMBOWdIFMGEyXV07h/9sMRPrbgzZuSUzPI5VhwhL/iAxOlef7EPwv
m9oT6gw2zy6EbBSkRJZOGIu1F1HU8mILFY3zYog61/uYGr5DqXWmmMq/H2y9p0w1
1Gu0Mrz2uSsqrwMVbRqKF0FRVeXfrs28PCRRP62uQAnBKcqWHtvrB6BgrwmdbTET
HOpQHICuJ8dqHKizS4cfctEwV4XF806YAhM4isyJIgc2huqYo4d4x/bcsGTs149I
tarGlOBh0YDHK7anAa8rhAO2aJDQ8NbW5LRLQSFI7Uji1HR4ltlZWUeXFqOwl1br
a9SbDUX4+385e6wKwfE29ujlMCnDoekUnoPBZlhE9saH9L+kt/c9koHgplJYbhtk
t1CU5ODWx2S9jAWi0PFZKXs9kh6sQzHRgibraSTfBIXDxTTLxaFa9Ms4LFK6Cpsc
dLU6FgZhYsWCPCrv7SdvvFCxjTB7CKieW5en2u2/quGowUtyGW0AlIXOv462+oHS
2JauM4bw8AcsIlhgpSjwPlMq1a7Cz2DKgJioQnueHBik+imD2xsaH+YYfHCka4Cg
kWP6C2+LaoEeIYipg4TBtLlNNVLSUofIrSAkMloMKkW2WQFAAywrVS+hhUoyY9Fj
mxLja6pgutx3b4Ld+x2rPsH+MEpDLFqSoT7NW71ahrRG/YMwMUQ2zQFZUYukpOzd
FiTigFhLenp0VmsNQfK6HYpXhMG0ZXr4Y+JJc9c76l6YFpbExZyFtpDwmnNZMToc
+t7rvdFY4KzHvfQMb55LpI44GEQH1WFDLSQ7cIWtOunOC82z16Y/d1m0JHby0OGD
aiSxSOmPax/gN6jJD20Kt8KadwuFksJrFp8A58EilgU9gCXsbXi3XnC95WDiDRQt
2u7+fr9D5Yhdc8aYYiG04Yv15I1mKgHqrs6s/hogo17m8Sz+ynu7dJYWK8oHjEUG
7IjR89tDBdoHuovxNXruvXBX7kO0ENzjHKaJSlPxdHXGh7/+U4l2eZ55f8g39O8F
uDMXNe0Of9FpXriSAm/vB837cH/MAqNM9vE2pL4osDUOn38yGSngkSgimwh8bIEy
NSQe+qb2MT6hbUmoXwnzacRJgLxvkAhxx0nnWXdToIwxaNqW0pQntEWVzSO6Sy2A
xI4QBml0veYLCb+F+qsSk3jM4ZUbu9vVpu+hOzFKPoeIB2cT9eQOrU0xXjmWATnD
Xn7ZZHM5IWebu99jztxEkyEfxGOvgBIkR+fjhC18Ual436beB+wxDywg38N9EwC0
6TfoooOODcqr7id6UG3daViPkKYhLTve1bu5oS38KhA1/ykC9bEHwBaEfF/tAv9h
8lyLyecSVj0+snwujsK8KNPmMR8gAygJRbSiF/S+LcJH6NuoSN8GDX+wGppdZeHa
+33uodGucNCPdw08PmbF2yOEQnHTylZuus0dMnD2eU6vSwS8IZ8BoLD/CTgs+sFl
OIRNBhp0s9UpAgjTdIJ9TADuP3SHYVDpLA2H90aCy047rsC8GasvarQmHsNrzu5B
fcZoqN5yZ8U9ysIbqHS/JhveMES9MSoIc5+ksreNilOJRJqoqEQhqbylEH5VrGb3
hVqqLpzGhoiEd3xCgM3OkAwyQJalrbGMR/a/4JeQD2PKmo1TMVt6u9GpWAV/7jwR
VC2S5MnsCymtIxIlAyROPbmoBV+oh/GWtV73fXmsuCCVxnnZmImVlKPtfq/kGUwu
h3ubTRZ7woIpb3NMezvqrQaMR5/83rq1gZtsaZAt03bdgsa5+3O3kRBHED9J5YiG
EK24ih4sG3cdNUOPsoffS9btm7Yg2Ca0j/ycot/WMUPodWH5Ocor03EpCqHwjHKr
yR/VWG6TxBZ8+hqBedzFO4glQM4326YOl3s+8UlBXKl6barelwAvSmKXcokWM7c9
/VC6vP1wk7zll9uuDF7CIFV+SO0R/9VZzwmuKUz8KBCyVunHQ1Srjg8v+St/fywk
DjVIxpUTMG34z2kwmE49SmdbcW0kioNqzwA6CT25/R88U0Vr4w6760Oeo+Z18a45
AAYpwTHY0qEiC8IiazUV8JkXGK2ofHtwpIfHBeuCdjAdlEF8nEQu+Ib4eMfWy0Kq
8q/eP//UGeRjnhOGW9paMNwU3LEbyf65IZ+ZFfghMf5ybH2Kk9cJ7+CLVGB2IiUF
yu4pYZOOjdYfttfBA13TOpwhgnmXoWtYmwGb8rHswML8+ETqeFUXP5NIk1RSCy88
kukA+f4KgKwQbOkwDiDhRoGTBqj850e9eOF4wPfcR+xTmCty5Gbh43B/W/EtwE5A
TjJxSdxN2gsaENytnVOdk1uby3YMBkXxYeeTrBxHVGRHvJ55fobdQmqDMnWH+/3t
xUGuEEZE+U/q13tKQjzwEU6k51YYZRrMYF08PwEpx1klEaaS00MhlJTDyYkl2vFe
68TgIlNxa0oIfp0KvGPA30HwIw+NclVqL6AttV+mjRvnNvJSA6qzrpzgRhFslNa1
v1GitIVFos+rXbp0sfXUY5iwuiHsIdz4BucceeMDUTSNjcynF+jvyZEV6iLL8TOR
Wa0R3/53ESiDIkMYtOirsyf05C22emQs2EOf7I0Oo9izkbgBhwezaJsS1TMtfOJR
RK56M7pOchjeTA/jyy+SrTWix4pAXx5eWgwthHi/1eJv550RSONOq7uU4AsoZc/M
TN7GH1dB7Sn4kbdqk3TlncU+AIfv7vUtby82LWEDDfdWEwC0/FWIzO/waiDg1XdU
t+6xlnaPJzls05YFNeGtbil6Ecapsn+tYlWWQ8D1703xfdVtDBiPIMUWxRFx91uq
/97U8wNPHVOjHjRI+Rz7yY4RksZjqC1bf06U8A0DhSg6Ifn49rXSB0n47DTbu2K5
gEQxftK9OeSrqOcbWsWnUuxzamYFok72Xk/88leTtYXs1O/FzDa7o3wwwA2RLNUs
PL0g5hx5F4Lwf9gUvQBe0aQyCvV6Ol6qqjsVDrkyBxATmlvnTsH64eFt/MrUyvUL
1Fq5Y+yzljjOMijrePcjv59zMw9j9s1wWm8O5RW1n0BDQ9hXVEu9TrXQBtM2xg0R
2/c57QEWctzpFYaAayTjwQdnjoGo7CIYal3q8dCOa08G2rP6sRQHIBQ8gCi3W+G3
5gu2MIUD4077AVmtpDzXa2mV1CydO8PmC9IiZExYnhfb5i4FvzBFxILIleLmtQMD
H4yX0qUpudUVog7uuYKTwYEfm4yse36ZYBSEXIEiRguSO84w/R9yqKyGxrQvxFTk
jtGHc1o5Zdkqd8fj2YKN/s8r04+456+FbG5knFvW5EP+RDI+Z1kzWtY+gLcPAUpb
ebPNX4SOBLDE7lEYwDuigL8xyCNMyaseT+t5JzpGOBlALgZnGiUtTpc5u4NuS+nx
kpmoa500JLhsJOQHVjr+Vv2aN8a0BMmkLClpafjmlcUrcLF6Sw7/Lz8UlNl5H7vS
4UZWMOvOqd2HNLKKtPV9wMv13eZqkwvzUD6HAflEtUh+7r4zyg265GgwY5iL9AT5
9ZoGsBUoJk2/PGoQ1Wd13MlF61WAWa8QerqrZIEYs5a9OFLV+2lcpVDurJpbjK3u
RVdGf59O227DhbcF2mHEryEgbFKbmgqp2u2YtvWPjh+bSImq5tq60Vxz8MxzW2TE
b2sbGMxSrhvbMU3h9Rb8+e2VZjf+VRHKFAsb5f+voWoLxGJ6hquLb3PJLcL3R1vJ
EW9306vdeU32bl3oXwoO+SkZv+PZv0uWuQa4LxKalYYn9TbGNAqINnkZhNRuKtDp
ZRhRy6hK6LOepLR3usLeZ6uW5/ZHH34HTdgywhtWIk4VGrykZkmObMARiQd3asbD
80hU5uwK8LVgwDa47iTUj7/FDFzzlYgkgn96/QL44DsplyT6b0tLkoo4iCVwNIbj
RuFyt8H1VJEOA+zEa5/lnqG4JhQ17F9YDqMmmxtaY9R48LoxhpmUd/qCV6tyuxTZ
jPWRkH/Zs7VFmxJTqHvwyXsVpSjYuWbgB1wlB6WYrwSh4P0Qct8NkNkw0oWC9CO1
A9ARK2rocP9uBRLsNgSCCFQJilCCBsvvG4nq2JSirIJ2zQtodwJX//2lBiu+SpWb
fPkwlEXWt9KLEOb3lGM+jrZXQGsDvWcvMwcxxaI0v65IVdVU1tD7pAg5HCnVsWGe
xZiy9dybbziniX2TNfm8+MNVH8IPrsisUy0YN0fr2bcVd4VDshe75OV5JqX6BsQ8
9xH0Qa+e8IH1vJArOg19W6sdBvTXP03YpUXx96rkoiRql4I9ju9o+MwyoM0+IFQB
yFMPCGMi1D1x262koB6SzOtVP7oUT9dRBMZz2vo8ZKKXFhn2uTaaTRd1dObzVILA
1Jy+NYSwS4A4LhEUNDn1H907m/85mMPWMuxtQELrihpSVYwBRPbaq9LanDF97NY+
fsq2hisca6zwXui6wtIXqdN2gTRJXblPKaENJ+tR9x7a2da5teHpLUKb9qOg1CtU
BCM8JEcxnzsI6S44nSq9gj9Fo++jcpQPkzmHojK8g22m171+r9+oPT1n/4XOCQG7
9pXt5Q+Qy6t5c6qS05rp5nhGSc3MsEIdgBRy5ExwlzknTlp1AvXBPmVyGvfotjpn
SLD0wanz4xlu+oX0flNqMaObygqXchkQBxC5F2O+Y5wrsGsACMp6WR3z3Vi/8bC8
+QkJKomxmgN0DF4XphAS1fJGb1ycEx/UzW/UmdbJYfvJUZ6fXnw1BabE2cEunuFh
z8zuRorLohWHKmxYlOtDnjr9wIcUFNIR8nQOdyoykk8wYzPXd+ay23vqMVDkFS/g
MDoMNEZfhlij9x1Fu79Rhee2SHahNWW9nW3tu9OjiSXvrmMFd8CCGnkr61dBy///
c9ZrSHIbQPwyrcA+P9xGU2fISSZFRO+qLZU2q4dknULO/vMLw642h9a+dUq/zpd3
I/t2eySoN8j+Jg01bC3jgZXI6o/bn9FSsf6nX31mucvX9x7r2IdHoY5IXsHzAkYP
YFwECg7o9QXXp4u1+tFraiJvg9lj0/0eVW92yfpNvy6Npov5B0O4R0B/GBRovk3g
i1KLxMkAiybMDVMnuP77csEYjq7EfPHtKgTor75WBPmV/TEvlFlOh51ZM3z8j+V4
ttWyBD5rFfH302Kp9GJ7vIN2NJOS5crPpGkMD/w9iWM0VOqy74y+ZToYKGiN+crF
NB9YfvNSnk4/E3s+GcsJlLZYXWt1dn3flEr+vACjU5pcGZwQF2BuwI9wmZn+55ph
csEZ6ZsNUrdicuf+2kCWqsSw9KX/zKkqDSIunBb82xYlQJbDehvohjkJJ28w/Y5T
iex1mhvX7Dr86PGeb6B1UdLU5jtk1OiVhe6mzlQo/8DYVkJHi8/GLiB1K8GtU5a3
jp9byG8QlGLV4DTdKK0RMh6q7KNS7i+h+hWhL6iEaeoRFtO13G4q8QQFg7xeM3Wv
VeC8FqP+pCnvhcxK5SHB4x7ZPE2XzMWQzm4tKOG7ipBcGXpRx9FfNEAdPJS7hL5a
m6aniIFFYuypBgGBDsx36E7x1dM97hGhvU0Eq1LkqKdZZ484r9/sECPdcc1tgC+v
znJFcC/anLyODcGiV+jGPzycw/FPHt/hqGOdfJfY2pnVJ0hpmkG6cAMaYAJ5wzwn
BkGraNq5vDznsHx4AnIjJy2XUxizUV1/oDk7lewY3Y4Dyex/8LqL/pGcDAU2TLbT
+EuewGrXEwg5cpPeGHoxu4DKxOqyEKCqe+WQFZDbC4l8vnJSFqAmQlAnHRwsNaoA
uPIlA8BNSF4ZvyeGeo1v972caqH4vzm2JLtRxkfho/OfwN/gOedbx8Iy1sEYHdF5
Ag1Tsp6MbRdAFBCVQK99uEovH6EVfRYHsvg48GBKkKrIDZrPfyGJm6kluvFrp29Z
NDImsrSASnvIVvbEM0AvrmF4/h3X7xyXUEB5hPQLEiNEvXw60vCp6pUU3do68dah
OYVj+imEittleYPynY35rukMLafTD8RYEmebB/JDo16dGRgotYELP/44J15ZJEAQ
2m3RpFua+vEXhFvpUN8VAEp+3waTCVJ50tkjN/sNrA/dK1/p/dT5fez+tNYxRxkm
B9x09X8GtGVjBxs1UwOtaebtpHiXKwnHgYoSoOwfB/hcmyncyO0MvFaDgYN513Pv
jDz7wsR88BNYAqZ8Lim0rByplL20dw5WdtOeKp9aHLw4+eZayr5QSakOB0SOqyqj
4LTQwU+fDfL+8ZmanAgBXxhqVivgR6rPMZQlAVdcF0isvl1K2TWULUJqiVxxpt0s
vjjFILoHoyoK748G5+g2aK6w3xURz0KV6lqk8e6m375oCbEz/0j2IbB9+NPcxgjl
KdUbUp4P7laGByb5j5miBYujf52qrUJcegXh/TdZx+875pVaiDsXIbEI6unLbRmL
goEuCt4cnUCQcBDk9p6XuFKf+Q2yNI4ds2LGw4CHNFPGNHvQu2pwrzQFGhdhg3+m
bsLAIH1BJG2zN0zaRbRDbRVMk6UOAKO9W5hjib+fAn5PeUPuuGH401iF202MvIvd
xauaZ2he3KF31x4O6MhQUa6pA3v/gFr67ohV4Mi6/JbKSiQuDik5nTdPnDZQ0Upz
XVcKoc+59bfSDiRFGjPltVM1kKzb4hnLwPfdo3kQ1cCyRVUzhuvRwW6f95kqhCQu
7gYhP+xRI0drAI8IG75K/NOodg84ssWPMlab8p070xlSZybIGIayR2NCUSqfP6mM
VqI+29arxiAjAL/vDZ57f1DJCeG4vXFv37AxWkfeagM13Cl3ngs/BzO1hVlbUh70
IEgdrCeGuZqFo0VDuj9VsHJdIYvneVW1yHrfF7bmVbg4RO1+9C9a+H+VHLqhsihU
yGFX8Q5efz5sNlElhFxmWiYgFsX5OZ0GGO0cnxzD0xJCrGv8D1pVkTabPrnPVg+m
Z0LUyqZAXiOkq+Me/zw7oybaeyEvNRCWnEd0W+JSvYGvBgEmPpiTl3Eydux2smiw
xJCHRv39Ke1/9Q0q1ebJWRqsXVUTbJrMDeG3nLrcajyM6vr6aleHOx+QlzKjAgZX
DvSydRvK4ao2tm/q3Rc8qotGsd++pmnqjrgZTOUbv1yGKQM73iqaatEU7umgLbVK
/ICE7IDlOIZcn0CbNeh1ux6XAmRTKEDmcU4lVu6Qh22oJMdj1pcdf+OGN31G/vC3
Gn0I2Oj+MImV/pc6260ehyiv+vsrlmmi5DyK9cFy0LJ6z9OGLOItWL7oxEVXEQl3
BgKXoN79mR3sdkZexre0Y4zmRR1zQFhFSvNsbrqrtBFU9R4jzZX5rpF5Boqamr2u
WLaCEIDFCBXU0u3guUF4ojDQIpOv+XoIu8JnVdM14yK68r1WYJROHbde6kaYC381
EhZQOc6F9ndny94X2pv/fOA/VzyluXFuDwzxL83bH9oqYxeBCDzUPbF/Paaz6z3+
XrjRyNcMCWDYXcpSyf+PeDppwhPU2NwmTvM2qR4TV8Dme3zvhtW1kCf/8hWotv4J
ZV51YApdy2ffTAaNat1Q9DvzRBFTV6UwTANuY7ZSdvqJvwJEtxwAWfcbI+pqFUZb
arYpgnQKQeU4Raq61UZZqV/NcRHhJlIbgArSgjUH0SboaqeaTPsju244YwPosh6I
/9HPgr29GtDWyJdCM7DRYtkj/KBo1JvUUc1p6WdD/k2jVMyqwP6Ck5TPUWgYpCAC
Tg+4SpeLXer0f+D7lR7HqmdIXlZktUy/ztYmJJLLC6AZjBYaKQsygfRG4TW0QLc2
b+VqNpgIGygVEWTTS1s2jv7N233UkHFoXlLkaxbhwB+tXim55RljM1TZZ4hnJ4Ob
DDBkRPFvvWGLZ/0t2jdzI6bBW33XFGRkmFAJpGNZs7loXJIjDH9tSvhK6wzyUuR4
gACZNzp6r51N1zrlaDh5YP9tZuLmOUTF2cBGbJJzjPum8FwgIFs6uAG2e82zngbN
fwsVeGveatJvWfWibOn8HN0iUmBO1E73OZZlPw27AK1WmMFq54G2/4MQCpCmxAkR
JivEk1wteqCL+E6XdiUY4MzQ+i5WeU2L0cnS9OSeRgJEgfzIEtkQiBzGu2CTgIk8
F+pOC5jnQMGmxtc2WYN6h4JcFTuMK4vobzxI7miWWYlcgLGOuzkXri8hHEySZRwF
Tv5U2PWOC4RhvLcAvN326qMIalZ4ThDIZnqqL8j0KavZB9LH5pzLc+YLtKHQB/Kd
NV46m+/JEr1BAV4EihpgUlrRLQJeevzKMrUyip0Iaz/Fsun7G+jYCbaWUkfETOV2
77iA0uTPSZVcBpBUC8GNiM9+GsUJXV9up/o8DYKuGJjufuUm+nJbu72+FIBjUhOs
1ZESg1Gy2BQH0gVaF7qMn4ddJ4UAUGydFGgL9dQgzsqpYegnnfg1tWac2LCCOhHq
ZVyYutHOIX5/kQwNCJ9TueJBKMaL8UNBAAZxCVMSNKm1X2BlOa5WdCZcP+aFhfyK
N11RjYvfOGPLFIz+OX+PbqLDGrmH7jXKvx8JW8BQRhmJ8GluJaLJlC6mURi+5o5Y
gizOHvDnENUxeIp4MnMJ1B9hS98nG20oqDL/F6O4RVCn9S69Jy2ez/7134Xw55KP
XmVWmNhW0/QktActvfGlJ/QvsEo0YNhfCyCEzbyUqZxkGVXTrtrN5MCvAp0x1bL5
pejTvyzbdvAAdAuymyIStERJVGcELVjNs6gP2QKdQx+I0j00JOy5bAvOu1ytkNYv
S+ZMN8AWPeBchyhK8a9aR+IVmKXOF6PVGputw5k9O69zcVzn99krbfKSFxHL3dqL
xvvXdxIwQPlNOcTXlwECTNz3dcutE1ERTbQCoN7YBj61dej2qJiqScn15UuE6OTq
yKihz0fKSTY4kBEi/i/QsspJKwJ1mi25sZWkFzKlVzeXlj4D5Yw8uPRUXQmtDdrz
GMUltu1nfQt1IF9qSfDHCdefLv8vEsc5yJg2XMEm/FGzWoIPhwxk0UzICjcD7IMK
J4FGS/WJ1WLB1Xuzotiu8oWuKG1OTMp0GvRsC0XsNO3tXFDxsm1iRY9QNxps4tBb
eSEYS+4hcGpwd/YrdRu1mB3BM+s8RmxLI+crTz0fP1R4/6+mscmSPX7hAC0sew5L
7GzfrPdb2cc2aPtw706/CLvyYXnbJgQakTiTjZMoBCdq3uxUN/0soxyT96Y3DOqK
O7fEwywV0HOUwPZXL2bZVaXrhmTEUphD+aDNA9x0PV3gzCa/jbCzmlY0F0b1HjFX
k9U1pgbIemyceLqawKYwNu69Lye06VDME6rFPCC1gAeBuGERUH5JrdiVMxaCh/Pr
kas3TlVIlDa++2Hz7Ltzv4DXxQyHY0L2PiLEhBWlq3XDY9ts0w2F+CwraKgzl6Rd
/it2qrBUp6I+45Drd6pvAD1tD4L/GuK6//f37r/9i8B/oz5dGogDO4vIqfKYZQ6I
5aY1hC2g2C4VAA5duOEGvGYIAW/w11UJJFHjDish4yHui4ns3LgHQE8/vqrSUjfg
0eziQ5slleUK24NDgOmK7tCNnyBTCN1nuW1eGuNsG8hloY7TQTC7qnaBdWog0kz+
5+dPitrUwALYC/s+3PxNuxucfFRWQNYnTq7oE1YlIfwXwzYER7l70aamIRwPYjsq
N640v+yQeeGL/FpQhBoRQr5mwF1VsFTIzgVa5Eu7q5AmbUEHb0u8X9EQffO8HBA9
UTOqWDv9yumGuXjE678JRNvgbgM67v+6Cv77rJ6HJFGZXfCRa1oiIGUUkUopSI4V
ZMxf6kW2KtiJYivj3olH/aLAWttTsXiNHgQUqqTDx6wC3ZrHAObMei3vQkmzs4Hv
5v0qKiWhMW2LmsLry7hBu625+P86QwduMkw6PMzVTelJgxZaxXrzOkuz4e+DxHMH
5epfC7bkmyw9o5rg7T+y6aDmCpmQqSR7FYTxM3LBoGOnJzamqtRE7IGWg4myvuB5
5R2gCI7Do/qISIVhfjC9ELwggy3/Arz1mm0y77BLK7DJIf1u2mWwnnP67l6/TPqn
jseHaCYjVESsFFrAOSpArBvbz7tmBBGvB8Q9vLGOyVDxSgrnaITRFd/oNuqsfa2C
pYGUTQzx5B1U6Oug5HooIuofKHHUXggpezzysuKvgyq32UhRc1zQxSBrBfprLBpq
BGms8ncUnyAb9DdgcV583MDXeFK7VH/6aSws3fa/YnPqvYvENj2DbsSk4hhf1G7Y
jLDjtZ+w6jsxSP0iK6Vn5cRU5MVxCZ16ApeY1177nsDhwCrT7AZnMaBoB2bNnsxv
Cka2Tj5qMDXVU94BO3RNB13UXmEiZ6fzB1/DeX10MBbXkxl0MNjo3+3wj0ORjLjU
vlslG0nCPissRnhEDuL62vpONvi/96y18dEKqhCMN7+w1tXKWqlXXoQMSLd0t4nU
uAKqIwxWHZvUTW2YOk+2zeJFdQ+CbUeH5IOcTzO26VX9ar2g1agkDyXuNtQxalJJ
V6LGYGhiv7CbMdECuszbHhZOXsRD6sQp4PQRdGOcBLuABjXMzf7t57T2EubTtrFn
xpgpJBMJEeeSZJWj/KQw2a8V7qkxvh0+1HEDio3RQoKcnJGSDEsybl48l8W3J1vQ
aJ+w67MOMb+pvo6ZLaSGXDQOjjjzOJfgmP7M3uZAkxFpAzXooNkY+dT2njlRgypx
N9/r9z1Trqf35RfKZgaCSKuG4gI3hujBpYZ2UjEKJ53f5bRVdiqNLhiwGU3hnAdr
cWb95ReL1Ug9VTKVkI2IwcZ26NsSoFXi9K2hAOxxwq4xEcOb1uZYDrkdpYR0EwQs
L6WQZ1qoEOfcoUBRqkLghj20rLYopMJAJ7znWnKUUZbzGJvhjzCHttG661MIuFWx
/4wfsfeh3def8ilsCZN1biLrMeZpgo21EWvBRhRx+xt/pqSRMaCTVQCfizq5iUxT
fvM3YaZT9oeg5OUV5M/9b6GhDUXQqcOLQKojFnSPHYaEMiPu9JJU8eiouNIQQNQB
s4fKn2l6CAEmTIpUf+2iqQ8d6mBMG20W2Txpos2S6Q13iJbFmscZB+WzGwq5QuIZ
pDoLRGGl1JlWNW8i7UdmKNvstpCu6NxcNFE7Q9jkRxjPk2F4/GkzAI0NoEvRj8IX
l5icGipLuq/RIlx8HNBCxy6FLsgqgYzRxooaNIpd3QO3HaCJOgD/0v+zGtVIOw5b
Quu2B/rtOQDXjslmu5zmP+ND+le/BDK2PsMBGKRDEwqIulu0M6FAOXv33I8Dy79D
XNjcdnGG0iUrnRbgGdL/R2ssSzbyJkNYhaoyD0YqGg//MPB6DdteVw7pQ7E2+wPC
hyfKeA8Ivyvxd3PRMddElP1FK9j/7QIr7h62Qq8HoVPuQiHU4jo4p4q70ER3j1Pg
5pgV94FrZ4qMaO5R7L6E70eiq57VhFUFNn6DCZsEe3AJplJKzZtnT/82jNsa7DvN
o0zP4ruuAxT8RpycdHVRxYh9otuXkkDCoV/SXSWSLShXozi5M2d+K1ldZ/PemghY
pa5MpbCP79q11W9ClIiOiLIvhDTq2NqnLmTg7SXqXh0FZNEhD2MhPRUnSglfuJ8y
BfvTbs4yYjr5JpvqFX27dTtMskVqiYGccVYuJNnNzoKTFPEzaS/pyhHnQKYr+0yD
OwYK7K5lsFEj5eWYDwbp/yPaIBcD6LrzUa/L3RQZpegY+PZdvamsNmIvmueDhi9w
CLRuAWNSU41ZkeBNclQqJWBqZl853eEErO/Qkw3oxg7sSl0J3BrVLNsijt4eTMTT
ldsIK0bsohesZJeYUNOOjB0kJZfLP6OJ8YLx+vhoqUQI22MYXOCIPLZ+Cm61rS+i
xvoF9kgC6NREkitJNQaUryUNDDh+FH6yaph/CTQuq4yuqAigBwA9dM+tx1aQhVsa
R0Cb2XIJGTdwBwofUPbKHz1wqFqAqiPsoIDUI8S1MD2tj740nxigL9LGP/rO4LPY
l64Uv7o65Sd0O+E+yB3pdi9idvAeP44EIkKm1RdRq7lvLUWxo9GiIPLzvOXqIpNZ
3NRqvcGwGnWG91FOE9VhACL3L652V/AHXyZ+wU0ZQ/4ucMuCGCuJV7ai8EhugSV2
6WH4sDpAwjbhd4FqnWfqFcHF2ZFjyasa0+X/uTYBBpGadJC5M7CdI0QlclFg0Gli
/HWc9HeNpP9VQ+SxgCWpaw+TivgQGuKjw1isCO/MsjCi4LvbQjQ2YvSnWlxjcwMA
hFjoyskU3VUzjfGYv3Sgh06HRoQW9EvGLPCXZKsctlUZdJXGSgk43fHHfAT6mn2e
MgEvo9tjGAr66in0n9Vu0bHOEuj7nXrXkLzbZ0/Y0Xmg8vPjlQ7J4V3AahyOhe1A
7j+3nWQ65ruBF3QUwJPxbNOUWl7CN7LMqXk2dLDAiRgEV7HnYXR8nv1mlZOrwSIz
hdYyugxwUl1hhgE4BOjrPdMbb+0mMK3XdhsfwF+HOwRhMMRUaN5/HeXQxRq4GEzw
At9nQHlySMoTyUYx5I7GFvUq7OxdBEMgutFCELH3Np9Gly7hyt8v0pu39RpxGQBe
g6BJW9hilj9kqYPe10expAxpjLnf+YYhimfS14lKIPYIRGX+sX2CANxJYIMLe+eg
78sKCfqGv15UD/9UlUSUmNhXaVRDYSLgqtZAy9ANxxczveTTpBbKvugW3D+fPHxk
MbXqtiUGRSOQs6Iur3+5oEmZBuDb5Ghiva3XKllA35Mg+oASU/F/s2SJPA2fjBa8
jtqIFy4aDUhTOIAII2XPIOomd2F+9CXmD0UYSfpf6M6+ZCufx2NuAVpYHKwjPpwV
Ohwigf/vC2Gfcs74a5fJZBhdI5NAIxi2kP5w1566cDDj+wLh1LPcoqmV6GkQ9n89
b6eHcpAl0mJxMjI/aEn7G06nw4Lne5x0jloW3CUYkQfX7kFWwwoLtROmjOkQe/h5
usnXtRXzaKhH62320qTHYfMt4k68GJYdUajlx7FTOn9La+TkmPsZTOWOGDqcCFgZ
AdwcgmcsByFe5oH1oiPPlqsvOwe31kY4DEIWF73BH650ZWz5Mp0t91/6+npN9OlP
IYSmxhwFxJEdlFmgvSdVVBAqcUpJWqXsiGJw6E5fI8VdNViubqC0UcFNsCZVJV8C
+bV7DDTU/FAyEobm6ShW1jxX8HCMj1Qow5qX7eprqDdYic1OBO16jZ+K64RICDFO
AIBxyPpPmptJHKHgpInJ5M7gj/HX2cQ5n/crkTULNf1JKNsouYhQybOgGKHekJGF
QL40ntNaQVsY7qcDG0l4uKR6cDfalaTOeoPt61gF17g1JH6m6IXM45oEH4idjxG6
Zm++LxvwcytkeU4q6ZpQ9OQGqwQ6w7s18uv7DWaPP0661ZplSRat8KClnme8r1VI
iG7mfLWCUeHo/+Ppo8jCck/3JANouyxPfQLxG1XxFr6+7GaUZh2dI68RFbMtHuXy
D6//CGh2HcnIXjYXKW3V80FHTP5L5VfQUoIR6gvzN6HZK6zMH4pr0EbIbXr9blnt
5rEE1Rv6MhRBnYRi/k4S0qs80usOLNcGkJkE+Ndq5aV1qgi3Py45mnf/e7IxAN/S
hMhjiD9eoEp8/IKVX+FzQHGNdfut+4sVuLh+diu2TSHfrciM+GbEbf2R8Lhm4syw
hLpo3cc4Qoll3Y0L2og0fzO0kXSHN0nZ5XZco+QpdIrEl6aPt38Bz4DdGNx8tnjC
0zcWUcB+Y+zbpw0yg2QFEhr4no+w7rVzLT6y/5klhbatOymVVeBO+D9UHP2iEZ/e
3zUdrFSV1zPeCYX0VL6L0bpcL+xEBemsVDy8ijFiFQTxPdQM1XTxFa2EAG3nQ4al
hJAxWx0n2w3lqsg4ZDQCwsreBpOzudcCrVK5EWL6MtDVeMvJO7nDOwS4GYsmzdMi
X7NaAzyNjE7u5SDz51EjUjsiqZ2ls+rr8SVrpYVCZJO7RwB8NLGe4tmGbPrZalDN
ZZRqn9AswaZWwxaEBnyWYTfbQgBgqjvc8iAKR9L05xA4R7oyORIMDLdjdMX54H8e
NAJn2oxawniAYYvz67zNWI3C6epbCmwFTRymtd8gmutOQmMuoHiwNQ4bmvWQ/LCU
Z9igKpiYp9KhvhJr1YoK8l7X/nqwUHbsB4cedPWtcONeIhG17oKGjARC4zqBHEY2
xNdAVkq9Dj5O8a5kUYuYesYWMisrxA1Awgk0vszm1oHKUHUmG61HSzsIBFI1ykGx
FI4lk103n8dbDFR/dqdTBq/9HrfEBTw/IAdpTzZ4d3bqD5aoAbkUUNdCGC9I+ynC
vuHf0mKUBCovxJ5d7/2RmRilMkXcgElJqAfEESkCUKODwBpRegBPdWtHQibIZd6E
UUlCiloHzFXhDAObYHO7oo/fjlw2TUOCFGzUUoSJsw/d607gyBY/TotAJl1GekRt
ZNeFA+QZBGdDD0A2h6epLxdxsGcEtddpG9b0SWFmqpE5XMW7CYgJ7/vXrjAp3nlF
giWXvQPAUWlfre+o/FQpEoOD+bmSBGOMx1RbYrY5Bu9UZlNK2spT7g/ifod8AuzM
W+XIsbbLAbFD2HkEWJVMUe928hk9sA8PRLGdSNT+w1irip/ncPTzb14y4QSNx6du
NsNcPZeXzk4G6qOtPHhTO4LPUlGqjYkN/yR+hSEhHXxOhBVbiXJoemDVpcVeurcP
ZF9b3WltXMInuakmZ+cgzyPgGaOwFIvpzYPW0I3wXI5vuVJ0s8ro67Yg6OPlg7Yt
y+v9lpqC9F/SGcJdFALzQtQ6UTcARpy+TcQahitnJgIw31kzI75M5UH2XOpDT8Dp
KEsCjzQCjRMznecDuqf6eNWwohPYnUNFSa0CSw6TRYPg4I/RLm8N+8ymnUsrEe7l
cnndlvOQLFHPCvQ40MTr52RlXElP8Ltpqw58vg9OXcaHZ/bbVLoskDnxep/TJNy4
Dv18ef6Bj5nPHahkeSOGmUU7KISjJIILxZy9O4LBG6zpfF3Y1LXgoZouEAz5Oc+f
T2chcqDl4oKD3aDYEncu7OPn9zLQJnPwOMboYNZ2l1SvyCx0sac8xIuS9S74Zfca
lwdJl+G+w1J275764dB8ZqGMLW8O1/SQt/I4KIZHVpOCqY4ABjlvozcRJ1TDYbej
01zmBFxzcBjtYd6AxfidkD3YkQ7ZeYzsD3S1D47S4YZofSj69PhDbIkXJjaVfxYS
g3iLRmL28m+bUFxSflQZXCdtD77xMG+mSsRUOvY6RIgbZk6zel6cxls+CCybSSGF
eIO+XwsD6g/FkChgiPS5qh2qufSvlLX+6cNDjptrOV9RzDG9nhT/jA6ZqpRncYAG
4+1sSYnERdeBdBdAPZOtqRGCms4RODyoE1I1NG3r50TDYs5znlShYsqkSRq47u4E
gWWBxzjob67yAY7wFP15BTlHl9nCtfzusTeKAWPxLTJ0JyFfFHlC0zSEWhY86n/d
fMsxRV4OLMpwkEfQNJ5bwikrpGV+FDZQMqrOE6UiBI0ikBLL2MWiTAdpBXPRae+G
Ef6KbheT+17BChW73rdMdcc3RFNaFoaEdO5BuL7145+JaPRIdr1Vy3c4C8LzfD/7
Yn/WSWeG1iMGZ44DqpYoInrPIH8NrP0zNuWkUnDiE0hxiOyEMZ5bOvwpYzetGdFw
iEBheqqXIScfmQ9Ause7g91j27cHmfYyU+wXgsJ9lbQ57LcuoI6ryCwE1Tme3oat
mDZ5AQ99H+mtvLty9e4RpoZtD3bvOhkhf64E3WJRV7s/PkzrZY4n4rqgMKiRBxaI
8jFBZsFX4OQeFdX8+znrCujVTO+i/QiaUIdCyaqjY8MrauvtfEgXJRBiwL/E4GsN
RZilGCqFa/GDyGqpnoUmnqd69ucKPzUMmfj01b8LG+4cs78TEIzwq7NLzRUBikWd
z+QfkLdk7mebhFSgi2F/I7xIna4IyAtgWo5BgfzPTILgwjWsfzAYL2ffdBHhvzgo
x7ihEFnTEaTiG0f6icGL12NPzYUqaxkbHGEkm+7u0i0TDgWi0eIk9zpvJaSc9kqz
zuz30Y60HmkcZJj9TVSWw7hYj1MWiVPogIPq2XSLLKRvR0eS7JGmEq10Mgpktx6z
HV82l4hvb9t4c5afabdtviFjD1smKEc74OpPwg5Zf8hhVvHhXrAJovYvwBuly3lJ
E46lgnU9Br7JhqULll8+0UaLSDTd/xNNYFRH0dbD/dPTdcrRQJkPTWkf+xeXi3np
pmojKNlVvSUFPgttuQapYZgkS2wb0hpiHox8OJzZ0e0Cmt4weThaqKar48SyXWIK
Gz4JAxg2U8SED58PqvoSWn2xyFVA6/RMfGp39+P09HbsF1L+BJ09CH0DStEB+HuH
mCmzVtbrXlm8J7R04a7LXZjItAe/VkiQYATEX04MhxPiZPOibOegWLH781ORY07p
8RYndYczt3pPrKjxI3ZwmFVqZxXdtcPMEdiKfPSizNzgP08bLQx2dNGR0ZmQkkEa
n94YQIJ50tgNKoZNdM8+bT8y4u7Jbw8IPpCqTSQhUFeU0VVq++4fZMRrWkcpCERN
E6KUTssye/pgekPmu+oa7RPTXxkrZyKYvVXAQgJUTfgKxW6tHW/NfgSFuW7CF1sZ
Xzh0kiWTY9WJt5Lr/KAYj9YnEGTCi6HgLoQ3p+OYKhdbNp/fjvvXTy/68FBkzJzd
2WU6CFbDg9JZfOtXCqnYdDRbGWkvRlOjsEGEs4mgENDYD6J8Xm+/3oD3KkdoqCit
w+yJHS8M3kd8bAm1ggMQGJ4mK2ROlMDt4dt7Xe/dF56/lJiNVABt7KimuuwKk87G
7loSvWpU32xmjqilGxuvx0KK3azU9odnSFDucKZ/d24sKNidNtXZ/wQeCwua0HAD
Unmv95/j3Fh749qmkwYCFsIgvLr0bwJ0KnBjL0y9Mq4bIFzJrMNXdwAQ6mSqnURy
zibv/cOn79NLFNAxdW7X/BPceML29RpXzcQgTVj0hNuBDdy+3GNKEBAo1e1OSmzR
HPVxHXq/dGIEKEKajTBZ10ov+/XAdINkqfR/FosMH8tk5mo5/5U2C+PgcvJOHAIX
h9cHLH/pVX9avuv+FcvJXozaRzKg0Q+koJtGinyGmlHRehNoDZBybwOju80GF5ML
Y/EDBQBbaWUPxDJ/oCNSeMTm4PBnW9qvoVTodxLVkk0ZV88XKK8+Z1m3CncHcQZY
agr/VsU3VZZh5Fc3khq6oa7ddG8XzykQVXrkuRN/I/9SxrO7vRnaZrtg57pz8IaV
C3SNDhobOFFiFP2TJdLhDHtes+yl2Smmm4n4natMkscr7djFe2j3DDccgrJDC8Re
vwCknOsGreRe4kPD7glVwvElCqoe5HVSFhZlnzdKgXXqRi/9onI/8mRonNoBanCY
4c4+LV2cN2FXN5CyxA6m8P34D24KWf7xB3qOQQiK3rvv9zQUuQhVTyeltMIUTkNZ
cSMYCAHheLRxuXHuo6nG7U7DO9VAu5bnjQdLl0B2JzjyfqyiBjdPIrC30Lo/zU+H
ayoxdw1Xvi2I5YGpPl8k4WAtcqF5lcRodQHEg0rjpce6MFtigvcka3eh5bcn4AhG
WurWgxAlejAPYARydgu/dbrcPohkKhznWOSF1/rZbKLCYWrtlTYnDaDDW3ooxfQk
whYZfrBq6UBRfEEQz8aE04crgVBYnLncsmc/MaSk+9mrRTbC7f+uKL1uLH3182Fd
UF2qh9LCEBDlvG6KGEhAxraIJHbIPD8UCdVV89bqxc5x5CwhDZHh1IblXLHTpOds
TdVixnQrPj9xtSKKa6TfyCiWj/bdUFts4QRoY+4OrFju0mGVABCOGNNtiumwxWT8
ZWU3dxAAGEcaP1/fVxhwUcOd12iwn42VcM/zVosy53JIH9GQEcKP26sRtXMhnjNV
KElp7QgVutOPHEQyH0EXah8+rKfOSRQtfUg6yRIgz7asCOrAR39DDVvCGcOZJBbH
yrlqU4OrCfARXY+ia8UG8IJ7E44WCXInXpnOaYu094sC+4MGYhNlMF2/vIPfqt6v
rfUIF9vc0jiUbi4eU76VIafd1VMqE+NK/HzKq4NpiZOkFE5Op8XwM0GbIB6ZQSBm
6monybOzKxakL5YzhA85t5HENFZfOemF5qQ3ByPWyB1ZVB0gb/7zpTKR84f2IAA1
vTWsW3KcfTOr/X0lnRFNHNZV1vNk0YAMoCtsCrZj50ZwNAepuXbf4K4JdC5Qlw0r
742lej8Dcu8q8NWnPyumrZpuuVMOpXn4uPQJjxAbeWX0zINlOwEYWeoBrP0M9UQ6
qohiDEsmTLjwdM1/wUdXx0NuhH9g/ePhubrnMM3mOOQjSw4P+lwMgNcjzYj48fn+
X9VDjMO8JMtXmDkXS22OBgED+Rb+cVuOjrcv3H/DK6EqHO37llHWsLaZqN4E5r0Y
ixw4FeBg3KXOTbsZhZCtlxG2IffF7ISGcgy5L9gxSCu75ein30X/FPqkVFsFCt7H
bwcXVgSczNsS1srDLgY0M/TaqlHpwACD18DXUFJOdDBUj75Hgwh1TemZ/5TGNw3o
tlCcaTgJY3o7N55qSaF7SyOss4zqQGTTmRzZPOr+BMOtgNwANWza4zDjWTKo7Ovn
OXfxBZWWax2SQd472hBw8y7Z5ne0scKQt9sMJ1WveMVNLMkWLTX2tzpHcJlZ54sE
LbXT2Q0zq/zI9Id0Ka17wJN0ngtkSut0S7E757tWMGeLp47tG2ZB4r8NdGhVFIvr
f/GYtEanS5cmy76/7gOUKloz3/KTwJNcMUmBIy4wK7pbM8v8SqsXgJEmc4v3XuPA
dY9tcy1MwPnSGQLH84znVKJh8SIXTMM3B+flVfN8TkjwJYTReW3ypT4cfJNIs/ci
yIMQhE4ih5cBiPxE4pCDy/M8agaNjgsfR67lS3LEg5ai5Ut6dXJ7LPTH8oCu1/3c
3DPOr6EvGHPnBWpHaPFlbfZcx5c7oMswcDt4QQZDv4n07XUMfT2oBisT2ZtmjlqT
hnak5/0x+meMz6b8/YDke95mQ3KoSEYeVop1iFVVmyR9o6ywn01xNgba0/gbkKMa
LFEZrXzWQ6jlYYEpma54k6ftXtzA5iwun1B8QQlVfM9SQ2vJUhwRhCYRFb6uh9Gj
9YUYgVPU7qGmv50UIGgtILCQKD02HvhzGuLnZi3S2s0nqcx8ShFXhw1EbgWnSLny
vGMytETingCi7NrstbwEPgOD/Y4sh7PDzFeOI4jkdVUAmGUywn46QsOL9cX+/4CO
8wo39MWwNXXnMjW4rw9y/q4tfcWjNxgasRDpkUz4A4wYf7Eh6s9qOjN48zWc9rRi
m+KvZh71nXxXkXhYQymzr6tNpUY+EZ+bPIlDkJOAUEYynnpwWkSvLeoU3dE5bpdN
IhRySerQtwQxtMHFvQ6bisgHX5mblQMRUo4ZI+0v91prgbBqKp9uIV2CxzcYwX6V
g+dE8Zhc4aOjnU0SvAJpmwW3WyYx2sTvj3EHNd7fZpsW0N8Pbmm+Er1F5XCyi0wS
3NaCeYVPCLnd5pULSNL+9PSZa6cvNN9RyxEQ1d+UgdU6UH299CZdoo7VezLJWAQr
TPeal830OJAx8cKpAYM6kpsXvGp6UrTMzGEc0w3mWEf/9ZgC/nau/nllflJu8Mo7
m3ZVCaaOAt/DNqig5M/INxGXiVC6q8D3+/s1wEkeS1N1AnZKY6100x/phDoo13YM
zJCCS5eo8PFTQ5/zz/KJsGLYG164/uYC6q3hN5NIFVFKQXcalYJK3162Kd8Si8NX
XXhp3vr6XKJXewWmI8J3plI3HaDDTlirnWu0Abw5fv1wb86E5X9UaRA0xJsWdRli
MBCPgGkFSvrMsnt6lBhqg3LRtCy/K4r9/GKg4GEDF7e/nAws+pV+HHWlRpjzGQZI
7PLXg2GKBJU0VsO9b5K2SFbJFWTSV5a2pv5dmN659NHLJFv2eBChnL2eUGXqWzNm
fuN2fzl88Fej+rGCHQFsaQ5KQLNBF+1Nysc5PvjUR+448rSL00f9aAHV8ion1/sC
2BwaPCDqsUJsuiFMH6bZTHSclXqq+Tw6RbfHau+J7MapKsPynXXZZQTODILDeVXs
gKhm57CjglZc1+hydjqoDwP72mMSbNrI/1bOZQw2CQ6WDt8GKYf7G7k8v1e7SUOl
6L9Xahjnc3SbaASckPo9Ih/IN+hRxCniH5WRyLkRBpXubqX2rkisQG5zMOFHm9Fs
ujfcoEfGMqx8WCzN2vNpDFR0kI0ii0YHjRqbZ6t/pCw780r017mGIIN0jUYfVlOO
+Gks56nlZLAbF880JcJxadKfRiUR4qu068qkIGFi8VrL0R8/gs/2zQtTyLidzpdf
9KO3+0gsPyQMWTyvUI5UaapkoirShVJ/POB+o5vxB/3It5FlK+0Np4EKv14I4XGy
gL8c/cgteXY3RFBXp9JQ3kY7bFe+TipfpFuxZkC9gVtbO5oLuN8dgKvNaLGhrNEN
lzANzCyXIXvxDa5CfDd94qgRb5jmPof345F4wHCXMDr0764gISmmbAedcHtznXN6
NlMU3q2/WtfAyF5hIpnkqta4D5Py7brLPdWHXFl9nAG5qljEy9DQQjDDlYE8ZkFp
lsdNZCafUv1krx8IiL/RJTTLTMXF7KhW8tGOL5e1c5wmd2IQtwjKPrph1RH32iUG
LgVSeYEpGUMz5pFEl6Z2uoi5dSv8+DoMErTlrtdhEAjBch6tKMgaIXboG6jE3kSO
cqfHoJ5matYS2yU1A+ozzWTpKx5H8Qhjo3pwfSSZq3Ogs5Y+2vuMvhegZghjgkKi
01FlZkTNPEHF02A5PsUYbMXaYKDsONBWADDh4pQueCgTRNXn32Rzn53HcgCSW+eT
2FRJQ6RkowAbwJjL9m6QMeMWQBlmJsq+zL8vmwScfJRdxoTuJyvSnsE7IOLBnRSa
/lCXBHT6pmhfSGGBerxQVyOVUCbO4OVX+MkTQ5ePG4lrOu/vWRXq0XM9uZGED+bN
ePD5yQeVQevcbgpcKyL4KRUwAJl69GCklplCpyAOnFDHwYQD5CtN7vnpap9T9SMy
CGwE5ADTYGuvK2vA6NaoTyedDe8FemXpwV9RMOtc+uqxL1jzpV8h/7b+fWF0SVoh
RFcZT/2oPRFm2lZZEEgTII1xIaWkfNyQtBUPiQW96dxaB/hA4H+thrS7FVMRNSiP
JDb58zIOsRwXXsyAycV7d2Lx/XqmQWnVnBZKDc0wWSr3ix77X8FePVkdOTf4b3GE
hdrgL4vNvGDn5k+yV+lrkiiI/7Nn1wj5yfNgMj9VirEpOYQjSXkTEk08w3J/SG3j
h3cZvxuckOcoWrb0aurr18An6+4PQdXPXuLUGydT9W3obCxhPpADxnsb05lPcrzV
WZ4U4ksSp4QhlrSg+tC8SRypqaRsj95N+/k68WWZPoNQTSdSTg52zClIXb7E+cL3
U2qU8vkayjiI5JjUK/qakMrkd/GzIp70OBXuv5pShA4ulMWwnsB2NPFHsbxLb08u
J7sek56X6uORbp/5oAqzO2I5v0JQIBqPcYzcOBzWpmX2FQYjsr3/sz5IEPy+zZ4n
UE2Y05VITMIVcuL5S6ZHcA7a0BD9NbCr0mXm72mLj7sS6vOkakvdgSRs7jhc61bB
pu1WjHwVpbt8OLxlO7cNRof/EWw1p7D5m9aTE6cQiInOBNcxe3Dn3pOWlA7l+745
TiqIh1kUuHDGcOhdqFPDIxSSGGHqv7eTBLu+XHJftogSSHoq0O0rZ0/gigVxQMXG
klFGXYflP+OZ3tkVjlF5ZOUvG2Zc08uZHPP5JrYpjGkPYNRXb2GhC0jS/khSGNiF
1AEl7Zwn3E9MHLkDST34SJr39l/9RBBSXz0x0QiE6KSdoygiypNV/Dzf9bgaqP5V
a/wkutgTzYhn7G1KPFl8mUG+owIOjQm9ETkKxCf4Pc2z/2sSsLijtTnYbmgJpUSE
3435DsTudnSg1GOF+H5DhWEJHGsfs2hlRi2LrlbYE7GE7PYrJ5EKHyi3SgTGAdEM
7VOiTPlH1e1wp+eiPXtQimkLJ41o7ou/be4tXyPZQ3rd9+KZAqrZt98llcCYg9+A
kPO3vgdf/pkHz4EQixGmJ4pCL1o5Mu752J4W/A9RXb68cm2kC26OFXRKXAJj+k+W
4yX1R3zdEZXLtVOQ2QvcWSpc4yAMgwOiNk2XjesyQL+uL91eB9umIpHMUVP22+NW
x5yE9luQgOdjOzvHzIgrc4mMmi8NcGC0klB1V32r9ApAcg/Eya4QjJGV+ubh4qD9
ELtlASnYL7NHfp5fsI6UXF52UeXYe9oqpWmht59hyjKYyYLDLUwIoTh4y2dkll7w
wDo7T0bCKgHbejEgy6rq7zMbo6d6ZORqNX8C8dE6gSxuRbFQ9XjaYWcKZ40gDDd7
Dc6J7/aMueQJ2PQB61Pj1Han1izW6wGc2C3YNAZKcYXbPvpeGlmR5UduOGXiujH6
FiWvNElQhE3MWpdFcwMn6EyxuF9AWTJvUACPnQawkoCv6TKL/80rfdBMw5lVLxyU
jJ/4uu/Ge7Adt05Ino1BucCK5BF/Bun1DxjUkTzPJTRX34SFEM+LOVQuIJBxExkO
0a3FsKHCAzZ516eDVWXW3ucuDIUK7ch1vqMrXc+QAPBd1Pw1oB2E6rcu+d4jYojH
rdX1TNJxkEYFMae7Loo+Qs6hxb+Ug1PaRtwc3+2LahsleqOp8a8dmKzzB1roQAeK
Nylo7bKo54cR91/1MmZeF+EkgQDetgewHGy1c6//pVOJPNe1qIhg+KANnRlwDH4t
FhZX+7xgz4JIk+7qE0/zi4zLJXwYXscjOgn0GuZZOVF54hJeTYqIHy4B2X+KbDD/
8ZJmH6cn3OlBcu4hC8pgS90RRYTF3cmWQu0WIyC9sDrZxjszaW361sGXMPCccSwD
bFLjD8f5s1MAKC1LH3jbd0KuAhfJ6NojZ7K978soK27aaQgMziY3+z6K4nvYcHhx
IKIP0Y3Z6uGr8+dI88CPSYDwJUJ2z4SLtMQpjS4fD+3NbVzx25JMVIF/zmgKrHMW
HQvrZ/AGEnROISUGGOFNka4JgHZenhNrrj4LE2wKPG7GNu5G8caqvwBBITJ77UPG
ADLDS22dTDvWhEFqzPHXeet+GbWf5P5q/MsBa/ZMLQead+45LB0mB+4mVIukySao
V4q2Gl+vZqNZywz9qtNJjG/yv2Y90kzDX6vsSg0osYFvl3px5oVBwSAAmEigVS+i
HXF2n7ms0NNEwNM/BycW49Pt4BQrNka7ryrsb4F4gOBnN5X8xSBccTED5+3WyYMK
PT/pWMp3G4MajFa7/n7ICQORtQWBPj5lIm4pfQ11CCqkEgI9SsYaOFwQCmJNTx0P
WNVUc9SgFvtudiE3qvkb3CTf/+89ruifj0KbyClox88rIP9qsjVJ3Yc3T/J0GafN
0WW+pBak4H7Dxcz6Mbbw6IrfRPYFzIJMep+YDytBcYsc6GuEp9u+7/XoX91kq5pG
z1ElKSXPX6I9ZUznyiw0ghGp+O+NOxg8l5NlBCaPCXEVQC28TLw9TKo7qkTL+fbx
52SnyVwjZ8V3Z9ttlBZyysghgdu4DuDKwkcPLtwq/8iVS/IsaOXrm5hn+2bpNTx7
58bBfc8xRf0JvmC0+qvU9Rmu99XpDn/PHcAoXIn2L7CEausqGygzPoBrrMLLHPU+
afNyAaB0KALSHxGgNdAjan+ilE7ZtZNmxRaV8TS67Z8MGQCnp49L3zyESiFQlw3T
qKUlQ0tX0xS6OqbLfEN9sNq/CWRc0+exRkSkYz4RP3RF05xN+4DvaczvXAlT1sAh
bO3hPKad6BUAGhHESrjHxOoL01qhi44Ug+G+5MwLAws5wHMkDBZ4bDzy10+e1+/n
wumVEt1iIxzdKyaU/7bh4gyrcPCsnWrff/d0GdfIXZtGPolM402QmQyfG2kCbtPp
/yJ/Ffs4gtSo2HKncOp0GMzshArPhHZb6nr7yhoDnLjYGnfr3N99Yp9Na1wN6FqD
Ve1GO6IobqkwrquWBf4bMioz/llW+o1thBF1hm71/aQwAS/FkaTi50gn9VaRuS/Z
+dyRO3mXGywG/e8/Rv2pYkHh9m0InamjDTZZshTyLqVheU2+vZ6RWKw3zxPoi+bJ
2//FIG/l3+ir68lNXuzqLLaGkeQE/03JTyiNijiDP8pPh58a5NfNICWAWsnp5qWc
f4zKj3+E/ur4LodYxnkJjut1WToJwRzGZid4f0FzEhu/OcjWTc4l0RbacoNq3eLw
t//fQctntdjLNMWmtWde3PP0rHM2sNqY7S2EagwnZ0XfzCbBKkLqWtzes7pfuWkj
6npxGhQzdo/BYAQBrE6qqrSjQvkhz+s8VWuaWLFSQagQp1dRwIOsufrS9VqYvgMB
Zgt2zpR9MHWEG7W2joy7In4xKSK4l2ZxyB9Y+LwzdZO4A0ptua4+qFhjRzQ6Uuh5
v8nd3rwXSTaVUBaAVnD4v2BWvDMaXx9LY6TjkdP+TsfDEHYB/kw7b5pT9q1gozAu
Ox2O4DjeeSJhKMsNah7bKAliWagmf6GOuR5NEneY9LbeDm5O0Ks/h65UO9XsM7m1
VrOQz7M1sYmPnVokc+dMv03RHtIFpMOaNmJ216BWspOKlsDxAmeHMX21hQ1Y5bLw
XUur7grSlPw1cAPKk5dajqoV82tS7sp55k1YMr0UR/lhTdCTlkEH+97saV3bWKXg
jb0FmVbFkPnixsXLAUSXGT6/lcMWeXulnJ3wYy9PYBxNR+4twe1QQZPr8sonKmt5
oQg3Z2S9fn2WfN8lFY05sTk9OlW+Wl0dipQPh9rnhD4TNpbVaRjvSvaTjTCT+mV1
nr4miu/LOYNg63kwzpt5s2NruReZe7ZW+6KK3iMteQEzvL7se34p1PpFMSTXT2cY
2h+cEOu82Mpzb/8cmMpFGrkSTUlzEWNbks5o8Fh56X3/IQMTgav/AVOHel03rz+i
Zdncv43U86gR2J0VuPNItGhEXyF0BGNd3V5n2KHgWB+ZRXO5Gn0R8GiIggGLgwpZ
WUogNu1ABtIYGQaGD3ZEXn74AKZuW0AsLBTSzyEt8n+TSulBfC2z/ml7dUgyIsJX
cgGGzJ3M7c2ddEgadtt75Bccm30a44DYkgInwqxd9WRQ7DzDavw1ScAIklmxq81b
h61He7DxTodZoUoP/IGN1bnmOuOw/lgT/IsXLgwEwEXHHiasewMQW8xNzVpd3lU+
mgfOCAzCchFcOE+T+yFpP3I1urFaVqD3ZZ9cE2S24vxqjsWpTcljr8UxnDCEoVab
BiQ+0z25o1o1HOnTR+ikmKbuWw12DrPj49By1XurtXns5tImBrqot0Ebb9fmdP7I
TK1X8iqQltm1izBC+C4HxCTZ8FKHFeg4ZgbA+cEAAMuko0MqaWZloMGVWNSIOWzc
hpE6GnVLw7LQi9aZzuzruOc11oTipc4cUgtzcV27eIn66TWpDrKzLpAq8LAwvp9b
XBUHJ1ine6+X1H+oSwkg0gIZd6Qu3qDvORtR1yYStGVYD/UakUyA8smAnXoeNOif
xH9bPgzLYAUokB6gHB7k4dKuoFMYOgB174EaAa7E1+q8jz/2QQ+OiViBKs2Lm6wY
ffAI17lehuROJHdylXxfvXjByKy7bDxm2K77z7vz3bA2WDLe9DBWKFnwP7QcLoaF
+kcM8g6bgvyuwIBOLheRwE/mcEvVquq4zVDql/htiOhVhWncVBe/AIiNk2aDW1Nx
mhIb7Ff5ISTAlZgigl3w+6P6h/gSx883UD7S4g2zhforG2xvT9DgPPTv8czKRcLu
Q/KXnqsalB/OpxP6mhEVqwy27/Sw38OKo8dPtfp82oqi8Bib0qJEZPhwULamJBIJ
8puiImFuc/FmpdtC8kpec4xV+NMs4BuKzRdFEPL2rcI=
`pragma protect end_protected
