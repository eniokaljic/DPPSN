// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PzJazo6xVoB8xptndiBViCF1W8WXCu7CNkkKdLWwfS4NLgQinIsjP1Nv+PLsXWGz
yLFWCGEKSWWKnN+Twac01Pu8l5tXZZfHmvbCUlf1dX8jmBCH+5pGshabMikPVjIB
cXFq7sfJ3jmRWx1QWuxYA+CHMToXRBld+V1fhNT1LFw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17968)
aCNe1ayoNyJY2UG85hapZgPZmOHfSt8ytFHST7Vp+yCxtXjg6u4pPLzaDbPu2OQf
hZWvrg/vUQ5reGZRH428Af0DRWZg1jvFQNWGBvRLzk9WGsyaa4P0UmkU+N12a7Un
nTUBHB/BmS5zDgO6+neh2WegJaeA/MgdxCu4WpyAPtEHHxutwHrL98Cbda385er6
ZyxKqzZ4Nvj5l07Z8jdGMmOV/sYHMFNRao8CPwbyesNCoIT5m+gbe4xxTEYzVbJ1
LcA7vuMBB69pF/NOnH46DoOySOe8xBLmmul5TGmaKZRA1O7dqK7K3UGXVsDb+zUn
egvBvTPJHjxpZ+rYPO4TNV0B/Yo65HscrSamsRX4w5CiQdAJmGYPp+6HNbalfhjd
2QRifQ8yDOXYyya04faI6tDXyWQi5GY8zZHLjvJagNPeZbRK97Xuj41kG78269Xk
W0QFCvtGevcDGehc0hy8Wa30wkvOixQQKPZfIP7g+h5F51USzo6XwQU3yVdqlxgg
amw4ECdJwIu3TDjYtMSqiiqp6Z08BavCxxBCjmJmgY/EFz23dPcoJWfh0Cqptna/
eWmKNlE8tv4fJ19gpNI+ybADGLTIyxgh5umnJTw/ClyspTGDVLDNNrSakzFZqk8F
Z+rlMPx0pwyMWxUjmZLUxtkEkg9yQ+geJi9Uf/vSWY/HEJmNXSiJKk7z+9eC7Iwh
jEF1z6AaZCRWHzH1xCKqDcLygEL18sCM+APZCHPYs6J2JpinpqM8IVfN9BwmDdpk
RAtIh1la7cw6FrnE3WATDUnbKVqquEC9Xj3n2LxyJtKbRAUxe1JYwldqyqykg3lU
7HXTET+S8ZuER7yDGsT/mCGv0AK4y8I9w9pFmaygbeyYew8OL30/HEpn+JO2pXPH
FYmKfAacLGLOohFAeMsy/btp4UtSH9ijh15ow5VoKwNSrugo090gU0HwPY6+SYVi
CDNcQq9+sc3Y75bf1m8DQnkfQcH6GmXM1j5ie5KFVOydxlH5Mf9VB8tuL4ftZQ+9
nO16CPYvnqy+SqwRwDKIv/g7DeTQcSXifEbJ0imFpp7htWiwKf77D7+hapXTxQOd
Z/hrXNLMv3BPDBUeD70nsCd7pqNX4tHpk5AOJqbGpLWGtwOTzJ5PN4Yt0uWKL5VC
7N77Q5+EL6ymyGEjZDfV+oIoJ2TFCxlGRl1tGDb3ZNXkxzZofP64xKqmfSNFo5ZW
cfDWtY0/5S4jUb20ROti0AqyQxl+6lXp0YubjHcnhVJWkhUriepFKEPvopVeFBYR
jXbvFMY+BqOk8lEShmGb5oXGr2NydmGqFRw7jhZKMDQn4cdDBU2jZE0LjLcy3fVJ
chG5UXiC3vA95koUrfuhsND9UWv4VxK+xO0F5r/Qd5VJ+LdwjmU1bJOtU/0B/Sg0
ShqOFLdOeYgon30ZU5p7kEhMfKHf3IJCZyrJGBco73lqMgSVJdAPk4EDHvV4VjkP
vFe/6WEJ5cngiptBUC483Hu2X0hFz3U1a7h72j3Dq14OjkhTKFL0izpmhqv1jTC8
M9Kh8dV4plad85BWsY8qulNU+IulfIatEuylLsHqRBApA5OXXHFwBhO8TL8ZC/iw
DBV+8PI4icJ9H5al0KcsboVnu7+DKlzuANLH+vUzL5zbJKtoC8jES4fZTVHJlrG6
4kc3mXEXPRBNrXPHsukIXdqJzxe0gR/gjzZj/CdtZMGb9FENEqovYzeuq32ZsVbe
bGUeQmgN7ZFuNFqnV5jla2dNbk/lurFZi4QDWl5yPrzqiEDpqc7nO8GZPo9JdftD
DbDRtPB3Xw4EBHtS75I5ivJzQkBlWE5B3UwMhWRUi1Kr4weBJ8f6H686xBWdCvGj
GUTotCEPo2rYnJjNBGG8TDo53VB6jPZWnXOiyTWYcB9h+Vxr7SfYZuA2zLjZfoO0
EuJehOFU16igYgUWg5iyA5Axcy7QUCrFR71tQHv12y5wF34i5sfboYPNdnl+Wh9f
sYhQscS/Lg2hLxm+WWG/QSUxdC2HQA6kC0krfj9uIcGwRIdYgraAI+PNhyFa12hu
ERRB8n/erxWQsHyWDnsMRL2xZgM7uwX+9el/n0ik02GiylZpqMdJcim/lpKgRDzR
ws/eiNHNl7xTRM3f/+TZpO28/1BqoWK+30oGoPoEgZWIxV6gDPbKpHhuytOnHuYJ
5aSogYtp0tae0ztPvBYoGm7H0V0xpY2nX4w13J4utbMvK1wWGP7rc+Ea9ngssttb
2kFidh+N0ELnbYsrk/MLZAyl5Z6YFoevUb1uJdh+sEDGbEEpHSnBEK6tjZuzCDKi
m2xzJYE0CT21ORKON7pWEZ4n65LcvSr4gsYPoKFh0o6dZ0lRCK1Mpbf+EGikMtLm
1uALchE/Kp55EvFP9DHdmjQ0/HJo2TMx3gxOo1kqC2uDzxk6te7GQWO7IqvStjnk
5rkcjwJzLyfKZdk1OOY3sPO5MIxfk2qTzQimTXedI6hN9pECqjxin99N1Gn5f0xP
kPiqtYl9YVPZuWmybfaWTisu5ubpRjY0XdKCeriDh3dd9YhgpAvCpoWaopWkeRDA
6IQxPxEyNjVxymnhLB2wSn5vcsUTqYC4fdmslzNIwe4ey2YT4v3ONt+J8Z7ChdtS
aybI4HbSfDLzxOOhwBFwAaaGBdFdZ5rTSs7rlGlRZXIbiToy++q8185ZccCSelzb
XiZ9Clwf/P4qdvnFQ9qFo3Yze4q6051WjCyHaFIV00qyR10IBn6oJmBGARhFEcr0
WixlbionkvHDqhQ8ocaVax22Flt59WwND26R6G+DceY+EnfUpWPK/9VyFPd/oNt9
kOvBWCJzX+34DEiCuOITF/t8rlj0pF2/VRrBbCVdBGO9FEk+7VnfRlJvy3uC+2W+
gNos3RdH8+gZJaQZ4HXzi+MpMoFykIBdR3Ov3u4mfz9zsW7U4waNtkTlrpIfEO5G
L6GR2FITXajftlz1+j8fIDQgbxOBVeqTPujDDjBXyaGPxuaAADrb15b/utPQ0pqW
LZTqxNajr838D5g9KlJq5rA5B5HZEvZQsziL2Zzb+ehD4j2ZFGbGnyADGqZE4SPQ
i/l908/BeIumJf+PBJYbWB52BlqWG5j2BRCbUrmxT84UI1kShz/ghhbh6FCvr0d5
5uUZ9jw29jQguVJjOM4WLRwcS6lb5z3eDl8QF4v37wTE+cA+6BLISyJHKfa/Ipvj
LqhNt+UX9WhUifhqLHbbk/TroOAoXe5MlmhMvIBCKARmztdVy2hr1UJWPtIBJZmi
U1roAaVLoT0Zy07y5FMFuq3jBah5lMSMnd15TWP3j9jzV25MgQgVRfTlDCA8PyET
vm0tCRVm/I38qmrOKSy8Puj72MpfBGINZQQiTeICIUrvd88DxO6O6UEgEFlAQAxZ
WKKQYSBMbWrNwV+A+qXFxEewfdO6td43b6BvqbPV6kQdhhSp1DmzRAfABR1rEaTA
35C9i34Va/USfevbbBjlbyeQmD+fyP2x3dqrvFXLOl0Qq35CTx2o37JsqA2cbDNe
JDSDCCsnICRgMPs/ZqsllGVEVhutnNdaXycju5pKmXkhWPfJ/nRDkr951tT+OZhg
/ssX4So5Rjyy8lB+G3ksV1y6xz3ePUfKh95MdLjkTDq+pDP1/RCo5ljwmmYIuFvp
VomyfbsUgKS6m8FsO74RSAH2fn2nC91hwI7dTFuVYtEWHmDX3yOFMUqtyKx2y1/W
F4qzZ+96gjy1gcKrjbdPav3ZTbYMjV4aNtfMQ0n+GwT3mdIkqOV0vBPt5COSRSUa
3rpznMUX2piEh+I7cut5GkzLpsPAlEMlHRY5YP6yV+aqeGYhTQk1nuz/f1oWWcmf
NA4Fm4rIk3+jqdiJ7ZGzIL/1i6UGgwvj01AMnZoqKFzr0uyZ5cRLOIgokJ5EKvqq
tNWlTYsN27pIquDosCuHy+n36/mE/lE4jS2f+3UCy8xTNkcqFCPnsXRtpTHg7nLc
7g5FG+gyS1YsUlqFDrYE5EkomO3DDXmq8YcdF67lIERmXg7wROxWn8/9ygcZU310
WbY725rNZNKqEoEcps1GsqFgkhc+oCQJP7oQ9+AOwMZvc7NraMMcluKMWil1bTgl
G/cQ4t0aVvmSHs+KB6Lqrdq9SuFOJsGX1zBJYKYDsqn8p4p87KHby73xQggEd/aW
9UW92JWsV36Cpwo7wu3ST/M9M10cIAZ4msyprLGUgOU5KMoUukn+NSEODZTZGocw
irNxf/3o4J8gPgCt/5Sq4JMXfnJpNUlHDYLX/t2fd1jcmOkXfEjC+rYE4qyVrPpm
qhBSCP/fL9RK0+JpwF+AILoLXjDE6fnzs6bpc+ZtsCVKwQCwYQ7Zzz1I4rzYdYR6
EnXWsBLVnD85kPszS3y6i1pARFJWPCHyfcKlurgsgkzsq7uHYD92vL0ciQKdHKU8
xsyLXJAR4bfVJPlzXQ9OJnqHUeIcMiITRx8ik8ldRwQH92TCnVG01TiwIfN28cSL
78HH+VQFASasFnTTdrFkEq6tTrc/cYmBLu/L90++3ggxnvXnaKEP6diHJLmSpB6l
bbtvWpTcJ0e0rtSYHEOpCioIF4p9vxl/ExKi5wsom9NVGlNrGYYh9KXE/fA+oGnM
WZu9UQf7GDDpnin1y+jZWNTlnoAiV7JKM//+wtVB6tRdSUcw7KYp9HlmlDKFDIcN
zM6fWUQrCv1xiLQ47eiqSXqMQpo37Xq3ylvWogn1SGdIHh6xrf7CT0fVvbgfa83b
pO2gBkNn0eg4tugza4Q7XnPFG/XkGEJjtnu8bUO/iUETG8DWYYqJ0y9CuU673889
9e8XysDbFPmkVABi6knIn6D0B/fJP4OZcMD2PIwy3MUs1Kx17JWo6Zk2LedH2Pe1
SkL8xa2DiMdswEoNcu10fc5Mav1rvQSVvV4dKSbohLalNISVrMzhe9HjYcHduu/t
Ll6NNMDGqpAgwUnoEp8eXYBfqBjKOY7nlms3xM7RQ0KY8OpbNXsXC3zL+41lKck5
sRF/rY6eoOPL5XCnFg+5UEvm0q4TVk266Wv6Av/RDBHdB61dN5OFam6CZEhv+kgE
FegoY6uy76HOVWTgu/ReOQcf5FZoSLX4bweWZ4HEuz81Lb1sNFvOjtYd0YIiejDn
+Gk/3j4AYW4cHNflYUUstm0h2TNEjTjbJc9FC5O7ydY2zUKzLOdw8wywVx//ztxR
Grgckrn45baiOiFeS7hggzA47pz8ad9HfRkxGXAqER9bSLxy9wQ/+XWwD/IOZXSB
ZfViGtH+XJBDgO1mnB6W3f/ASeC7BMJCn0StWCh+8xu1XzED7Necfeg7p9NZiEXS
K6Jh23pM6LrmtC67RBbcOlV7Gjxw5frntIxVs3kA8gr3lZKeCsfaE1GNOhtJJd6R
WK05hckGCYT48wKcIUNrzWdvfcekNczEMjTexcovP5muMVlMBg0kzYxY9QYW6Axn
m2PmvC1yFdBOacKftlvBU01TEHpim1QRPODyF7RGIQvDI5ZrPMxhNHIKv7AC08FA
Iv3Fk/wutdD8lpdRLEpa56bWs7u3Rcg2qBDALigmFFPjwzGpsQsSJV+IzS+jVHBx
Rgehr7n/Y9G7sRmAmVPkFEHCWKioM4n/84AF/wRPhqdj1uQpDAIJkQyRnROkRhVw
7w6rmB330q+N0498U1FAUzJsQd5HWgtCOxnG19RvFNrbnrARsrvDbmtiiPmj03wJ
oP4g5yCzWNifmz45RRrbeqIprsn3mk536a/7cMttH+qaqx6oY4QXPuWjEjFP89Pd
P4gi6bBGaCQ3036vqRvZNMWkPMmMPjtDb8jXDTbR4QWXC3fZ+NcWUGlsnfQLL7Yk
TX4cL5RfY9hQgXFsf3C4DCZyu1vmBvSBpU568nXpGGvGusc2Kloq7F8H0J0WdcQP
1FTq9hgt+f7dLxRc4xW98SaclxnIX8Jg0U+ukYV9MVRp/pQPhe0rN7iddEGXGyq/
3jui4plKKQnN4indlLn1FchzLk17RJpQAG8P3gy6Z/DvUM+XBw02EsLOq5GwDWkG
+dUCBGTxWLt2oqdD45tIQ08pY0z8nAi87JPUf/9A9F/lclXcGTjplDi/B7HwEfy0
zoQPmkg8xBgyUhq3dz6dDm6sngBUsFOBd53HdGnEPnS0ymQVWpI3v6t6Pko4E7pS
4ukmNl+Oq/gKEDSI+aurMha7J2igRw2xo2yE7SOPoLJexRSS6ogXrPP5hxlLSDLM
epbo7zlvRLhUHdsiMVZJ4W0FFkv6v4CusQHouAUNwr+4ITV8ouKTReMFeNRzmkYL
+JEGMI08QA1gTHbCoEySxs3Y3QkD6dPHdtixaoedTjyNr511UtQG8qWUq5yAV+Ox
1c1tczVZ3HzZ1l3GQhOay/C2R53NEVf5b4YVj7g/1dRJL9eC6HpOEDdnamc82g8Y
0F1NsaOx19AeYQ7n2GtAdq/HafOYDMCwoldVgVzhDNUWuTIgYDaus4pbx0XtipUq
L6pcQjWr3/kQRCK69deKj8NT3Bg6wsfSlh+ywmoDVwQortC3eJ2cgYGBzmEZYfv6
93eISgACB35vH87FeVwGuGEsNjyBZJM1/azv7+FVSWfqse/RCYYgnqmUWVLFm1wO
o2lk/mjHzdINfKSJ97oNqFUlFrNWzmknKFZvpeZbY63c8B9HPTzpceVryxROEf2N
yaE26FGAoLynEtnpgmD90eK5xOujf3vVwYECtPaxEFwpEiwiM8CSKsOm5ZMKpKEI
gxNwWjlVEqkOLuEGyEOFkyTXyRPMf3LvTEpHF8UUboz87h7aqkMU0NQYTruq0BF5
03K0EScSf/W7fJTfw270Rg9wpDA6e2t9329lq2uMfSqU9qzl4ZPAzl2M6aep3zV6
qM5XYBKPktzK/pbZblgfWhWXeZxOoSmyT8I9/lGl5UlbaX5CJ8OfhjGt6MuL5eYr
xxdJ2tOvcmk5R+/ZSWNLFzHNaTisbUNY2v9r6GmUL2n+4as9pu8g4J2vp6jrvUVY
cjuXk/rqAjUjRryTP2awJrYvldHD3Lu/zSx1W73RGlHBEk1lWF7rR31X2pMjoASz
5yXXG4ct9zH2yo1HddNClYmSYM/0nNHDcVbVwGeCSExd/cdh1EOII+G9virudf2P
ONx6eLuM4jSeQF0hevdYUtZuzBkm3aFcL7qlh00bZANbIzOZ+Y/QB0mosayJhsHc
kSJ6RzAh7++V0vfj3Hfpyg1nq2Z4qUCcKGCoCg9ETBx83wthQJRGyQ41G9u0CXKn
YcFXHbX/TRsQ+PYZbDBMGuGx5YodGSv6/w78AZZBcNaVp/SuWYcfrTbDbxDeShrZ
rlVKnzUBOZyod542gXT2UL3a7pHfoANlDTu5K2Kk7pz0rDUETsBz1myPM7mLzY98
t6jB+feJ+OQYrsfX1oPGsJxmKFKwz4FODtVzrS49cMM8F5eOLTcEoR1Zuj0wOwvH
Ty5clKqFzyzcCSQVQMebCyeKPAqa9tCU6C6NHermuWs5qm/cb72ofcfIGqapDmnh
d+PQn2ue4G9Ki1bsny26/fWnmgjzsfD7LYdfa/LbQ0uj8vm0ri/l7ao2Y4PPwH7u
L4ggrN+ZcpBa4E2ZfFHqxMJzzcyg+tifX1N60J8AkmkblOtd9HsdbiAqMWwRTKUe
ObH9ux/G8LFSdQeb18iYdHKiV5vu5VZuoNTjUeA/ytZYF1IDWu76I2RAl+RyWkXp
rfxLtxKtYv5xgTH9TgmYAPZHmpNORvRrOYSYhUwkTMOP4jTAFZgdHg6euFQuXbHs
Swabfqx7sM5N/pT3YryolOnnRWLvcHlFQBF9fX4OWIQD62bgfCO70mxCw33Giwbm
WQXnYVI4lbCyDpfm7GtMvVHukzH3Iz0dSleLIh1UHQR8xnn+zov1D9nIqX9t+cQ9
CD0FO+z6XOQCXRQo2roDEVbedK0AcsxCXzawQRvnNPZW5774TC3/PgKSriZ8t6xK
FzLnxOGBb1qx4uU9lSfr7pa95WDfW1mi6y8Ug/y3pnIxXdI3g04S7Cz8eLAS0oXT
aMSALhQiGq2D9JdW/DlL0nd5+ZxOH/qDcnoW1bjjcm1D1xjQdzVwACREMl01paCZ
Inp9sA9Gh0L/wzp4gRUW3XHxEOZdUIkG0FNAoiVmF6JBkwzOITQrroF6jOonYktB
HfhQTqlA0sP/Urid0Squbf1VTSY/Tk/HV2KqZaiZftPb4/UeDBITIBt3OXwH1k5H
g/VSHlQcUJFULcfQPwPkiq9ZnYoXxaG9j8MP3q0FztAdcesSxsVP7Q4e8AO/XZDS
qvWCTSSaYf3NMqGGVPVZU0I+Ik9no1C/WI2X/diqARfreOmaoZrQZRGFyIRJxVME
ZGSPxwWsFF2zokhdS0f8Vx4/VeXQeVhv1uNJ8k4FyY26WUF2Z8RULo6dw8zup6+6
kKa/YzrW1Plg3RDBnGK+iiJnSom2xohgvjEhFBnnDptPyx9cSt9A6Vg5tcAvHFOg
5H6S7iHWgOI7F5hhLERCkcO0Odcnj1sisj2xNKSH0q0tNno3DUZWTBpPtR43A9KI
ZrmLqa9330YVi9Q0VPG1A5atc46yWnlDHSEUkVysCGiWzyu3Nns/q2KSTlcJpxnA
DLCfL1bXZRE2WQ5n4esSg8yPF68fH5vfasgFT4a2ZFyduvTxJX/Wf6eVTcenqQ8r
hHGAAbItTkKKtsDxcwXF566yzNnBv4tob0xentaQSWxYIOzR1HgXzSAYekYhJMmQ
sPobPKqw1AjU+YZ3+XEtR6T+SxCrJGtTgnVB/1YnlwDIerezIvWQzSZgf+IyiRF0
97y6MOvYGq0Ba7h7i8Pf2b6DoCQuXLN00n4Uwv6DvL/hkibt6/5dwC7iyeSAAuhO
gyIfJHKux3a0BIK8OCGoM5wW5epbhlq7hyQv/0h3ukt72oK45cvpPTZPk+WUR1Cb
++3w6OitXyRL8mjs+xXqBUVfrANUJhO9EKkCyv4SZ1gHaCNu5HKr6+BvmuIdQNUj
GngmyoXbsEJj1DtvxNNIATEeAdyCq+EVZF4YgUzNZ0sIXQIkloFFBwDQcs5n/71o
SmAUH91O/LmAvGxKzRLQWKdul6iTPCRHRN0DQmRwuvyYQ4U2fb7YhDbSXfCC2vXv
VojS9n4Ps9aG40EgHM2KxPayBmEYSATalLWnOtyAhxrSI49nTL8O/8Prs0o0MGza
RhIyE8mLL8TfFlIKu0J99FxuAK9vSB7sv/FWVb5b8+pN9C5T7eXQ1g8A2YkOkqwX
p65aAxyN9ZkcznyBVQOkVr/lGTsrbDzAqSwyhcuVFoJY2aIi9AUcLlMBt7jIteo6
tq0oYzUMx9Xg5pXGZU2et2vLTvtuaZflYG10n/g9/cQH/D8Q7ueAgcujfz1++NpY
JwxwlLJcMEYatXlgk72VM8Ij8SPv5whHCPZNHP5aL5GvRpG1+mWNvwMESsEFLs27
k3Wuga4JwR+ZLCTYAi++NEEcOscwxyKgV1bosBwl2lIhOxwkV0FZ/tPJ4lx5/4IQ
FN25yVADKPrQsC4lYa9Ojy0IPreRqb1QOch51m1x8Oo2CkE2hAkqvKIdPomv0znB
pEnKXWmmjZm4g4co4kf8anZX1ZgSh0GezTMPFNd0dRKHT5C7/MaRhLSxH6Abxn6C
tKZUGvJx+UsmPtGoZl4S9vKK6G5XpAwDxgIidYrMR+kvM2OPvHiRNZK+supiZT2c
vAvBaBFFByXZWy+Ocit2c5QhCp3AYZZIli+4nPKbwofWrIuU0qukGJ59TCy/OB9D
RBTjiHWd2ypAzdiPGXSYNRfmIGtQhMjQ+eQtuFCAMCHNW8g2b0pmiLowuuUuNAv/
giyZosSLgx9xcIWp0XlmHAfyOVRnIjnU4Tc1xZ0Z7Fx0+Xyq7Cj0KFyom26YU+oU
XUpTowd0uSvXSXB0gGOjLFovxs8OVl9PkKpZc1hYolbdWa8l/6IIMPK14ohhpnHL
382cP+rsKd9MCoRQK4SS2Xz6r2cWe6WvhONzI60hwRzGhAYkjXarMZ6RjJJDxKlv
JjHOhuHH87N6iEVUWzy+rYVxVRAPAj7SWCz/2EVNFkv2HjDTaQdcOjpbr+EQKRCZ
EAkv4ACRiaF52oe1xCjoiAs8kazb495F+vZi9Auyil9N6SBi4ThygAZ7Vn2toA8E
VbZ+0rkmMZ9x87sn4GsOjENbvWmw5uBp0RhYxkhd4mjBUsmkIb+cU6DXtcP8P1Hr
sCwfvte2rsmvWfyU1g51DJ8p09l0HiPzTsgfZvbiHlipd239PlRZQuBpd359kRzY
MuxcHAgjGNabQ13lx9gAFzINJXpmWvXJFLQ59xoXFuJbbNjIemnGLfr+AWk7HJdl
auBvmVjeqE1M28BEDh+eVfgTC9YAhcxqvbgvXQSgDD7RZx9zXcVUtViASSFuhnVu
9RI6Hd4FrmcrpIcm1KbJHztqWs1WhpaHEESZQiw1lTBXpY/ZsWfuPYThrj/h9Wc9
46pQBBT94Qq1uDtHocv7Jxb/qXJfG8j+tYiPNWlsldiMKZzHJcCEpqaJTY6qi19i
JqTMxcPhpgwKT7MOFLXmE62fz3MQ5vYeK2yN8cPqmUUxO92CLWRsQR9BlJSCGDao
M//bFFUatq0i7me27PJCQrF2lStiRiBK9UQoNBWOpL/3r8yuJet0RDKF8a+cAoCM
mO4xy6qUspOHc/4XVlSliO0B5VPR5/jvHtaibJ0qYJrw/zoZOk/DiDxcZyT1bLXp
otysJHf023FBXnz6SZ4twDyOSJpBwjfJ/kTZOETMC3/vzo9sRm6gQehbOvILTaQu
dMOI/tq+ZmguuaBIqMqE/Qv5ExfYYfVlyv5EbhJI4WC7cZC1ltXu/ZYS69eQNvpC
ArsOGSCGhId4hUWDMT4LOdSWJbsgf84Dy/x63o2IA4Ll+0rUeQdKl6oflzw56y/y
Vyu+9TWRq3+8ropD4KTKbEhQdnrn4Go6nGKqSbjE3zEo6Si+jhcPRueGkiO+TRhR
ZMRTBsk7Hw0vYkhl3caU4XLQ9xHkFOWDQwob4fzae5srcASxtWNIxxwSYB4f/kA8
yPoyhV++KzrdWmNDeXV1wFAHQ3kg4hW3Wzc9zQYe/ha5JynGHYPCtzPZC2o+02PT
Bf1PAMWdbm+J5r9L22oDNRC1mXqk/7dNA6LYJhlgq+rrYsjRFhLP/mrmB2nlWVIm
Xg9ZoP6/7Kun7LHwhftTwaw+S7MDK4UFp9bB4447A1VgMxdkECdk40hcMdmbnHJN
IOUtBqhrDCE3RFSfOR26qVe3+G5hXE9nxYDH9XBwU2qlMhmtn+LVOMwVndsr2rij
yOoFKnOlbvyVCzdUeRIsMiBWsVf5n7GZW211lR3Ho47HJp4m/tWBomLtiqkMKzSr
92mU8zQLtSNWJX9tfW+RthLm3qs+eZ9kgoVXlq8thSpNOn8yt3qnzBzKBVIwNQFA
rK0UpQhH2w16Gx8sCZkUjGtQmeGPNHvi5Auo+42tl6kaJRDmKDTJ/sZndoiE4v7e
79R2mW4Cw2nqkQdRcl0/YllslQ4H5cj1f6f2ECzVXueBZRQ7/OxOeDyjr2fTxPAD
2fgXyUxnTZCCt6TOXaxoWLZtDh6VcAWNVkOKDEC6+BSQ+NIwnRc8IvU2rrWlERub
+a8/TSWK+eQeI2wlwxp62Ci5XjoeEt5N/bjSe2L6OaNF3fT9hnyAhC0HhIaNENt4
R+Mgsu2a17zljVkWPLCvuCuW9VDkiY+EYMmfQ5J46qt4EGcokk3Nn/ozIcj+3oMc
aPAn9Ipdf5q+8akxudKRNWH2338lXOWHxKoo9OWq6bgkyloafGbiwCOixrZF+Mnz
QjeCHD2iYvGIYUFR/fSqpV2wcAsyFNTpHSaZ89YMw6TRheBtsP76uWWOjVtJkzr3
jJ/P/VSmshqWaZVTHZnSZ1WJ4GcwOm4tc1ZG5Va8kX3ea68D9Def0xpOejJdIe0f
oH38lG2bDiALExw3er0s3oR51N8x0LL6odvEBUeEGYgpzmdzluijS+Lc2sMmDgy+
xvnPMTIlodtwL/8zlTYeIxq6i0Lw9x3Tsr6+ND7Z5mXGRO/APNd5KHDDOjDO8q/R
L+4MAeb8kmnzXrkVATCp8/N4C9H8MgVW3vdSat/jAS9GT6TTjmJcThSthbyXYxNQ
EziCSEogMwq8SWLXoPzXyL/PzcT0OFy5j6eXxmJTdeiFVFWuKYHeRljo+k9yxuPU
zw5O35ZOtDz/zzngKKfVL4nOixGH+zRwbhRuDhTJ7LnS+0K36e/CRt4ZxRKaHVbq
HM8YRm5nn7NlJp81e4YdH+RMqLXsQhxBgtgI2CgWYXeCYrNHKe5TKGsfx+qMfMeG
TwHhRbxPkHJK5tvpn2fuq888pUfePvMrIM0cfkHUGr7xYRGcUwHZrCuPotcELcxY
FdpJF82Px2OptBbAhHtyTe6iFwK/6XV7N6NHwjNZCLvREgvcGxLpYUPD+TygJ6N2
kgL64BnERL4xuENR1j7NN7bLQIRuacfyoZDLCe/RUTOdXo7VBpjm/l3LJWUXyqK4
Ad+rcJ8nfdQVc0ccQGIAuYJRCXdvx3sB26xZFLRyAvDYe9GrY3YDCSUdk/24bY1n
xz+dLpSVoDmjRECHJ/VajtB7Tq4R92PTUu4KFXbLKxyio3MRL6aHhhgQgHUtkGBU
JZWk7nlUo/wJrIEyOqPTa5gOXS/I/cCFw9F+jI0IkKsVamC0CeuFvMLRyTWn2EzF
VTF/7DsrtjkDyJzjG4NwbjmE8MQiDSHTmw2qfdi9jVk8agGH5oC4qqjX0BcA5HaR
0ld886cguaiWfuZc0mc1oZFuwxn02J73r72uES1R82Dl2sG6/6xWkDab7pCK33iS
5yXk5Oo4/tXVEDJUu1I0nnJ9MPdwMipRPdwsaVckfGvZqPDXy29NxKXsrsTGcIt5
NoiemzWRMPKlnPM2kyZ+Oaz3mxKWkSs2nN8snbA7/lBUuSNsd3Ni01OKDer6Erdo
1PljpdhxLMkAwgiXb+WGZXPsFujF2Otq7ds6K3c1YZHACkJyJWNMbyjLdtYrAvaS
jrjQLnV6yxryfRoC7awv1eCxagsDK1yOWRdoILvANy08JadbT+VA4pd1zjx4t/Ga
IKb+wy51I85OB+cH8osDrDGXpdd0+TPvHHTtvt9sCYeK6F3pJOgB1vWZ7RW0GqFU
sm4adXp47c12qk90+6f6m9mERZVd8om1mPuDBTAs+Lj6w8iDg0sASdCWUy35zeJ4
avEu7c3LjV8h+D8qLaD+uhxMsDgoY+Mg+BtFExjHrUPrZyMR5H4Ni3cKBAflZ5ep
Od48XzVf9a7SXt8uwa1DBOaC8lE3aZWrFLdSK9Yb8wSRnoTmgw1SKgBJMAoWWxIo
9S3y0ET1mKm8vFBlIQcMqDqWOXs2MGktEF0RrSq7C90PNMbvEoK3KpQ538WT/9d8
gH8K1V2NHcKXKZe6dMRv+hDwQJepCkSlbdk/c+jk4nejHGyzjW/k5x83WAytDQuQ
KYv9xxK6WxLhmVlHafQc7T+seWZzWdlLWVscL7LUde0VuK0RcVW5q/DSFivXDysO
qJhNO8OH4qkoSQhwshlqcPbZDIijjSlGlJ20MWp5/xwuXQzWCQptsMj+jlJXI4Xd
QbUm/Kw51q8A+3NJhYiMFMDTYlOWINLhjXaCaDGhq1eKyj8VCM7eGoRUNv5d66oR
KuPFPTv5lJqRJPkd1EllzTRJDK+4g18mq6v/e7kEWJP6KLEaDyA3suYU+Mgkr2nn
VkdZHvvFyshYd+Sx0utNpUYcId8H9ISgIxka6/f1zGaSKfOguppRAN8Bti361CmZ
lNRRwgWbEeW0iHmxN7C4aB9LRhgtmIk+TgA5wJUWWmkcMpSVFfiSpPYzzxYP1/De
/nVEVnarxZdvba9woaQS9hw6SlIJBrh+yxVGPuk3D2qEvSpGkhYQD+ZRwzsP2ZSg
IhVkCusVowkbkwd9sJJ3BMj6yWkA6MuyGjunXNRZGa1bdtiF4BZuNe7VH94iKobV
ruUs8wgQPrCBpe3SM4yHJ+JNstylVQPnztU13okhqi5TSNa9FuKGajcdnrbpB9Dx
uM9q0jxxGszdxzmNCU4cufuopn3qDPR9UbZIbn0haLlNZWGjIdbHn0QLq3toV2wk
+m7hmiruC4LFSgN4XEtjcxP4kOCs3ua3a8HLt/giA0enLApoav3ZAOHvXeQyv+v1
Fam/wl09M9kNC/uvzUsUidiMLmarklLUk7GRjfQ+YtHw78AlbpKsmmo6yVIyoX6h
zS8R7geRWz0CQf2KQ9w/quCiWa2/NHoA5IHpIb5ZhfPjHfpsbkRZ5mCHr5/IEl2i
rZ3ZSC+DeDnnakmFRkcM8+m/5pmukrKfjt/hy/n+ohX6qY2/YJwyFTGzv14xc93I
N13GnDKyRKy80qyyr/FyGTk5kIqVrAG6A3RAETFhafyg3npYfjhyJdx1H80b7ptN
xUcl0VoqxNZRENetyCXzz462HOvZl+FypBcwD4OK4hH2h1zu5EBDgWemKhMoqvXc
9VlDivvAJpX2pX7pvKDsEeQz/syFv+Fk8OyDYaR9LzOfxDZqgX6tJ3NA42Koa67y
bqVH9RnqcqWSn+jm7YUMOMZV2cHEMsdXEYlt7zioQ/DTl6e9og9kJUt3gebEB9e9
jAHMBarjnS3PDpgVwnWNQW+aQ2TZvgHUid6dP8llyHVCtWAhTnGfkozG1tBKGwX/
4p8BTGqkVsvsbUY8KrEZbIxp69tzkWSe44FEFREW8ZGeSUM0BipSg0TlU6nQnVwC
Hy4yhsfjkne4htD8VWpN39QrWaQ8GRs7jCLCo5MzozXxDE/OjWUq4W0U2SEnYW2e
mvdktxnb8nz/aVuDwssnHwXdHeS48Yi5MsY+NZiu3I2ya/98W2e4ebhd/p5xz89q
NCCCXRL73+sXvarZ52Pdq8FsZlRYk7uHciYP5A4fkkvJlXU1Uziu/nc397lKnQ12
WXn45TmEp7Uj+GxYQjJz4LQGvC1+GwRir/DBDAT3YNwlVj8WrAReYaK4apRVhB7a
mO1Y2xqNPiElg6GzudIsa87rOE218FHr38oOARA+jYLtsGUeLJFh3/BzyJctfB08
bVnWYMd+XiYJYqTRb4jhk7cxgOYFgpJUfDwvo7gkJK2EEtR/GmhsnC61oSuiMigq
xCeQ9GdADt540c6v9EACydim5a4/zlbS98B3AZ9rlHMhHJ2B4JMouCxkvEjats0s
XVSnw2/+Lxu6CLJ71fpD5+mKS9EWQMcPBhWdR2Z6mnBI0iCBXzoX81BvpLrENPKR
tYF61V0KZYWSRdemKLu4bNqdDnfvPoHrkv/fXs0oajbe6tflrP1Oy3wDPTNCxasT
3LWw8NAbBvbUXzBGGwxPidLycNPLsM9TJJm87/TFyvz5kSHQd/626WgUebo643NT
bmxK6kLUlugv53FfOHLDNRMyOj2bZoc3n/KmgTuLD5yeioxPXfCDYvWuyBoweSZO
bPShfLbYPGCg1X8Q7khQlP1kFCYq8b9x97lloUkpxFuuC5zUcZkvGBTmlPLy6ghF
nRqgq99CxhhEutLOX6SB8qJ6mnqI6HGgQgND58VDQMWhUIXXyM3Jvag1XV+YNlcv
RnnksYSGqDg3CopPIt0FZYWA80AuhHLZGktaf86gnaNQN5YmthyRGc64jw4hzFP0
y+v7YimdWffiHxeRtOHWrZLFe9sJaAxBIGC4PRHyh44S7ZaITAIReFO17yjmR7Ee
wPlHxkHqDVi8BnYcjEYARuBbSF6USDvM9Zi1EzBCy17lYdCT6Dt7WuILgKLi7JCw
ricz1RLdEdhp6dyXWA5jXCfG5jaCWQoWMDj3N8abarvdNro9PPMP06MPje21nI51
ShP6LH405xAkWDRBZoo1m3B25BFiFZFHi6cBI/IskmPwEe6ymT188nVFfEBwv4sy
/gkz9RjnmN+AKg/tq8nC8Cs3mJ8qIs1v3++zUMt6j1iiVVSUy56KrJeL/r+/FAl0
unuEUAEEBwTW0mQqlI7FSgbjMvMx7+gmZiQ064UUUDCgn2BZv0X+gwOnA4IQWbG1
dnwW6DSRH8CFVlyhBW7OBv7t/voJJ/kcdyVvmE6Ch3ZDeHWTnSx4+3zMdSxhO2Nx
TxCFpIoaZFX60DGjNRC3S/roWODElHWrxqxtUZJPth2pREwFX07768u+g+XQQK96
9/2j1Nc5zA7M+k2E8I8kshCjFINOg7BdfxeidzGF19r6mDtbBijww1WzWaXoyCnY
yO/ZB0h+JGjM5+icT8itHBC9PSOr8ZSuVh7ojyMynaGsNumqm5OOqO0eg0R1iSGQ
nXcjCS4HyAZe1K4f184jzJ/IsuNTjLpT/mi8GCkaft/QXEmenDJtNRkxoUfevr6V
q3fZfs7hzenNi/Fr/9iRopv+B7QLwVOKATNCwsaaPqlc2iPNcnKqPj6HpLvUzc/F
DldmFkTDdfOJ5fo2tMBXLc0u+QncVqyywC15ja8sYBwCadj09axSpng1Pz0N1sxz
FNKFJ2aNdGT1eFQQHeXAzIrAbnTjNnqeW8saAQ3dA+eskheBf1hQ1o56m3x3V4BK
h7Dz5izecXaHsXAkyQJ7zMoag+Qj5wjlSPcai8kjq7K6fmNaOABiaTCAb/GWbW/U
mv3xrHq1WrWbtFXFQzUATSuR/rLxbiFn2ILHnT9E1rxFkypqVCImZJ5Gtu0xLsX3
4R0MJCk1d8vgzXfRCrmAzNqLav2TSn4CAKQvlYf9j6GUlWQ0hMLoy0UN5HpF8WqM
wRdNihvZDOgtjk5hijppuWOxfk9aD95TbDxpbXAIpdN9VIP6Ui3lRAQsmxdOGZgu
4OoUG+QP44wVPgM7uhqC7ijy1BWQLAaL5RvjupL2qpL0ewnw09p3DEsoehJCXXx4
NJ4nwNL9OArz3f4r7g5Tkw67sEUZ1UTifw9GIHN0viXvvHIDuPvqhW3WI8Ozk2WW
8Rqdf+4Yxc2pfnJbI8Rl/k4NvR/79i7og6JzfZsBGLizfLvox9vYaWPVgxtyb4J4
j7XIy0Tlgz1mEGbWZxfLHa3fXCuiWpA7OPZYluyLm5q1fpcYS/0iLb1FlIr5YB2U
395kQQU1t1v5iRaziGoOSGmzMcn7H6bCicx6J9G9HRUiy9W9bNe0pRbp9Kz0xf65
18fqIk/LeDBz+2HQc6kRlI1wksSSj3S7NziMVOaI4QWtAExeCdBySrl4rY8ZdIBM
5RM/jd12syGpANIbFH3ViSHT6WSuJIRTAZ09BHRiZcpb3siFBUUqtjKhpBM7BGvN
eexjXWAY1T6/2b4dN4mWmNrbkQAAEWLvwsKxmGwE3Srhr3bN8Wj6NY881DzWKbuf
Zhbffh25d5cOF0uoL/tWFsoHtYSGeTUn+9qoqy4t9dWIlG3Fby5uqyorBCtqb38N
R71T60Sq5vR/difSJ+MYguK8BnYYViz4dpdnBg18jqMszMsHMgBiRvGKnYdAEkik
BbnoxTS/AIfDdp/AUSiX9PdHGlPQcYBH4yUI4XBEiY04oxKnAwcPpGxxt1sU99na
dILj0ram15OBYzICnqSXLTSwnQPZDtjpYPe6B6xJBV34sO+i7JDprLw3qReEooM6
IhKbZLIsyobgagzBm/HGAIiX0gvMLNklkelNSGAEUJnf360o4Esaq6Ed5noQSIMX
OXwnVGv0h0cUt/j8KnpkYTiRPg8v8EsoqsQ9BJ8XVDWy/jQL+V0AMztDHZhuM6on
fac9XpqiIsggPN3entYUJH6t82K5LZ5S11wNMFh/0Mc1uxYOa2mZyns5WlSpAkvP
6l87Q6iQiCWb+rECe8BlAY9tJsjK/tujE+bs0ooSJVh8rQjg08TTKH4XGIwOGtfj
8xyhl5F3LF/C7jMv4f3LS9GRszD5JVVSyxzzIofBTCoadJrHz+xTaiFJX6Gba5Ak
XR+IXNAs10u5YuKbDapEK14Y/9U/YaWUori01x5zcg9XvKRHIHogPup3Xd9rJD/t
qmKTQyTmTuJEiG0Sg+ct84rQYRBwK5uHTpAQvPIRUXjOqwS+iS1PIeKBJKBArMPk
Lh/FqzZITo3uRUF7I351+aiaxsTDbYBlFwJYVbykAcjT1Mv4cx4Tz5Lu+OF/noQY
I/J1Q1Wd1cAezmZlBA6j55pWMdTVw2JhXScQ9y0spvt4qVP574P6isVvMbld9Hg9
5CAKbMk/mbf0NmP0zd5QUiZG4btW6I3FRNzu5wzqXo9AOsclwDvbaKdozDf0IKQ/
Gdgzh8iJMGQ8iwhtG6WJyyjcyuCtp+VfIXxpvX1qPJ742yywG3vfIZdgcm3PI7FT
QD1tyUU3idZYQEPVWv48EJk+zbfmeNTErsILucLqh8Rl9IYtcCSwoL5/63aLLVAp
1tkk/aFw+25r2TR199eB1pJYA5Eou4DAT1sK+u0PkNcv+LFjQPTNm6p1yu3PYbPd
GxkdYCaN9n5CY5FEIy6OuaLdRBLdY1Jw8anhvhgqfm/HDgteNbI4smqlWO2phcKd
M6SngnIR5xW5OIIavVcxw7ja/1+HGwpYAQ0SXg0eotKtuMC+i8WupIQV4HuuP669
51GZ7WpCpd1aBiGCKv6HmY4N8tMQXVzYSKTHcOVLDUEZdypYsuq2R8ZsU2xE56Pc
VSxGErlr9MwVRpITKii5by0lvF2SklxKawGUWAcicQ/Sebn9Uhnc9gFF/900xV4D
7KfIJd8nDWhjA0hiJ7WJHNouugUL/ZgWDKJdZ0Y1d+rhuC90GoaXpEhQvBglyZKI
/cNYIlxGA88Oizdr+nlGqHrsWzME5y2mFjmaAqX7+AFK8XL+nNcOcR3CF1aKPPrp
0ojx5m+giXKkgysZ6tUZBkRYTkfbuFrK9dY8fVFaLVZ5MW4eEW+N4i3qCRn+C6Zy
Vv569vVX9OoFydcoAxORFJOrc3F4LLhAnNl6MkJMC+I6LJ3ha6HJ+0ZMtTlcyqbp
esIl1HzbivaCmXkG6t+DlmQCEm1TYfWoXKdx4XH4GtCw5h6it99W2Z1omYIJwHxX
tkpKV1Cj0881lxZZ0yajzI5/ZkJ+RFjNxsM9LGVCQX/wzrRvsgg3cr8vqaE0/pI6
PCw5jJIN/bCEkHcSYLCGR3Drvy/Pv2kQ/IpOPTgRSUqFjpSaW8fJCxQKRY4mNgBj
4s5iD1R3ckE6jiUbzn/sQO6U0x+X/0QrjtQWt38VEh/CgKPDMJFJuJr218kxXjLw
tAVB7IOp+aRqMAQ3bM1y2C5bUKoWjQGDW+vJz3m2CR6047ulYN4JHgxgrGuJJF/8
woCpQKYYzFVq3bvOyxBFrX0GcOEYzEOjlrcoYZ1GGooqVy8MXjUgfZDcKvjFsZGT
GFEMYVkXM9ZXAvbRBdl2NI8UYPaAtAP+Cwl6nAZyzUgMBy+1wEecOlAD+bvJ1oDq
xH8svmTiGOkpFECBNCQXaNq8jtBDQbvlSna+mgiCFo5dXVpcwUPJiuJtb6yxvsDg
4THX3DHsGKXhE26uRPhzlqbYCSXO24s1eHe6RhdcfsjQPJEpOvrTTwjWCAwJ7+pH
x3Q9f2cva5ZaRsGz8ly+XtmtiCimQV29KPStGcwJ8g51PDMxguCJN4HS1t590/qQ
B1ffHYMKp5l2QjCHyZ1gDkt4WYD7HTnRP50dAxjy23ZBNjWtumz70bI2ZrDQMe9O
hzMfWe8jEjVcd0iog0moO81E4fDzeC+JjpDbh203QbrhsKhWfRzxHoSoIXy16SMb
8A5S4OmE2ATGQ/nmg8DMh3Fhg16btZFIAzGQtJVhbsb+sOURrnhscxHHK1dZPqDs
Ba/dwaFHTHLaDHSgYOyzM181Txm8azVYJmjQ+7Cl6RDgVCjyTnxYi9Onq55U3RHD
yqRwZiANiUpEtDTz1Sz4J2UZfU2nLLLHwUYssUFZ+3Y7kxSGEPkVy/0Aiwl9wbWd
T+LG2YKTylfq610flZYwodhTR/+opSDKTS7at5v9c1lCN+fEjMyJ9NkmZj0ABiwB
lTyRglHtct4buILjpbURag7iOgLX8V1Olyitzx3ai/i1TzWdiC2qf/6G5nSQtxgq
E2Rq3wuYlvrHxnfZLWUhSeE4j35Erap/EcDRD7CMUw1WsVyRRBrYAsD3refzgr9i
2BQHEFpSpL6bGrO/8+u4DRlrK6zRE5SksNMFtt5ubSH3YiCy+OjrrwZOvZrvmBJD
+zu2clIOpdv3n2/LtYHQ7xD5PsIAP0wvDc8SuHBUtFL+3b7Vd97UHck9Lv35cFi5
3MvKXoiq/A6kNLPzYn6YJfxw5G9owt/Ko34sL26KYBffDTgZx0yZc3ycOSo1tt7w
cRcH7dauhJQ01RtH6swkei+dSFxQIfQEO0jlugXRixtuVnF9S+EEwWrmt45rGYwF
o4JrdoxyrqJM912Luv2hhDf9z6jMQUijO+BQD/uS3p+75KBTWXDBwP8ZaGJehDmX
2t/enTfoXD/GVmmeZ5894S0WneHE8AOI7md4TMS4IZ861DX83zZ/rYhbG4+bFmDq
tHieo0QqZNM8hNyCNcNN2oR/5ImWHz+fMI6hrAyU0TisqluZaH9GMkW8KM6wBIjH
5UgpqUVm9hJt5LH+WdwJlZ1BiwBV4VkoCegNE5LEuMTTMAj+GHhtamgrLh3cskST
35enAGAIgvTWCnxgdkCsj1lt4hf83GrFIt1+TvBbNXFGgsGxhP5kSu6PPUo0Wk7p
MDTDLYtdrQFE37Nwsc4UFKE0GorpJpfAvUWmpZSY0U1JRx61Ag+kgW3I+nPvMF4B
n9hAN1jCUr4dULGOQGvaODEkmH0tSzlG8AQ6Ey/Ai11l09dpImm6+08MMu2NgnLk
4udTK/8+JNlSAVMuVI3YCWJKSwrhECHXkXHmtJwMXvlreitGhT1DPAsI4LgcW9uj
O9INSOcpYHzRz6r6cwscSTLpryS4AaWTcg26q6LroOu0BbtNZgMEGKfJmHfb9z0q
TmqaKyO5/hSXaEeb/8KKtZ29Iv9SymkaPrrs1LawlPrmMOxMBPzv8YD4C4U8XjWJ
ZsXNECL3vYOEtKdyTJEsSGNAl3VS+vvBT9xt/dau2pI+wOVuLz2g247gJvSltuI5
G1olAZDJ92kj968tSV+Jkp1GRWvNM611cvo54pORJ0CZ1d4OD1ieZI7kTcpqb3Mh
mM4yPop0Kk/BOKZ4YtCggOKWz6cHbX9cTJF4nuIygXu/1FHXER2p5s/YjLWN+uBW
0N0IDdHiHnX4FxsfzwiyCEfXiyU/V1YH6DD8qJIuIxcIAuWXiQNQIb7tHjGw3ftv
SCYRQ57tEzoid4rOJnRzm/8XZASAzFoYsM7rWrYgXuAPgmbYr64ac2zWwybk4QVI
I9B5JdSvjyZARFVPRFOEyGWpjdllLlrBCA/n9/ul6BaxkuOjaeX36yWSg1HP+fT+
BjexvZ6GMhNQS+wm7EfASgQb861kGjG7mEPO+CnK1spNd6EDZpxxwyFX13ax2p4d
PTo5AxbD7wmbUTPRDI/QfvMdRcj8AmycIgVdbp9/7+e1QsfXSNj+TQMvNOqoOKxH
dxGfSmUaL96ZdvE81Tkj4oeZurfoi607ObhG2hktVnnrEXef+YPM9rzPFzYeNLnL
5FyJ9yIsnwWAEHzFWYDCsYzmwcLjf/t7XBjIWkvp4Kzt/1942qqkWdP1miS+8YNL
m9fr4uFzPgX+foV4c0XerhnSzHXQvfIL0XMweokdueWgaHkr0mx5CmtAE5Rcyl3a
/I8WfBc3PDrLCMVcizgKUbxmMrj0eEjoZvadVmjzfCD3xI5dSYyY5DmGCKImH1x9
TQMPxZh10eDmpdWBFlkbWZ6+/bBdJm7fsDDYgAgvnezvs/3gsp1xKPdGZVlxStIo
T6M8XEmbFDZ8pTQxNlJYjGiuFjrCyAQdzXt6dxb/ELFtXxJJ1AGesrMGPorSHyZs
5sTajSXHg/UXTUxxw1kgiR/dPcdyIvfxEkPnJawKUDwEQb7ErPJS79VGmrCSoknH
+GsuV593K+mQZDqIdMEfvUbpT2wjbVCjE2tbUvShAzHjdsGUB27PIhz0lMoTy0Gu
3pBzv0U81QiTjkUAMZsj9NDHNmGZI3rhpn1/OVjUBFDTDt3VbdTTk5/xnYKEjfS8
/lrWq+QUfH2KP4/RjYvZcw4Z0xkGIY5ClJN39dwU7kwyAzFnlhm9IO+t+VJqA5zp
z5hoyMS9/EJ/CNx0DGq6/WJkIE4jl61l0HF+gebuUEBuc0Z6QKZoWhZm2sF4Z6kU
TjbpwYDyqk/KYkY5brIjSKGzF1gBvGPyEO5YqMNKFSChjzMDR2tHgxF4R7NYKwE4
QW2/vnoaPT74yZBM62+17zjqUsnyVz1Up1EQwZeApJQkHP6cOyHUFfGMf0cKvB9s
Z10QWglVgczPMJt+Hbe4r8jHk3QM6VBQyX0oJIPsUO3G1iv1d1e147gBprdZgFUF
RQw//564/wXzz3BaDuTEgIJsmuNyQhtpQeed0GStHXIgVSoENYHcMwUPI5tDrawl
VmZfJVeobRmilCu5F3q+y46j/yBGYazOnIUbL8oP99ei/Fr8GhWyPJ1OmYVivqPK
YhN4YW9D2IbuYS59QvEWKy+pbXRQN9o0SsNY9FoOYF5X9MJlVQ6kUBd9B85pNiyf
6iZjbJxRyOOF5TSL7i/fv/PIJeUUgs7YrCvkxwiwtxqvvAjwIgTp96Jrz9xCzP2U
1Jg96nvqiPjnLTGjMHyviejS46rC5Wqo9ZjRMG3/T9JKT7tZ0YeWAYolLD4p107t
KQfP8VqQ4YZYrlWBoL7/T/gLZg68W4vvAaUAelvwzkPU7q9Pyr94hTceh4rtqf0v
Heo6KbujBsP8A3UmYmNDqBjJCFvT+Sr9aDB+EkB7SFjmMUpTYjdBKbTNqm0wtZRl
Wb7GMMOW5FS8rYraZRMitdb2lVeGsCvrkvEDueP0h4qysCpxpAH5kPhnVnis/wZG
/xMB4oumN4fM8NbVlLef/92WRj7mdJtCoMifmRk3yMR2Nggwg6pnZd6/s4EtAlHs
35rAh9i6rHBOXJ1u4BAllslVp1j47tr6FWQgRiCU69n+CAR67syOs3Lo95iL3M5h
JWQ+vs6Vouv1DBzIn9JRnN0zoP8VVBo3R6ARVbO2E/Sjlf87sS6kmJIEuQbxlLjy
/Tr1rSt3gPQ7rtmn68NStnplrD1a/+YH9ObdnD6CV2/DoYjF1tC5rAnxaiSUghY9
4BY4O0hKz5PrfFdpBFlw+2y9sQ7iWzPBGhe3iL+x224dpCQiextkJpABmfOJKeJl
qfPmFbNRA2nE1Jz+10Hil44TvIjG77Kd3Se+avTtpaSqQDkPRG9yhj269P+63U25
4/bog+8sN5sD8SvJcxA18njYE/IDt6ceXdMdrijSfiBYKKKRnw//J9VkND05th9d
/XWFs2Bg9PUkV+ttNMkCODeewoI9KHgE4Y9MrZ85UkBiC9eMneR6kXyDDZS3hAjq
SY+Pd0Xkb9tnuplBLkA6AVAuRtVE+uPEwN/NjtKa2LiaXqkgEQKTb0avPbGn5LUf
rgzG4CmpOEgWc/qwB2Y1POhzPdHV3jDQi0IqRWdRCAZ+S+4xQ98ZGGR95P93UEMf
/xz+JM4LQyvXtajaVi90leFat2KUQgx6e8rzAHI9K37/XQTbBkPUInYTYPN4hbCV
Q/q4kvMgLCYw7chQuEa5uWCOY2MWzrUyil4ECNC5M3CQg/YnMVDP2cZtWBcZxTlM
HfySeKMuZwBw+f4BuPQ+yB4N261xOwbed8RhcfcOgslbNJdbdC5FuGo+BNuU+OoD
0Uf0k8HKeexYgRkAbmx/88Ano8DoQo+6ChJ9BtemTUh5SRdnfRNb9FxZPkO+mBz6
SMXziAGUd9a6LmPzkjjBEy0j2nWK/d7TGbuvpTDbMXPR47Q8MitSRfT7fIawRQwT
vKwIa9FBlotPXbSJPl5+oJtXCMlVq0p+E+LcD7jtk3Vu7f8nRb+L9qtzOGrDFRPO
2LMAt6LprtKaYrWNsXDaFOIXB/43QKGa+X8s3PwVwQowz0481bbPnIFcn7E52E/P
TIwc3IgWHMG8pzDTAO7eBQ==
`pragma protect end_protected
