// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kkWJj2mi5pSIwemIe0Qz32kHUG1yNILA8o1ELYAcz1Z4hozcVTdq8Cla+g5SAUiP
vOtpXWuBT2v9oQX1Acr6pF9DgvS4d57Op/h5+1VoKmzvxWp2g61shAyKVhAuGgUz
xtrfqpNip0FBUQXG6sSwzKjccu65WhwjRBL/jUJdNpQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20352)
ilKnx5uK/JyKHQ0/YMNsdcXehmQESlQ+5g4FWAUmdZiaAy16IROFgtHrXFlOKQyl
ddA7jR8PeQQwoGpu0VMCGcjFFiCuRFjc8Eey3aVa6vVV/Znv0H8JUhEwHVbzvFFt
W+P228Qv7T8g7VNWDY5MJZcEFm3q0aslQl1YocvWtX5W5QLjUpqmTLsgcyMvT/9O
SlOmrQN+K8bnaT/EKBZeaQ5hQcEjH3VnB8QJiM2c2wuC6HYxBOM6wu9VTyz1VDOf
0t4hKF1CZkVauz3pi9Rr7jPhrmDX9mN70arwwL0v92Fz/QeiF1T5HYyGcde6hFC3
+M8XiF9JrX6q2lP44JTzip1Tvy1R+64XBzPtREB5S9PaHcsRZL2Jf8KFzIY1v2Dn
zdAbaPd7RrpCMwMirnisxIDcoi1vJC0CDsVgnwyXFGSTIOR7wRPNkyu2+vooP3eD
vFpRa0IHoRarae0Kpn8agpYZRhpofkzc1IrQjG+33VeAUo5YXroKwN9RlIFBrjCN
eLM5LZ3vsJyfgIQx0pKm1GcS8khU3xEwH+ttVZpA1O0EIQYwna7CMVYEfrQwfA84
usJ2EAz57ZeW6TxCBhI4wM6LrDzsLnTEPxYQPivz9oo5/JwSwROdiLALTAiulVym
rOGHQaRaSXkQuoEv/+BjwRExUouFRj9gHugwHNUI3v5fNA/QOb24G0X9Rgl7gawO
UB3rk679mudwVMe8oL9IA5HwWUng5dfVc0zd/fUs7ChScOdia6Es5zBM5uTTJUzc
4Wk6JEIUOAoDVxTqj9z6OEePwNKHI5VfyTrw3wqVtu6WIMWLtVTGT/xwH9Rrhhnl
N6T0bRiKEsFAgREq9pcKU09tIdaDmLrruT293/fsPvo8AY2UMIMMK9vqkQ77DOD9
kVpj0p/puC2bp39EOskWJe+gBznep2ETgEQpeeGb6wvs75SAsJjJOGQ08Yd8aFJ2
WQ4sTpi0mkWWzsLcgTDO6HVU4hT94IWgnolet+f/MVdBfTmM0qpdAd7uNXkQ70kE
6jJEEDSe18G7jq7bq9Fm8kbnqDLQfuyhE0cTLZho+V2U0QZ8pmXAbSJpEu9UVzmz
+EVI5JId4EuMwNvLw7cRGPdcM26kVe9tL85ds8XSfq/EI5HljI0KgRCGwTm7Rv8I
u7224UEWQ3PDhESFkAAJHGrbcxQpYxmbG9ak++5W9XGEKgYxsBYUc/Zxh9RBS74U
rqqh+e+ewVM1nLl3+G04JYy4yQhdb8YCJFiu1QP2I5ti0zPFfcEyLoMDj4I2i+0a
HTRHazv7FWRYO0IofNtrX7c9vbHyuGZ4DEzTUyd/oxBCpeqw4S7azjNnS4a0hzfF
G5OL2aBZsk5ojSpJDwQaYQ/XohU73hEFcdh5bjkxTU8EqAMb83w+Crgb+i9azEWH
7FzmBt7D+NpgJ9tMn0rsEhG/xD+PC+1uT1hNkKQd9bnYNyftPgWGv8WdMN/V2Wb2
cgEpXKSF1shtDeBJx9aLwtGzCkSpGccxvae/QFiFJ23mUKUceB6z6qPJ1P5ZDnxL
/Wk66Jis9awT0+7ryUl9RUnCe1awy6CcHRdEqrB/1BKes6xm9ugy3KrQEPQfURNu
JFC+9gQRW3WT+6sq0f+QOFnfGvQ9bYsP+P1m/PND2WRq7nPrtBJBB8aieemJKIOd
B9vlxP6Z1e9/9vItEfVqCGX0VTn4Jx4gIklIT9aAM7cd6J7yd6Pa4EtU6gHAtD0u
LhNxsAGZuMdG0+urxDH/fJN5Lhu7SaogLc+jC4XqzEy+SQM1hI6/YA2pRJL1QPHd
KeKY6g5jizCEuMrGjaNuiKfmOpkPNiDlfU106Gt9pZtXVYbA+6ORX5n9gXhFrXTt
tr8m0+ETTBkPG6RuytoejxeDbtTi0oM4zwl6/69J1NA5GSSGUXQJfW118mLCoXq9
GLogqxFJzrZhZmmXMA7/wB3zQvjfGl4RWwPScvE+3OS1mu3WhbPdC5El7HGmfYlh
kmuAqO2LcVWceBV+/Bc+wrduskqNZ3Yf/MlgDbWw7ShY/nXZwbGQFmgxcAYG3ELX
ZiyC8potAc2/ono8LSpAWPoKi9/JF0Vnrzf/43e5pc4y/0cq+XzGdN6maBzl51zh
93XdexQhXQPXTg6o3J7qQczY3S/AD4+goCUg02VzaMuTl7oFAIOe1L+VR0gZjG3O
7JcFJs3L1QvAkzonOVnvKYN/x1JLvcGOPDf2ZQVL9KfjBQiuEiuz7pYMTWhFizmp
UzjfCgZu3kywSSFnDritsgik4ZEgS+kBSbnjpKM9IIHdtlMblFpmI1HTPMwiNIGr
Q5adIsISNTgfkZO6/rDg2SJLZ2zF0HzETnmMWwSIG5Dk708N1XurGepiJ/ymwFuF
RdYDzjTtIoAhOshDY/kynilxS6pD8Iba1yfjQa3zFHOvXwbd4mUmnKRkgCzn3gZW
nE1E5sfWJ1bF35iKZPMpRMAeeeQ5cW1aJ8PUIUubQZSq0w5rkQaMb7y5GbaHODAU
7Qn3LCHNt7iB7O2/3fIyUPvEEGeku9qkEKZtPTtDelVtXMp2Hf3OZbqTKy+n0Ops
7mxK4NOzHuccdYaCX+GLJjKbsQDPsu70ofZVmwrrSeWDci7i3/J8rGFVBpDcnB66
slNZnusg2IHk3iWX4h22nHMyo6yWIwIG5qAt2wP3rEM+4CDN3I2W12jqtekjv028
rfJZ45LAy47FsD0sNXQeOsUnwsBPRc9Uxi1joXQZzpc4GZ4M5UG+1G6STZax2CRt
XqIQKaNIoV+RpGt0U9OvuH66fmbJxa8vDnB+46pqgyAS9lAlOA32OelFzlPnErOS
V00b1L7BdvKa8MkH/M1D2e0O/0Dhs8c13mhm11wo4xQmRf1qAoC+O4SQCOKyiIyj
rLcK1mzbeNcCm3FDBB5UHUSkdzz7TA7DGtATRmKHgjZY+pRNTN2NPXmogTn8sn/e
YUJ/4lrRCcdbLrqNSMg05/4zFVML6PFQmX5T8YoZtxuhrwXYXGX69BfsefzWSHah
h4Wy/YFL3yKHTb8qnIaSN/21tChvouIIlcTy1aPxvSORi6JRhYFa6qdPxNTDnoGd
U4NNW9soSzJ0lL+lUh1LgThBvvmGrmKi5p4u6ppm6UjXcwEfcNFOPJc8r001AEDH
+OWWb8y/p/Kf/q9Dc0439fP34MbYudfzlrJv9lHGZQzYhI9NThAQosyKwO1Jbihc
0H51s3+6r/oMaDfdCgzAmVtLXH1ciQoiXmJxBn+w6BvkaNeSBuhPFtXqo8WrzRV3
iNr+5l1BTC18KXwmWHFFOs51HLNy272lTb94qSZw/g5CETT8kGsxXNaZLmS5xWFo
Z71LK6cAGt5bvXzZUUv/0cr0o8sX7ryBZGV3Dxr0/SU9UZ7S10s7uDjQLD+El5G1
PpOSkc9gHKQqnfOMzjIy4PWMXBGv2ka5CUvycdzC+H52yhqWvNLC3FSJdv1dOYgX
/nB6t4NDT7LBsF0gNN5IpYlbzMPFwGs6zbdAPJvj3/0rAttE18UZTHxBFFHN0jro
E5w2AmVJTQ7hAM+DqJ4ObrvUMVMzU6m/i2gfvd8mW+ph+W9XrUvHUc11MphG21rH
oSfZB+ndOImxT6sWs2ycNORz0Da/sVDRj8IPb5oEefyxodo028eeEw3xzyZrGAeC
p3CMVJDqfCGQqZ3ZmS3V2yVHQcy2rgeVbdviNels0GSv94V8GdgUH7MlVKBzaGwT
ZRR3hqa+R+DqVaylWUnKHBW4RD+TNTgwEE8kjO0d85TRO78bqqq8zNx5yDRJlel1
NVYw7qjYqAQM0367AfidOdPGt0PfiSYbis2ObgG893LYVVQK2dchgAwvus0CVqw1
jvYICsv+qoMSp2mgPDxMAewjmJIlo0ll80+pHL92CH7s+ryJ4nVZiM5B92VuzVmp
Drv8jPWwqCu/wSecOu1I2A3qc+2KPayAqgx2/xFsehYL1NHAWCTHcKRNaCPR3CRD
hiO3jgwS3+yJ1SToLCEuqmnkq7sNZYBSHz09uGx6+uBXCycIqvo6vy6siZIg9iYx
otrmPIw6mEy7fGn22r7/K5K4dzj2Hfo5BOwU10EFzvovtlNC9TyQlluMp+59QuS7
Za90sM83tK2RnaZ34B0NsLxjSEUS/5ZrPaTl1Z8D28RbKsdXcRzglMsk6FYW33AF
UvYmylLop24896snuNmRfQmyLtfi2OK0sax1FF1OJhrtk80OAsxRegDGqdKvQI9V
n0i6rpSnO1HfvT1cETdgryyIHjO7YjRFxFzlNPZRYe1zeZcPcpRt/tPJzDFlzHtK
2IRNOYTvsXL9d79JP1BN8t6OP4zk9jQL/OoCVQt0ZIYU6pJ5ty/UEj2vvN+rwgGl
tzgMP1fdYbNK023DAkR9NSwSQ7RoN0wM7Vxa67xeqdoVwkjGvUqZlc+ZthaVusKj
1cOq3odBtM6oZEq4dDdY3hp6WiWPBff0rals0x/aPhN2mKf5rNq309ydCeKzltVg
c9hTcKcMJ94DDccBzwgqn0eYUBet8oXx0MZvuHmfLxX2eyXvZnsBhyU1eAdJnllS
zRvvdVQEbp6pTrdexAnsMDjuK+8m3zwIUTI0VLQ/mxLi3ialc3R3lP7/VUV+vPNu
Pn1BQ+9L8SxOdt5vm9DlLKGZk+YtLr1/1vVDVO7O7pA5ttv+IQSaOXEifYf8URKb
AWFAoovo27iR3G7Fe5v2avhT/4SG8/rryH7/d+GX6OfKDnJuQeyacK4K+r5D5gLr
W+ZZhDRBx8iHzNT4z4u+VLHJxTw6M6bPvSHOHhQMQjSJEXgA1lScKk+1pv+gydYC
k/lhw/IzagvhV/SWb9BmP6qHAlJW3dUhHO73D5klt+m2uYLHry20/rOTwzx/7bCr
ocIDB8BimpYhyxMsUHlSTFyB33TSbg6UBA0GTQor+li7gGTxatkAz9qggg7PMvEo
igeB5fvRTOHzqrcRV/XMLCnvPewBR+/b12yAEfF8tzRkvehvQM6r8FyLVq8Sdu9t
gIyL/AYjJT0A4Qq2jmN2tPDvw4bX8HNt+Gu/FHbfwVjv8HA+StTfNZwR1/wrjYlI
RilKpoxEe6Td+49/SRphiAyfkAwk3kQioVv3bzerUttVcDAY/P8rkINetqPO5gQr
auR1girMWc3Ne5mMFCewfBjE+xJ5tS2+3Nep16R8B1BNaAuJ0G3d+jG0F7WRNUdT
1Kg16/uHs8wbmB+Yk+mlu/fHPQovxfZnEgdNYs+HuKiRSAVN2AI8ecXvqGurVjdB
MftTzEv7d2dDmIgpB7luxzyXBGOq7MdKRODPncHNSID4w//Ogl1l8afRVS4IhtBi
hmGH070yku5/2eRFc5moKIVUTIWmGw9YCFntxdz4uSi4KlK+oLZeIZZbd4xE0aQN
lE/wATY+uDvx7MJ2PFlFaOdqxOMSDMHjAi9KcY5/FINSF6wQS202CuN0lymqZ4jw
mA53S4Prf5LrILaKxP5ppGVfclMux92bQlI2B2cTsw7eFmYhjG/Mxc0BeCadGIDR
+9A264yit4YaZkjH6MRq/b5uetq9K/8T4v3vvYi29z8sQ2wwBbTdFbZB7NoaATmp
hkPYVZ42ax4ylNKxzkjBY4Yq3ddadwGwV4wvQGcb5pjuDw3w7n5CdI7gb05XuH3P
QAWbiLpQttljMtKDiLvimSCvmHoc+2kHHW/S7pqXr0VMQ30pfBJejC01ilzfKuZU
Gw4e8LXHl708oiTMVT+X1RWTGI7siIro4bH6l6NdhkSJ4KQrqPJt1UvMKYwH1zzv
A7eWaWaPAZviPj8/JuWvp/XZZrlYHPRjp5cE55erWa/5KG7sRvGueVqj9UC/ogOn
WL7zpe9gS9CDA67NCMX40JG+JSpjze9oKBAxyEqxT3KeUzcR9ZKb5lJZZOI92XOn
rxviETCdmNRu5yZd/gQBFAQWfUPRTg/U2bHhtuG8DHqVtzg1KAhcR5th97xMDGOt
4n2j3a8v8SV4QUHS1tRQ61rEZa+idv6yhVSXxVyDCiFnx75OiVljbmnm7gTAHxXs
MiyIERHg+ghnmwFjTHKd1rtJKt7oyFZRFNBQuS0oKh1ttdeFVCpEFzWnihHiyiDE
2nyaYbyqwRnod80A2iqDkapUoNy+Eh3KSidlBTcsm+BhYKd6x5yepTCy+X4e4F08
q4IujQbL7bSDjGHSSNQbLgb2aaZ822PpdPsMwv8iv934ecZOD9yHA+3YrwFwAOhl
79W+mJyBJFIaAxByLGBATBXn4h2BhmXOHuldhd4KeRSS6wBqfr8hBrJ7rU70CkUz
qNOi9+J9CxIkN0sJCi314qjY4S43FiGqN1RAk6MH1V0kkOT99zgO9snZ/iyZPPsK
+bX6zKD0XMgaPw+uEyNnP31hvUA2XeyzCnjjQyHX3dIzucuWY2Y0+UZMfxhbtH6G
2XjfEck9iMmmwFXMTgcBjIU/vCiy9EYBcYFe6+xRI0OOIk+ndZrojt5gyPoPmJoL
rFxwcXA0OutbsDJ2gqMkf9IBxXixF8NoFooGJX5lxoCoUJxYjBAwsUm7Wlusxe7d
CxtsnyLLHNLfmF6MaP9uoEfBvwnyqHFP6Hy/97uIaxhiC+O6j3BnCPvzRId1BEpG
X6IhZ8WZmYWvBnheI1RZRH0Cw9MG2NCpk/8oGhHO9JrkAWZiqpXpPtSfn+VXnCPP
tWHg2TpJIi/1FmsA/Slvs31WQZLd6q1PwQ1Cs94T3J5F1DuKXbhCE43szmxZlfB3
zeNzw1D6FIl24qNj/ZjnNTBaesySJryk73mS+CcQs00SAwYj23zsjzHjrgtRcpVi
d1mY+F/5ZVXrrm2Xq2rkOTyeqmDC++TOllwqRw4CJPHMP1zkJTExObP8JFtumAxe
TwR8qffcZF8O0WiZ/tcutelUSdbWSAMbLemTT+nA6U90m1Gsx5RCbWvAX3YEUZks
xjJr+j0wEM182Q43rGNOKgW0UIhx2P3wTXYlb0Pme5AsdHxJ5QIEyxP3jJLmdfKs
efc6UJMXKmX98n8URJPGf1nXUgGL0GCVTjGIdDHtHtx5761uiLUENEzWXw1KvE8n
zi0WMKAI54ONZbCKbx+IpwXq4wRO4ffzrhHxJJ6N698ggNC9ZqomMJF+aFwpXsLc
ln0nbUxD4mRCKzAkfjk1BAO+rXsiJymFcwmfiIqzaZ5UCpBSC6nHVW+3U+V3TOv7
vlkDZcHoTRzcFRLcho8u3ftaS8iHf7tOaM6EfkUJ2Jv0tc6vtJpdfAocxvWIhP9K
0dSXAU5atB5W2YFoE2haH6nNr90NIeOzB14CvtGB9tYoGPGtjdoY6ksKrQ8AQwQr
lw5bf1ULA0vguUKkp1FWWfA6udHdgSCr6KY452QpHHrSfeXUyDr8XPpwqilUiV7S
oqSjF9mq87nbeuhDdXNR0NOPuMyXJMNzJ/R/Q3Oiv53qHDWhTwpCItvWvMQLWy2j
SVG8zfeR9Gc8sW3OXx0DTmVAiwA7MuM7bsmopuDc8oF8s/C1eESy5a5aBCRiZgKM
ik8J745hyT/47Woy88vpwLGm4FYp6lL42fvzQQOYAX3xyoUsrq0s2WKuBUlNhL4Y
Xut0Y+KuX3VGe3iXCIQiQQYp3Qq9PAQOUvzQbkRDU/soAUCE6OmCAECP5YnBf/Tr
18kyGANPiPMON/WwT80Qm9pRxn7gdzpwHGk+iS/uxkJJ5wqehlCKvMR54JWaDxye
CDjpwUNJL9P3dMEJjnrq0LBPVtA0ole2wVLjjOvqatPTc0YVWI6cYeetWpk6E7fL
Cc1LB8rIYoRLrjbQkcV7JwPxeN6ymr6wU89AebN305um8y/F4fAuVv5RU67mqHjc
iYPuousPnWFYWIcLsrnaY6Ee40DhzJZWTU9WLVyCYYUnB4xNse+y8tZhFVcK7UdT
Oj83r1q/s7mducUc+CpschN18gGPD+ksL7qUJ10OKgOwziaObPPPR3veVcZgE+ez
coBkLLnvfelRwH1SOzcDEaYQQWh04CD3U2J52s5Cr2KsHVoeFXYOvggeYVWlur/z
OxsdJZNvftJ7CKnHOfq341KpbshP7aVGWvFBV3ACHY2797Ge7gM9rpW7f3QDKwKh
ObO24k3v3kSPpbg5hldTExqlByKowMqSHSWOumjxROaWJpIMALpGa4sqwvTizNWY
xOf5ixI2gH3PuVtJrhbo0w9DF/KenJKbpeWDmTWjUqPU7LO3VD+LcxrQknLdbXd+
rNEqfqpepYPUHa5sJSqsxEPuG513+RzKFq7grc/tZSsosYB4UnWQac4OHr19wlwd
X+kL96R3jydqNvUIG12kaw9ULNb4gmmCLZvVj49jDNa4WMKJqDsMpOpEcaPEtBZt
csYvbIHVFiOheKTJnqeiXrbtbI8ddOlZPoZsCenX2UE05wFYn13jXzDcM22os3mU
T7iekiGCarr/ZHmT/9WyEr1uwA//Q4kR9nnCdLOnV3q2iXfHX93dinTdlG9GjtI0
Ka1PrPhVODiPGp9xkPe4grEPQ7Vm8yIaTA3pHoq1LXRM6Ttcb2KI17c/N98Ns06+
+OwN/HSN6phFZ1jJXUwU/FCVUFCdTlCpAk529MVLi5a4PQVZ6N0ByJUsjrNllQZu
vJR7iyEtXARMyPLrc/+GkWzhBIG7OjjF5wZ970hI4TJi6YJDqiTe5AtgGYGS3I48
N5pQ9o2KahKoQYC6QgXOveHfk5oKzbL2cA4U7RqqYLwvS5I+U4Wq+o+ra5cse1iK
vByTHKuNJNgWwy0ID8yvHDipBvDIrWqkrgT44AzGbQ1bau3iEtG+1ElCuRcX4gaw
hAEUKKM0LgqLHD5BbFLBY8VlCQJ9uSvd+ry+6hrT9NMVZAwyJDBs8nXWhj7f4kaY
llAaVTSefVj9YFAwwhWeFf0euvr9wgNKDd+KRio6BAjMUQJo/BkoU8spL3ucpCXW
9I9BcrSPzOjqlCjNsZnXLwNt0hiZz67ul662w3LJNTHmrqpCaFLUb8vUKh1VKU34
FFEUssqjir3RTGA0z0qzmCJvtcNn8Nx07S8uYBbhi0wg29MrkQy2oE08DrtaBt47
SrqR9Z6wu6/ZRQkJTsQ6Udk/IfX0ODnA4RIaZN8N+XY8aj9/sZqEvRS7DhJ5luFf
Mwf5CC3NDnhFZT+XqgsBD51ziE9cPryz5h1loYhcEqnURyE4UX46eS9hafvsF+yG
uhMp914ZmJPWzNFhguRXJOiWcq/JAA4Jn3GVaVVQ8R8jsaGRvbKNgs8cHwSusL0b
IqOCP2lNMYJ408TG4vYkrJHZ7xWC7gwkEDs24pKnBNy5US3q82mvzUrdSlhECYQM
4y88OcnChwuIy9ywuyyr7LD9S+gtlQFvItaQpykcd2TB+JXK1H1Ml3s635zVETXu
yRsYkmJPGgyqVhjNytNII4mJuKeYXN4EUR7/vCf1b+K84mYQFHOpcPqZgyXLLUeL
AZt8/oLP1T9C3kutcnS2VNtQ6S/5bZcW3lSACFVGJGQJ5alAea7Aeu+v3Lrt4HIo
PiSbnffu7wo+Oqj771v+K7DBHkY8U6UKdIfYyqFkDq+6k6tIn9ityC0Y46xFeggk
ulao14b32WrYAcpeOQhgyio8mHRkw2IdOmgITSpenrm2o4efMVczkdoGhAOuXT2p
AWNk34jfMKa1iP5Gfk3hhkaJFlrz6U84bEU4XYZ5LiERpHpWCMFeqxFWy6zkQYzG
RfugUOoOAvbLzKlgFsQfgauKRuRUJzs2ysimHLY8z7No0nlAUdBYXjTOt/XjeRdv
uGvEmq5/NM2IQGL/rmnZsN0VaR6kz8aPNRw4dySU2ElvUo9lUsAMm/LG+PtA/7Mm
N+ExbAXX8VKdiwbevmpcxvVD3eNu9dZlpliOkCW0nVcWlodwBHq4TVmtiYN3AlBl
3cPPaGzHwEHQmz8wG4fRsquYVWHVpqZy3k2rAswcdmLcZF6gBuHTdT5FCBzzZq2r
eCOkr0Iwado0SK7vwNzJ0svQdWl6KsyHCPY5GOgCKHjwF8LB6tTa4TwJhzaSdQC5
tTx8z4ELO8Xwy/6stRbAO7mBtRzSDJs3DhxPSsyRLE3NhN9OVAHekBxycP+EsIoV
BI0pgP/13+vJJuHNstoTM++ZY8qUUpqFZgEqcFnFuM9f8k2wfVUKwD6pwmgx3gH3
yC7h5R9IlVlc5AhjaXNF/NryZ5b3TGFRDzNvALHgD63dBMM6F6CZ3STlqj9LXoVF
qYuw7kf0MM4yQfKXRalH1MNoV6wi2XXycb2ujyvdvDDPwQzHT8hDNBG83XXWiUjp
6lDnGxr7Tq6DzvGuMn3P+cob2E/ZwwYpSXA9X4Ays3cPkl1EzehRpXouiZcy/T0t
2FqEbIbNB5fV/Ef3l/Az7sW/iEgh3+ha+6S2hMpfGPwcqPuNVCjyrhCejOTL/jIW
06ek/mZJdLB7gWzN4hN4dRtcjfib443rxI10tskIQFIxU4cIXutbShQ4OpKawRjq
O7vGu0SgDYFQ7zMer7sFmje374iA+N1mVPTMXh+SrDrNEK8A9xK/0PS4TbWC+KmA
RwY+OpQWjIkb7f1gho0KFVECy7WcJeLUNGmpckMdJvjTy5G2dA2UN5J4JDPvxktp
GwtyvhTSM78J1SaWysdNvjk1Kv86LxmHIyEKIlDCCjy9/xr2kGANKdpyuZXYehtw
KB5161D0wfJvdfGjtUYfYAJCqN+nfO5iXyHeIrXDX67GjajVdoAzTDE+VWIVGp0g
2I13WPGA2g0mIPqn7aI3dbCKzS2VtQVyol/NAY5TOrNOvG5w8fW5yVc8Vz4+cWPH
Ovueg6kSA8ak8+RxZO0Jl0B+HzTPl5aJyNvN+0v4fTKcgwT7IrXdhLEpBVr362WR
N58gLRcfaQXnR3h6bA3lg4JsfRicz8ot4QFz661cqi9JDQOE7M+0MyAQAesUTsg1
6Zh1tjPN8R/2gVWFhT3sDTfUt9CZmPBAl3T7aFffMlIJSWlBtw8XdlaaCW7+Y0oe
fQOz9pAC0jxZQF1Kv5FfzH56wGUuUhB0tPQ2TfXSLZwlB9Ac3dGmkUO3a7yU6YS0
eTYbbIGvPdR7XkhDcPOx76WkM+pnmVMaWSmtNjeRpSfOrIYrQGe4eQZsWuwPNaon
nrmJCVVMlHb+QxNek4iXJX+NVzL/m250qWROYrg3dys72iiX63eg3zY5tcpFDPjg
l8bhwjgFWd/7u0hg+QTl0dR3yVfrMDnfgQzIzgf+8hcg/FUfhyG6bIbJZpiCqGxb
A3cwerubWAhrgrjlF84sIZAf1/A61zh/iavtLYjRgNM0KUtIdqKaRQSILFQOgJ/X
nkvX46cQWdkloMujjfEefFyO/8ZMbt1/ADcz0m47fxUYFldef1nKIrAJUG0euKSy
ymvlic2yUGAvPyeGehTazAUC+C9j/pikoD15+ucUqOH+68avvzmw7WbE+vvMHG9n
sb3XzA3a+8K3aj56gmK+v3b6siSIiT8eEG8LqDG4URQvVkTFjRf+t33ZWTNoZRHB
g1ob2m4tHktSSLlDnf4PZWcPXw93tNbM0rCVqWEHb6fmKpWkM8w+LuxUwdooYXqi
pT1QWZmCVIVieNkx7t8/51AJix1tdKDiudHKyuSgxTUmh0+E3+e/eUiKWl4AsO7d
gRg6sjHnMf+wDYdWpAYGZKNILc/4glbTyFnjqUiaottwrPFtLWrrpUyMbo9qnsaP
dCA68Ka6BkFVPO6WMIqBe/7Vr4+dzEG6TQo0j03yVsZmAWVog4S4qCI77HtnBogO
Dw+01pI+90AjoiyklZax1/Roc2ta+2i6w+mzn1MeHDvxBxDJVNZMns8CeVUlyt3j
tVYMTNBTYLcoI1EAMkcCHKz9UQLsVlh8yuroFIv7wgUwnMSLzqyG7DoW3/Q0sxtc
dLs4mRCXb40wd8b20Xr3K57BZi63/VKZ7ozbGSl76lamJrJCJQN0Nzt8cmSRLVUN
wxLYtM0GaUSinku7Q9nhvXs8mE5GbbQ56VojvZzYHJ4nl77Aj0H573z91XfN/+S6
xAsLOxFIKiZDI3P8woFiH/kv40CixngwBzsStJzu8L5P4idz2wsVhiOprdCKnvCJ
ncXZqLybBOs69HTLQWEK2vcDvi8IeENSG6NGX5KAgShgxw3FwYnr/frUe2bsnUsG
ZR/8ZC446tsua2nYEPt6Q54BIxt5teQw2eSqZYbbLNswf3SkU5RGlJBPxHwYXNpx
aFFlTaEFMTRbBJtwDusqCnmyeYvpWR7B2TRg0IL/eN/Qa6EK1bt/ZPdxPiv3HsxB
+sbUdpP6SXNB+waXVmJ4E2JjWKsxa1soVK9cadQepfOg/Oopoik9NOHkGiCPnZGO
ycr1YX345NMF8v6Q7HVwd1qyWwIt3Mso8tKVzqy2wta+IluPOwbovasPXp8sejbe
paagyYnYFECUOILUnug1GXyqZLsDhb5ncTDUClWvLQNKau6RjA1OegkA0S4w/Rgs
tAq2LM7yPhE6Y3hlJfqgH0hyWunJP6p6ffHKRCEqIHLerP24QNHYEYrbUgRxha8W
TMPPwung6HJMudxlGElte53nOEQ2eh75vWxmFZSWU/1ThjVLGSaEPl2VaNJXONb8
q32+C6floUj7+Js9JIvA+8kcZGJduWXhqE2A1+hNHTARKzJwZOxWgTOTUwrbvK9o
H45GyAj+v6qt8XEfpc+QmpMdNo4jqSRm9D3n2jxv2EZvxACbAmboRgqrEDQl9Sr2
lGfLRBV7YSuK2lsVe398+NT/bZcxS6El9Jv8nIdL0rDacv3G7f0NI62bNBTqA9+l
TgD7FzU2EXYuNWUY6zdNODiyxW9bykw+6voYnApUY4PLvTRDfOpWl66BJqvW2wgp
Zr6tKGDwR3j6uRSlclAqTBBTVzfVELdbcM7/1q0KKjOAuHuCxvKvN1MqCOz0cOKV
N0upZCQB5nq3r8r2lkumgotb6t3WnMis+PgRkl7ECzLUFOfeGdeCadZoIZOjtMFz
C+xmWqw9J1m7BCHTE7ejZxdomtjtlMESezWn516AybePcONcDF3z8sT49kSbFT8R
JZNTFPyhEnUxgxcaqy1dD5nIXVlUQ2hp4naEjB/f20By6idsKFKd67XNQfTyRjRi
J+p4f8Jxc9bTD2CzcuWEZ9zoAIGoWfGnCZPYYbrZ7hQPWYApe6Hb7wZR9wIwkk2I
SlxnoX8tLSFcoHn/yrhohmMabe6P4bPt5Zp9X7swqS0uJ2AIASDZ8LcrPij6bPqJ
EEaj/b6LRENdvxPHUTtHKyM+R7AlQFlE2vvNJvps//SkuyWZUt+SXOgKZ78qnCgo
nnCINhu2TS9E/XtXjZxbj+PvWRnMqhjeHHycUP3T49n4833qucYF/hjtQkiKKHr1
Ny6ymiJjmMTeZpJcf5BC5CLqbPcBkCGYQdP9JSzwEsaZldGSbV4urUQgzpeR4NBS
CKP9qpKZzJvf/vDd8vEDrBJFdEnqloUYEw/Nh6F+nc1cWh3y9/0ht6KPSn0PTfzj
4yv2fWMCoCg+mvbZklgipLGvQwed2bfdELmV5OLaY0Aclp51X8IFkC7Wfs0vrx1p
kqRlNrmWjHUSufrJrHcbjITIh2kY09l+w/9M3Cd6jAyI3ti3wni1c+5JUKbZjViJ
eUBDDqO4rX3CdbSlKgUb0HrF4Sbe1BJFnQQV1IQgGpW5EJg14gSNAjayjiSeL0Ob
FQ3Dj0m+e8y8SjcEph+1K7DfZIe64V7gMOf3WaqLz8qbt74WKPRKpLhflD8iPZ3U
jPfNLbqSuSy6uMsVFtD8iAkjPm3IkMnocwKVdVSiR580syGhOkT3OVktPpbrEZ3C
3HpzxPIdHEvi4M6huPn9DtEah1/Gy8ThVlWcaL0sHfAYQ3ok5QPDJh/SVzRc1fC4
n6vIpnTad9gKJ6glQNvfM5tmruCK6tNOQzJ49h72i0aBB54N36DhOMiNzULiAgcu
0mjTZUXXQG6Lg+SF4lXU6SPSXENP3cHoCj0pLF7vUoRy4bauTC5i0jWupfKwaYma
jI6B819iCl1Srhu1YPRHtIH1fLIrSPMa+WAjuxGgjLKviL1usxw6v24V7lA6bZl5
LnpW4coPvEcka635mcRQiw28sdUrqOZ5CdQLAGxV2NE2t6lJQnhNY/ZQICXf+h1W
chjr8skgM6GYdBK6/3ou2MZ42Hgp1HxWCxJPSP8Tzq+EgEJfwuAp4O0OotJR1f7w
crUgeOi1dNgQA6ywQQZfe3/6znmH2MyOjiC0HuTsu3h/mLFTsB9k4VITs2unKTHT
OZUa4Yez5UQOkutJdam6Vn2yOXBZMN73i3QYsmqO8VWarASV8iQgcXHJvd7OgKJO
0aXRDY7KuveQ0uByxawEhCZ4Ss4j0synUKsH6RrD6Dvrr1i1L5QzvqflRpyEK+5M
xJlMB1xfArqgeDX2mAR2Mba0F2P78+G4CkeGd0gJ28U3hi++J+lKTuNwQqt44XHf
QK70h3ub0cxF4EoKiAmH5YEZdZQKa14VRRzFZJT3D9fN+p61gMiA2wVYuP240gXg
EEYT06ULCt02d18Zo6WpuEFmfg3CIJ+dposCorQG4V/MFjcuOj9FxBlsxs8xzULg
UaP7PEBB7vgrJ2PAVcAGbJyWSgWuHf4CN7SllKDM3A9yH2Kwk/gZPqD3wZVQDk0U
gwe1PBSm9hY3gbag/OiER7OzsvM7/0r6J4vIMbjxn5LgvDhFOmrGwVuLNAEE1zam
Pe2D4dJqYwsWMWqTYWTEKJ1P2pPw3qgBQz2OrDcpKLQqVMtoLulw/Npj4rYI28q8
5UUZvKwExk7TRuG/c0r2/Iid/DUOXuVGIbYwuaA6eOwb6Dz06xTUiGNwEvm4IaIH
xOSDZTa4oNlaDlVD+7MMt8VE/HG2QX6Bia40QKCe9m5oyc2wmYm9KNHC97QmW74N
qRosW/ZEcqC3N0c9bhY+88b9+LMhK8UArJAOtL6+YGpd6dtC15GfslN5cE4CNyT6
AmACWLdL0ADGPS3nMDg+2wj+R3qTe/WSUOrha2ci2JO7W2FfWmMxYXPa69+1V4WQ
dhdHvfwGjBgj0Y5mb4m6y97a6pu2GDGFYFXWkmKyOgxCZJQmAi1rSItYGR+dkNo+
Fe8IZnGeZhuT3xxBHHtcqYXh1RRfZxlYNN278DapxmqgwLkVl1iy8ITS0hBgMbBl
7PysJFn5Y+ZrncsXmXP3XaG930sJVbOVA6NhZ9PCbyBnm2R63gYx9Yp8Gl93o3Sf
ZNDgK1R+bxIZhfJ5Q2lkRdMpRLpktr+yHghmq/k2RehL1UjvxHOKb4WalMTnGW9W
p5Dpi1GYjuKtw4j9YiasS8vgfHUw8hNTUBCEOqayuugyQka/VjTwE+YPK+qLHjEs
OBbRFpzc5uBELfM8KLZlDCP4wifmaiEMLybRPvXxf3R7QIG0AsgO6SgyNdAuJHoy
h6LKyOQNGbysDkT/krcWArwTcjh9Nr52Nknd9lEyjrucl/r0oC8GCT0R3XYqke4J
cYtmaMke8yeAntcJ1FS5lRyeuQjWWtehf6skpihJBoMppR3JQp6C0W3k2eYHdKx6
gM14XgBAQnIT96p6xJvY8ZCQLYGbAMd8W+DYv+WQSgJb5oLIbyXPThTNpOZDzxF9
NyXGcdkVztWZ572mAaTi77lpLX6HPxYwfLQbgX6Ekjk7jbJaCL3AasftDpP3ifiN
BiXdTicMULoUoYnE7eOv38c/qrrmfhDrktEi2G4aHZtr5+9iFUfnA2x5cUotCcQE
8mpi6Vx/STCJYYi3TF4VlVj5/4YZDk5yZ6zucA65wSmPacxGxyXsnqvK8QJoWF2i
PuaF4PkE3glMLgOb4bDkrVVFysMJ9mNRSOXkxxP/n9GjhKJZ5EPNvWeu1TsXETRZ
vlzadO2aXV8UmtgTPzaX/Eyvrgssj0zBmaYs8rrt2D039SJcSBIFcm8L6Cyazld9
U49BEpn8ssmsz3a5VUMJua/Bx44ilVvdb6KpGF7XvCpao7ByqfrMPRVW8fa7pQTk
+9BXhJ0pUmAbfTzeRywAHpK1C86Sobegum7MCQuBLYq6hYa5h8vgnc7GXFawSOAK
zXkCQcyzbwlUEgZbFhD9l6EHFFLkF+zZ24QLunwkTQibI7o62hbbitzEOpWIEwm4
P97lOL5zcRaUJ+f1YS8NJrocdaIEDW5VSDXF4i44QgsaKN/aQBDDlOh7vjQ7IbAj
2F+yfuKT09qnscqwi6aeNRQdqnoCoy+IvBg1o+IADR/9DnILbEO1g6ytZmUD1eHY
Kzf+FBcMb2RvisorPbHdrf3BN6BM17NSifCmPknKDBTxTDPnLpo+M6ySHg4PLIau
kmPzSexmLX7Y3R5MAGZB1suHg/xuilw8LByE19ge+GRqhLkqcHxYcKVg2AYt7LjP
CTXOt2KhcElKCCYDppc3HFt86K/5fe/nSmyuQc5TDQ4xeQFRg6+eu8/89BnM5pFa
rRkS58b/nAzJWPgfCCDwTd9OnXsUy3t8yESziZHmRTa6bSTrAOVoeaXPFI8SGBfy
HDDKE06G2pu7zHG5JteGBLAhK3XE55MjnkK8+I+VrWm1YF+O9zt9/qLPyIDbjoV1
B9vt7rinCLgD5esZFLOGC/G0skPNL2tK+1cgOEAbIWtlSKzmhBYFo/a5J1z0gQ7u
Ho1anvBeyfLxpy6jC441ye7ieArO7S9Wl7y4YOjPj6LCkDcwsyJOPyGB0A6bS4/1
ONcw6sy0IbSNwj5NkCLLzdOwghnpTrVUd4sk9B/YkYvnlf6uLJbITChHxJsEXAYZ
NMLfIrLERJuS/qykkbezMHX1peaLprW+ejwpvkg1qsoIz40+/yN6rU6a6WW+6QtA
6rkt2oGBkmKqzuchDBS2O3QwRTbWwsFwTlYzmCoLj6AxTjgRWJFiFsShds9jTXvM
yn+fOZ4KUjHx0ZGn0V3tELk7Uj7otFopoIDvre9M0UI4hWFWBmXeLD0VES55m/fg
yFjvNIKqTIIT7weNu8eFHOqdfr4otBsBpV/YZQ7YmoOQxIf8soH/tCHalYQ+4WCE
sVlEhQ95Laaeg67pR/Q6bt3hG6Knpw+jTK++nDiz2l/1yJM68UANUfX8tTi7YhZF
8QRYIo07XMfC1cTd6rNxw94UN2sncX0DodkuyTnBK315VUrQBYGcXNdEXuwx5jz2
cDbzFD7Ss/eXsFxenNZWCIzmsEgEkdQx/9psNmHDZOoqYsZPK1BpPxPes3X6scF+
LYgo995rZgsk5hJrVUpge/0fVIvZ1p2xtTP42/bhvwL/jmHA+eddiL3/rzjUCPWy
b8dfZQIgDvvGFWGNs5xfHFYLqr+JmrSXH+yLp5opPzkn4NZI76M3nXKi/C7kG1D+
LYqqxxF5TNVQxYDXLuSOG+oX1Wdztn0mFkl624KzrHJ+fSo3gX8Fkf2DOP2MBwP7
c1+BrZcSxM/SmPVzMMnpiD/jPkBzooof1SuuVNJYo1eVNGxToxNcln32/yfio0fi
qw8NEvLS3oGUPOQJgitvP9snYvUBjYk+Yueevs/eI2gmIrKRMW7LoANorVFc/nas
Ze/pHalVFvx0lUoiXRX0r7XTjIpzVbv1bVFTzqQG+a6j4ZKjERjTBrusdcAmqOm8
TI2hychJAJKx3jx+7lBTK8bD9DxTIdOJiX32jEHpos6SCqzwdOz7v/nN94tmwc6F
TuSgPcQY6jdTcnbMIDVMMeKamaUa21NhJbenPzcjAohgolrvhndWRlwwuxhcQNaT
37hm20LQHSrSu4Xflmgo5gCqFCZQL1EmHeLToZsQzHC1N0Z+Mqgm+pkjjNthlVwH
KIbYML4M3sSDHB0eikvGZLfYhtXZjMSsfiFag79fdhPNWxSibYUvXkrZ2TucQKEu
IzmOIfJvdWvKIPTYUDn0Wcx/2wBT310Tqr1XfZsxAV7RzmKxZ5shbfsRTahNtlcX
Lr6E/0YpxRtBKuotsv3CPd4ziS86dQFZE3gUhjiRmMnDdEN77Fa1+2j7bfhMvSuY
oQFCd51186/xvCkSopoqqzQrPAgQ7sQDTd0dfFvkej+Gv0xuP+0C513zEu1lTsiU
5brnRkUPzX0xiUTZ2mD8Iz/Xxwie31jLg3kda6ZObdX9Kzy3pj3UcsjyfzRnJqJ/
0uhht381E2oRX69WeBomdwPuHPiT1UVBTWkHQJBFfRbSLImvrFtiHrPgNKsJCY/7
wTvRfakJnjSoZiTJsm/xH7isi4vRZ4/1gAPyiqHSaUpOQhiOXkg5d8K0DKYJa+WE
BOYvbqdz6zy7AYRqcvVUIFvyWi5hUvrTG6Ke6vNXkoEjIdVDCQ/jfjEij6v5ozDx
W0qkFrDv+wU5X2jITAPHdQGlb9lRKN8cxJAKBjlQbSubvH34VeB2Ht+fh06ZfbZq
RTR9wr3RqJbalrilC8MKbkpSTeBpl85DiPJCKKHwTkqxlciuURhvaZC5M//FIi7m
Y8n2CuDkpACoPVS9Yis1uaUdRBVldXz2gycZlzVQTdpCYfHk8xHutpyKF94BIc+C
P7XGx3G+GrjIrKFIpo5YIxrMXeS8ed5vGmlGxUbkYHlqK5ComxPOhsJXw2rfm0ud
yBMk7T1BMiNnHFwfkB/uIQBIibKD5k+y0uORrVcb4ZPLbyi5sX0AJart6k1vcrZc
PsjxXbyH/gVsguiARNimuSfH6VsMjBEwGK5kf7kTEP/SqBIUjixJU8gzQSf0mN37
YFiCfUe+lRGQW2Dpinb6vGJespBTSms0buQFL8iK35QXuLnB4Rsmt2now2q3TOik
WCXB6qGkemznSDCsE3NHJZirNt5jHK/oC47mPfLhwe1UXlT4IOj84rVUGnb8hHC6
2OE/M084gWvs46KYqLpXw20nKZBCpDTWKItNdrjNKFHCPV3aQm9UAQ6J1NIBQ8wZ
ccRSZAV6ARNscOUoLrRfIGFAkuK9yOH1pIfJF4lN1yPwcLxHsUGGoQ3zTc5dTEDv
UHHTFHY/7JCvSM7LY72TmptZm5Mw+jJu6C68ELKfBJgy+jGtXn1U5X4AR3j3X10y
chewL6+pGOoLOb9RPiTqYET+ikx6+O7iRGWFPq3+WyJgkgDsKY+zCeoSir2YH16O
jXmnkvTEiHjXgKFgFOlZllcSf0CK3QIL3lwYLOQ+1lwVXw5rfsNmHa9IHbW739/n
1+yAAiqXVTGJphtkGUd+RCae3Q7ZlanBx6HT840uW9vKAy5os3XD5tYf7qajGsr2
vJTUCxjgB2EjjVcjmB1SzO+QMeWw0+RuGNIvW6AhnyHRRRGFnU9KTzBW+/uMNQNV
7ZlFgq9EGCB4BDGQEpAijW0SZCRn6T00nWoQpZDbPesV7Q2PCj3BMaGxFWRnFnx/
sgmgEceXcX/C6nzJD0e282LO2bATdaapTKiAG7z5H1ekN+OoxthMXXHn988A8fJK
unoQw+SDhBogIMnmpSTDf+qRuUEezrN/ZsnBcIGHs9AxLbuTpCn57YPNFES76U2Q
cTCtesIq3x1N+3qOsi81mvle+w7CmXMJ0vJeveAtkmTwPNKcAMaRAR0M1KzNYIja
CS4ZXucOBgwCkrCiWyW4CyGq7fnYZY/Vux4wfLbB5QFOM1P8YjQNsiqDhiV/TReM
OdeEJKJgU9lrrqlXJoVQt3RI4TpPeYBl8sRIjebtJmBJhYBrBFUVl893JDgQeAFO
QteuDi60AG8clfWZ/o02YZbGTyet8+g0YTZQzy3I4SXP3D7ILpnhV5Q+Fl3fTo5x
hg4+Nw3yGNd9oaFpLFgP3G1OQemtZ/PQP4aSgiCzc5MIYIz/5x3Yj2b3JqK0Hroi
mzg7eSbHJn/HertzgmRQm0HN3pcwFsWpgEsMzOFXpxcIBaI6nnzbLNKhaukiAg/E
PdAs6PqkE9709vlBuLjjEAknqHHXak3Qer2VQ0T+4in58UQBveWeIfq9HKR5PBmo
N3c3JM94d5f3jWke+i6jdUJBpEaEWaP0e1yZXJfa0FszUyKL6APDOUu7t1a5I09c
oewl4T+s+ysiftY+ObaaMukYieW+fdGwFQqg7uYaEXUn7AYViiIIm5UDSFVOEiVM
9KFPGH2ONNyoOUf4WOW/F7JZN8otnoIL/lok3X/eM0ddKj5nF2AwfIsKbmHYxfab
bJBtH2q/KFfNjQO235vULhOnJLViqpAiNAbArDWr2tCRShopJvUcD7aFKAJDSJHY
FvFnfu2EMvfz6QTInQZMbb+ODAmA+la6TCW8SZERibZdUvX2Zty3ZRzzqWFNlpKa
aZkFFeRSSY29/zgV4MCDfjRo4BCfmP3mxg62WoEQbVhWv1sIEhI3GdZGjlhOChiy
xwivU+GOA/zPomACLbKcXpnHnOxf40gYEay/5czWZz01+pwD7bWZqOjNoZQY93Ca
frf6Z6YfC0HYg3e91YHcwZOgf/6rD+W8tpLcCBAPd9TUNMY9x6NA19X+GU0SGYz1
/Zd0LTG+bst5QCVGV/W1eXGerBa+Gs8HaTT6+BdKaNrkguVK4BLJj/MN2RLZcPpj
MzGBMWbBKDri8V680DjtCRZWo/oCyD3xzFqtyJmv6KcDFPkLXIxheeJdzteOsc+t
bXJWyk6/f+GP29aHeIlu3yLzlDl+GSpd55Va46fpOnnFdHdIC7GvyCUnE8kxpCnQ
W/cQkreNHBE4KirTzNKYAeO741ITGhu+YHBrxu0lKlyAN9PH5NuT1Ww2b/o5sk9T
9ykyYx05l7gyI9Avqq5fjWyqlHRN8G0p3uyz+JgWVYKNvoxaMVoAV3ELD3T6xRba
Bxfgl2JICdfpyjZEP8i1br1T86nyD9YnQnd45qvpfBuea0Up274clclJ8JTRk5rD
OaK2vEmi1woSg+1bzfzxWRj07PQAtPQSskQTP3Y+I9Loe9XdefeN1CXn3fdPXYQh
cNvgR6SxfJduT/OtAOc1+RVPpv+cMDndTmAac1aToJGPV7FoetDfEMEyXIvZ7/mv
fRrb98UM1PJ9QKW1jQlapI/F95rOeDdmDXvv/eGlpERoPmI/gICs/4snXhegRm/I
PhMalzaztv5jtHBiksGXaGuTR5S1qZ4Vb06qSWJwVxJO3enmrXAvve3wmh0NYTV/
V/wHyJ10z/K4gUfO98ZJ33ZiOa0idNwgehCqrVJKc4S0+Jor9U/dw6W5uLOpJgjH
C9Ab6/2EH97CK6YZF4N5kMRtd/zT39CGtYwf8iVpc+dSGR90TouzXlZ+lWsYnORn
oVodXQYy5d4dtpyZoWVXvMT0KWkc6SlcCoBvuKtq6VzLGKWs2O6mj2zrWT7CkFnI
zRPJ4ATolZcwuqvLf1hbyk6m/imMJ/+M8m+I3ZQBsYlGCZaz6PaD+SrqfEVjCUok
LIPBTxKb4CIw+mjJSM/IuCAUsNlzBRDAobrwc6DvwFR9bvUnfwmSYRkx6gxoBnhO
jq1MnFKXj5tIGlpb4n4Ni3RfwUt616CIbzYtjPuBDHySHfiz7/sGy6tVfmmzJRjl
tGxoKdNgf1UPjSWhgfOuGH4MIMrrRHzcDy7IT/Tl4mQWPTamhMbia64Bji5bCez1
NqlQ6C7pdFdI4YLi1llkkXLwfp3stujXRFqERHS/5EMl+Mg+XPk5aB0Cv9rFJwJd
tB579KkBPvwnKcpC9OpOzqo/lIOy1/rOQAUmo5DWnhjh8EtCd3t5oaPP0RrabSuq
gR/ZYueGSMeGnQ/UjKyRlPoGzOs3w8kQwfIZ+ATM7JXlnqOqDVo74yajOnTqUkxH
B6paBDNxN4pUIdZEYvFsNhE3/BL4RfGe5KltfofyoyyEWbEOaCm598hz5HEIthGr
bUHLb3ULVbDm0SoDeTnd0lR9WJwacY9GCdkrOzZoqLfaZZkl2VfNF90v7ftWtdD1
Bp6SDEuLsPaEFsSQO/V0owsMZCTU6iUNMRR831QLvvbFOjP7kIvaGx43ECHld/qU
pfHLwrBfW/0f4VDye4hOMTX9pyyiFGps4rid9vl5DucoHqxcEp+J6trzEU3QqI67
NmbAwVzEJjl6NI9Pd52hou2t3dZVCpp9Bg8U07LRgrkgVZGmOdAa2Sq5jn0X8/Er
3VnRwmkOCMvoXxL8f7vhq20KVGvLqRSvX3jk3yWANyXxp22JApa9Kbm8R2IAAO/Q
IwExGK6sNFighJNtMUHbb5rHUlFSMhw4hXsX6oO68JqdgPWQKbmevFdrghxUyrB0
HyVqa0Zp7RSm6kF6k8fvaLb6U3Tc0u6ZpmE1iOphhRGNEDGiu/FmzHBuVx8C9H3w
1cs+cTzvJVyn+rreFhxh8u3TZvratMV3mXOOzOS7FVbXVa3k1eAS9Oe1To85ixTO
Q5i9SkFj2VAGAvnB8GQn1d4F1cJ6IDgmiKGCMBJideqkC43lPHI6+RtJhtuCGbX/
elQzYMKaC95w4A5vF/HU/tTIM/CeIuWycGMwFFvVR0Vy3hRDR9JdvHHALkklG8cM
aKOFTDnReSmLlAKmuxdQW8PeXm0ahO31iWQTNVctOr7rmm0YYVpHe/Qi80RFLO+v
TOdPHVW+CWAzHx2ZwcMz6d1/xixSCNvb2BpTncDmqP36r75J9iKeRW7Og4VjcFWa
XUDB82CpwGCW+i91OFmiWP3mP48cn0RvJJ+WegH/2vRaD5YAsnMOV3G3UnlnCO42
hpevT02IsVLPcdwNTgXO2/dmV+0n787MOdU6nib95hs8Mwr8pB+XeJ4x5xPyJ969
eP7unQ87OTMCpvdTPNQ+xG+2ECecBEFY8zomJhReRVrTR3WLo3YXXORRFqnrxmF5
qCvLGacnyZyVdRN579IAEsUW8spt+TMxTLlwN9DrkulalGpmtdfzr/lfZjHs1pjU
vt9NbSUAWlMD7b5+TLNLwe/3e1c0hmxIf4KeA3eew2xl9DgKIjRnsW2MzACt2FUq
JSvaH6cfEq7EMxeiO4nGG1YeFsnf4NdgHFXKP3gLc9+SIfnhysGvjgZwtsR5HH1/
8SfdxPY2FfyEs5woxjUmatC0I96bfEuNgdfRLoblon9Lg1MJLgxPMxhbUY2Kpeoa
B2D+/FnvHQccgFnnZNW+k28Zk/lK4W/ThASqcra9ABpIFI3PKGuqD9gsFUYd3LPE
5bCRAtMhwCjFNbXZxFcW8Yzi3KkLOIM/oa9KlExv7DTXzebxOUJjt+sIWOtPz6Xi
K9VW2fahkZIsjCwa5tHn/7uqfi6bQ2crCUkmuRouONPuQqYnfl9d9vtI4NdGuqYr
T03pk8jKQjCqyV+rhgs+hn6Vs6wnvYhIriWVDVuA98MNDlsgUIT+Q6MmIzFXz5W/
g4n8sU6FDXRHWTDi7MLnUot7fOxHVSwwdHWULPJ5EHFOIFqPp5eCcUA46UcMo6Yn
HNU6ozqOPzxLwc8z8FN74K6D5iso4kYD8xUknDv9STOrLecT7OzY4D/BrIImdwvh
8bkjrgJsS2xuappRLFCN50JnCQgo9L0IsOGhqN+JNdAPO60fxHS9G2SwEZa9Ikzo
xinMDcJ68e9BrcCeWU0upSbUhOBFQdDMShouDIgY/G06ZBp1CvEXDKd9ExqOKwuC
ySlJwijEd28jJNY1Ipw2bZWdkRVPqEJJIm/c627xmIxHYQu0RTBH/5TFfZccpeV2
4X1WbBGaaSR1+1hDF2Z9aTDyoL+s7wZSflE9cABacfoxxms3L1/HgtjANHMiG4KD
QVW+HA41SsRxF5H8iru8lORiW8K0zVDXtpfcazHXh2t4OEUxEo9aKMdbvmMrET9k
7kluc0jZAmv5wW5CRrvFkdOGLs+Pd4kuywuSe4alApiKhZz71VCZljPcs49BdZbQ
zFEB7MqXZFXQjGlgT5JNBC243iO4/VEby/CDAPmnTerFZ19TrOIErpaO/R/c1W7y
1d43YeILv9h4Zdc5/GgP7bQXq3/dL5P70gpzuAhKcuAehqX35v/2R0eMnifHI67x
axBW20gJghu8on8Eb0mU4hPhPPj66k8PrQaeFmbOCZ46xbdomG1uE1Fa4wTliKTG
K/VAWAUG9tlkNsipUUNYxBeT/BNeCnGWpfe1LsHidhzZmM4Xz3HJ2YNbiJEn6kXp
53svWWLuUJ7yANKD7Ryo1QAdBBW4zsR81YcpGjg03b/ZTEJ15lKlXTQbRqEnrNZS
fuSV2rVe64EWyblJ2svHLsQQoaFjGPYN4jqfpbtkSMcrE19PVzay3C+utr2WggMR
9HEHbivIIywjDUJ6qtRdTYX2si67j+yPSbta2gOTDtE41YCEFCY9xsCtfKE/bBG3
+F0AdmY21ft0GbpupPg7meD+LGJtzBYOBqluf+lSqIe1f5VHao47FbKK4yZh9ymy
z6irAFk1sF9gabbUsODwDkGMO2893JF30EDHcMc2S5AqpgNGSwMFgjgQFK21rIkD
VpDtm7FS0zRN63EYGKVTkjxTJypzAMZ65bnPC4TedpE++gK0PuLxxzIf3sA28NCg
Y9E2Z6YFWj+bhsUgBsvS2kKXX6ta7X8A2KHn+5iEBCTRhA46SAMOtyjDkUs3+/Sh
Xz3FfpeH36+xlBWrp7degfJF6VJbHjbt74MS0UpKN9absmnthHzG5mleJhLIb9Xk
JAAcWzHVfLeC/yo82GllM+oGWfG40yDbJvCtYiItA8Ooalp4Tn+B70BmZtILrZ38
nJQ20f6Z0kLmD2r21lkzY9Lclac7NWPnQGUTdHruASwkXBXOdhiFLErrPr/7cSB0
8fYPtDVGmXklPXJC2ldLaQ0sbXnoBOYeXCuajkRKUyVrVn4lxogoiQ3NuJwvWv2i
7bp82RxrgwGstSNtbpm6iNkqZ54iBdxYZ+/LnxVTojo9jOSscpOY3OL6U6xHGXnS
qk4iNhSwqnFQiYep+k8etCrP1AOSjcFaPBgqLImE/xGaqDIvf8Ep4vrPLtbNnTz/
+3w5MV7Apnr+yAL9fil3+XC7XvjgFpWC6gqd4FVOGJh0CQA4CqvT27iUNHxs1vcb
jD2NdtVyt9dJDxNQrFPnUu0HrBZdUQ4nh7ourgKQ3W5mRi+0EDhUT4HFdWAVan2C
c/KOaXq8u7Fg7plpOzpLXsTYoqxlxxg7CPo+rY1Z5q1mtad5VVtu4WO2s6bxPz3y
9+/GT+XPxYPtVt35eOjTip4NqHmCxCVYQJYmaNNsAYdHiHN9AXADNgFImiK8483w
Yp0AzQwgySkH/07rYvg5oJUUVgJxFHD+b3Do7aU8hXMm962dSSj4A3z6B6DhOno4
QG2bmXcnLR6pcEGlQZnFOVqtbzm1VqTU3k4mmIcN1Im8NMMiPNCASpOTJ5Ks1djG
lXG6NfwkA76SwjxWYrivIlPWOqxU9S9b+aZYRjiMSJXZMeEs4AU6r2XqDX2Hy4pL
FBSbS3O1WoH//81ONOdCA0ZaREfZnt8+OaWtWKuayr8qhn8yU1/isvuEE3Iw1B2Q
LcCabjOcnTaNS4Ex4QgYZ9tOuW0xGXMeo6SbumSgL7dn7LIGtKQXQWKI7FMAQHD8
DuQP4FdB2/B38aSwtAx/uuI+CYUv0cxvFjK40/Cqy7ktm6VhdeOTApYa1QJOpAWG
+VZ/6LEDlg4392+vlSKohuHbgKyi+EBNCQdKIMgBYQRvE0dtoA8UtFD3zxauoQND
7ITYZDr6xXRuzYSQVgasEMN/X+tcB7+BEHpO2i9g6Dft+9Q5dtfiNaQFi86X9CUE
w2EtygQpDAjn+jcEtOnAMHElsIY2Hz726pka7GTyo63KVCyiTGeFadNWb0wJEk2v
/rfE2hDz4kdx5ygZQJ+GHLKH762GsbTWy4MU83RlEr2s/zoSysIWpjWhZSDG9d9v
ppC6i9mT4CCtM84wmWhEI3ne9qhrhYrG4BIj+ow9rI6Ip88fgvZxr1iofRqtdbbA
qSlFstsrDH9sL15Oa9lWyzYhG5AsZtSFG8+BbNneYBK6MGsV/ckGtzTo4ZT4Hco4
k2163QBO9iI0wmRnZDQ/06TkDERz7pou7NmGm38vdgmEs3FHlalFUInjh51MakJz
hMbTnXkOesbLhlou2P7MQZYvy6xFlQORq3Cu//VFNlmiOeXjaBN0LuyFFUlXkTVV
XSh0GrKvyi9qK73LLPjT07DdODxC1og3kW9CQgARKpzrdf9EVM+pFzvuNhaQ79gW
/JaXmoiHA6tT+xjoFtkxmeu83x19HmoNr6uU1n203Y2hhwl77TLRjl0IAtlpvhOZ
+bvtxYu/Uwoz+wuxyDxN1bL4wvzlf1Pb2qxMHWMSiucyYXHSBXeC2TGdrFFlZsXV
/1pLz3eS2JA6AYDUR4bNhXtSvME9eOV9IPTcrNussFbh+wyAz45IyYDuVPSD5UPt
fU21lmi2HyUZdoruGIbv5ySPNyq6rw1GJf3QhXWC/Zh4W1iHD39zD+05iEAzrreO
8kMVaja8V9Jn0IH7B0Eu9P0xW9gyO9P5TdTJChDxrw792J/uOVzohxdGgilhsYjq
eo24IczvBHiReTBCQID9gVOl7xu/XWXYlks64qgPQbtX9T3FTNkAOeKpSdlk7Q3Q
bZKGJMcres/WjNEuMfc65gxyvwU75PUJGziZe3L63XKtskE2EtsMLuhyc5Z2T1IT
cyDmm1UhOUH/rO/PnrltDO/4xkOZaWqahjsDO/uteScaOHOhsQb1frQi35umYMwG
uVK3faeF4aGU1ZCoJSLCEwMDCti+4rN0FoA1L7/YXq4tL17k963UN1WvYRL8tI/h
LTFIlo2MbwhAr/IZzSaxOA2AcsLCFaEokJBfaG0EKxXQLc7wqFNVKUwTlPbrSu+D
MfyXD6iL3g5f5srdXc+VirbcaU0cyCgrPU6z8uKrKf0QH+gG9JOXhGq23XWtr++n
SD07nSHdcGY8WhBN5Wyf7iUV6QLzWmGVOixSXxhitLZvjYHolVX6B80gD3RJIYcr
2w0TI9nyBNOMukgzuhe24tIrkHAP7hQBgIo2cE1BOPGidXnf9BLf75ShpuTCL5lx
W5Da4D3zIILDrJU1QOUOWJRUsh7+AtXYrawv36I2xhz8LHk+6dPr8JRg/AbqhyUq
/llaHVuKxg02xyDRCEcVnM7aJ1985MrxVDpvvCqxE7A2GKWe6ny90vKXlE2D200b
Ddczx/xG8VOdQ63T4YaHxX9hMenlG7+pLv2OfjPO7M83cTFfgELn2wpwT5BIs4tF
qj9VJIG79cUfr2Al8ty8nEno9TvUuTbLMvsnsQdp8AeVWvRxAlida/65UepoKIE2
tT6bFWyRcylYYWm8VwQdVlN7IRt66HEArfi4Zw+uIsq4v/XJQyKb66sOf+56BdvT
`pragma protect end_protected
