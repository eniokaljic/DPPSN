-- megafunction wizard: %10GBASE-R PHY v16.1%
-- GENERATION: XML
-- phy_10gbaser.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity phy_10gbaser is
	port (
		pll_ref_clk          : in  std_logic                      := '0';             --        pll_ref_clk.clk
		xgmii_rx_clk         : out std_logic;                                         --       xgmii_rx_clk.clk
		rx_block_lock        : out std_logic_vector(3 downto 0);                      --      rx_block_lock.export
		rx_hi_ber            : out std_logic_vector(3 downto 0);                      --          rx_hi_ber.export
		tx_ready             : out std_logic;                                         --           tx_ready.export
		xgmii_tx_clk         : in  std_logic                      := '0';             --       xgmii_tx_clk.clk
		rx_ready             : out std_logic;                                         --           rx_ready.export
		rx_data_ready        : out std_logic_vector(3 downto 0);                      --      rx_data_ready.export
		xgmii_rx_dc_0        : out std_logic_vector(71 downto 0);                     --      xgmii_rx_dc_0.data
		rx_serial_data_0     : in  std_logic                      := '0';             --   rx_serial_data_0.export
		xgmii_rx_dc_1        : out std_logic_vector(71 downto 0);                     --      xgmii_rx_dc_1.data
		rx_serial_data_1     : in  std_logic                      := '0';             --   rx_serial_data_1.export
		xgmii_rx_dc_2        : out std_logic_vector(71 downto 0);                     --      xgmii_rx_dc_2.data
		rx_serial_data_2     : in  std_logic                      := '0';             --   rx_serial_data_2.export
		xgmii_rx_dc_3        : out std_logic_vector(71 downto 0);                     --      xgmii_rx_dc_3.data
		rx_serial_data_3     : in  std_logic                      := '0';             --   rx_serial_data_3.export
		xgmii_tx_dc_0        : in  std_logic_vector(71 downto 0)  := (others => '0'); --      xgmii_tx_dc_0.data
		tx_serial_data_0     : out std_logic_vector(0 downto 0);                      --   tx_serial_data_0.export
		xgmii_tx_dc_1        : in  std_logic_vector(71 downto 0)  := (others => '0'); --      xgmii_tx_dc_1.data
		tx_serial_data_1     : out std_logic_vector(0 downto 0);                      --   tx_serial_data_1.export
		xgmii_tx_dc_2        : in  std_logic_vector(71 downto 0)  := (others => '0'); --      xgmii_tx_dc_2.data
		tx_serial_data_2     : out std_logic_vector(0 downto 0);                      --   tx_serial_data_2.export
		xgmii_tx_dc_3        : in  std_logic_vector(71 downto 0)  := (others => '0'); --      xgmii_tx_dc_3.data
		tx_serial_data_3     : out std_logic_vector(0 downto 0);                      --   tx_serial_data_3.export
		reconfig_from_xcvr   : out std_logic_vector(367 downto 0);                    -- reconfig_from_xcvr.reconfig_from_xcvr
		reconfig_to_xcvr     : in  std_logic_vector(559 downto 0) := (others => '0'); --   reconfig_to_xcvr.reconfig_to_xcvr
		phy_mgmt_clk         : in  std_logic                      := '0';             --       phy_mgmt_clk.clk
		phy_mgmt_clk_reset   : in  std_logic                      := '0';             -- phy_mgmt_clk_reset.reset
		phy_mgmt_address     : in  std_logic_vector(8 downto 0)   := (others => '0'); --           phy_mgmt.address
		phy_mgmt_read        : in  std_logic                      := '0';             --                   .read
		phy_mgmt_readdata    : out std_logic_vector(31 downto 0);                     --                   .readdata
		phy_mgmt_write       : in  std_logic                      := '0';             --                   .write
		phy_mgmt_writedata   : in  std_logic_vector(31 downto 0)  := (others => '0'); --                   .writedata
		phy_mgmt_waitrequest : out std_logic                                          --                   .waitrequest
	);
end entity phy_10gbaser;

architecture rtl of phy_10gbaser is
	component altera_xcvr_10gbaser is
		generic (
			device_family            : string  := "";
			num_channels             : integer := 1;
			operation_mode           : string  := "duplex";
			external_pma_ctrl_config : integer := 0;
			control_pin_out          : integer := 0;
			recovered_clk_out        : integer := 0;
			pll_locked_out           : integer := 0;
			ref_clk_freq             : string  := "644.53125 MHz";
			pma_mode                 : integer := 40;
			pll_type                 : string  := "AUTO";
			starting_channel_number  : integer := 0;
			reconfig_interfaces      : integer := 1;
			rx_use_coreclk           : integer := 0;
			embedded_reset           : integer := 1;
			latadj                   : integer := 0;
			high_precision_latadj    : integer := 1;
			tx_termination           : string  := "OCT_100_OHMS";
			tx_vod_selection         : integer := 7;
			tx_preemp_pretap         : integer := 0;
			tx_preemp_pretap_inv     : integer := 0;
			tx_preemp_tap_1          : integer := 15;
			tx_preemp_tap_2          : integer := 0;
			tx_preemp_tap_2_inv      : integer := 0;
			rx_common_mode           : string  := "0.82v";
			rx_termination           : string  := "OCT_100_OHMS";
			rx_eq_dc_gain            : integer := 0;
			rx_eq_ctrl               : integer := 0;
			mgmt_clk_in_mhz          : integer := 150
		);
		port (
			pll_ref_clk          : in  std_logic                      := 'X';             -- clk
			xgmii_rx_clk         : out std_logic;                                         -- clk
			rx_block_lock        : out std_logic_vector(3 downto 0);                      -- export
			rx_hi_ber            : out std_logic_vector(3 downto 0);                      -- export
			tx_ready             : out std_logic;                                         -- export
			xgmii_tx_clk         : in  std_logic                      := 'X';             -- clk
			rx_ready             : out std_logic;                                         -- export
			rx_data_ready        : out std_logic_vector(3 downto 0);                      -- export
			xgmii_rx_dc          : out std_logic_vector(287 downto 0);                    -- data
			rx_serial_data       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			xgmii_tx_dc          : in  std_logic_vector(287 downto 0) := (others => 'X'); -- data
			tx_serial_data       : out std_logic_vector(3 downto 0);                      -- export
			reconfig_from_xcvr   : out std_logic_vector(367 downto 0);                    -- reconfig_from_xcvr
			reconfig_to_xcvr     : in  std_logic_vector(559 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			phy_mgmt_clk         : in  std_logic                      := 'X';             -- clk
			phy_mgmt_clk_reset   : in  std_logic                      := 'X';             -- reset
			phy_mgmt_address     : in  std_logic_vector(8 downto 0)   := (others => 'X'); -- address
			phy_mgmt_read        : in  std_logic                      := 'X';             -- read
			phy_mgmt_readdata    : out std_logic_vector(31 downto 0);                     -- readdata
			phy_mgmt_write       : in  std_logic                      := 'X';             -- write
			phy_mgmt_writedata   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			phy_mgmt_waitrequest : out std_logic;                                         -- waitrequest
			rx_recovered_clk     : out std_logic_vector(3 downto 0);                      -- export
			rx_coreclkin         : in  std_logic                      := 'X';             -- export
			pll_locked           : out std_logic;                                         -- export
			gxb_pdn              : in  std_logic                      := 'X';             -- export
			pll_pdn              : in  std_logic                      := 'X';             -- export
			cal_blk_pdn          : in  std_logic                      := 'X';             -- export
			cal_blk_clk          : in  std_logic                      := 'X';             -- export
			tx_digitalreset      : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			tx_analogreset       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			tx_cal_busy          : out std_logic_vector(3 downto 0);                      -- export
			pll_powerdown        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			rx_digitalreset      : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			rx_analogreset       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- export
			rx_cal_busy          : out std_logic_vector(3 downto 0);                      -- export
			rx_is_lockedtodata   : out std_logic_vector(3 downto 0);                      -- export
			rx_latency_adj       : out std_logic_vector(63 downto 0);                     -- export
			tx_latency_adj       : out std_logic_vector(63 downto 0)                      -- export
		);
	end component altera_xcvr_10gbaser;

	signal phy_10gbaser_inst_tx_serial_data : std_logic_vector(3 downto 0);   -- port fragment
	signal phy_10gbaser_inst_xgmii_rx_dc    : std_logic_vector(287 downto 0); -- port fragment

begin

	phy_10gbaser_inst : component altera_xcvr_10gbaser
		generic map (
			device_family            => "Stratix V",
			num_channels             => 4,
			operation_mode           => "duplex",
			external_pma_ctrl_config => 0,
			control_pin_out          => 1,
			recovered_clk_out        => 0,
			pll_locked_out           => 0,
			ref_clk_freq             => "322.265625 MHz",
			pma_mode                 => 40,
			pll_type                 => "CMU",
			starting_channel_number  => 0,
			reconfig_interfaces      => 8,
			rx_use_coreclk           => 0,
			embedded_reset           => 1,
			latadj                   => 0,
			high_precision_latadj    => 1,
			tx_termination           => "OCT_100_OHMS",
			tx_vod_selection         => 7,
			tx_preemp_pretap         => 0,
			tx_preemp_pretap_inv     => 0,
			tx_preemp_tap_1          => 15,
			tx_preemp_tap_2          => 0,
			tx_preemp_tap_2_inv      => 0,
			rx_common_mode           => "0.82v",
			rx_termination           => "OCT_100_OHMS",
			rx_eq_dc_gain            => 0,
			rx_eq_ctrl               => 0,
			mgmt_clk_in_mhz          => 150
		)
		port map (
			pll_ref_clk                 => pll_ref_clk,                                   --        pll_ref_clk.clk
			xgmii_rx_clk                => xgmii_rx_clk,                                  --       xgmii_rx_clk.clk
			rx_block_lock               => rx_block_lock,                                 --      rx_block_lock.export
			rx_hi_ber                   => rx_hi_ber,                                     --          rx_hi_ber.export
			tx_ready                    => tx_ready,                                      --           tx_ready.export
			xgmii_tx_clk                => xgmii_tx_clk,                                  --       xgmii_tx_clk.clk
			rx_ready                    => rx_ready,                                      --           rx_ready.export
			rx_data_ready               => rx_data_ready,                                 --      rx_data_ready.export
			xgmii_rx_dc(71 downto 0)    => phy_10gbaser_inst_xgmii_rx_dc(71 downto 0),    --      xgmii_rx_dc_0.data
			xgmii_rx_dc(143 downto 72)  => phy_10gbaser_inst_xgmii_rx_dc(143 downto 72),  --                   .data
			xgmii_rx_dc(215 downto 144) => phy_10gbaser_inst_xgmii_rx_dc(215 downto 144), --                   .data
			xgmii_rx_dc(287 downto 216) => phy_10gbaser_inst_xgmii_rx_dc(287 downto 216), --                   .data
			rx_serial_data(0)           => rx_serial_data_0,                              --   rx_serial_data_0.export
			rx_serial_data(1)           => rx_serial_data_1,                              --                   .export
			rx_serial_data(2)           => rx_serial_data_2,                              --                   .export
			rx_serial_data(3)           => rx_serial_data_3,                              --                   .export
			xgmii_tx_dc(71 downto 0)    => xgmii_tx_dc_0(71 downto 0),                    --      xgmii_tx_dc_0.data
			xgmii_tx_dc(143 downto 72)  => xgmii_tx_dc_1(71 downto 0),                    --                   .data
			xgmii_tx_dc(215 downto 144) => xgmii_tx_dc_2(71 downto 0),                    --                   .data
			xgmii_tx_dc(287 downto 216) => xgmii_tx_dc_3(71 downto 0),                    --                   .data
			tx_serial_data(0)           => phy_10gbaser_inst_tx_serial_data(0),           --   tx_serial_data_0.export
			tx_serial_data(1)           => phy_10gbaser_inst_tx_serial_data(1),           --                   .export
			tx_serial_data(2)           => phy_10gbaser_inst_tx_serial_data(2),           --                   .export
			tx_serial_data(3)           => phy_10gbaser_inst_tx_serial_data(3),           --                   .export
			reconfig_from_xcvr          => reconfig_from_xcvr,                            -- reconfig_from_xcvr.reconfig_from_xcvr
			reconfig_to_xcvr            => reconfig_to_xcvr,                              --   reconfig_to_xcvr.reconfig_to_xcvr
			phy_mgmt_clk                => phy_mgmt_clk,                                  --       phy_mgmt_clk.clk
			phy_mgmt_clk_reset          => phy_mgmt_clk_reset,                            -- phy_mgmt_clk_reset.reset
			phy_mgmt_address            => phy_mgmt_address,                              --           phy_mgmt.address
			phy_mgmt_read               => phy_mgmt_read,                                 --                   .read
			phy_mgmt_readdata           => phy_mgmt_readdata,                             --                   .readdata
			phy_mgmt_write              => phy_mgmt_write,                                --                   .write
			phy_mgmt_writedata          => phy_mgmt_writedata,                            --                   .writedata
			phy_mgmt_waitrequest        => phy_mgmt_waitrequest,                          --                   .waitrequest
			rx_recovered_clk            => open,                                          --        (terminated)
			rx_coreclkin                => '0',                                           --        (terminated)
			pll_locked                  => open,                                          --        (terminated)
			gxb_pdn                     => '0',                                           --        (terminated)
			pll_pdn                     => '0',                                           --        (terminated)
			cal_blk_pdn                 => '0',                                           --        (terminated)
			cal_blk_clk                 => '0',                                           --        (terminated)
			tx_digitalreset             => "0000",                                        --        (terminated)
			tx_analogreset              => "0000",                                        --        (terminated)
			tx_cal_busy                 => open,                                          --        (terminated)
			pll_powerdown               => "0000",                                        --        (terminated)
			rx_digitalreset             => "0000",                                        --        (terminated)
			rx_analogreset              => "0000",                                        --        (terminated)
			rx_cal_busy                 => open,                                          --        (terminated)
			rx_is_lockedtodata          => open,                                          --        (terminated)
			rx_latency_adj              => open,                                          --        (terminated)
			tx_latency_adj              => open                                           --        (terminated)
		);

	xgmii_rx_dc_0 <= phy_10gbaser_inst_xgmii_rx_dc(71 downto 0);

	xgmii_rx_dc_1 <= phy_10gbaser_inst_xgmii_rx_dc(143 downto 72);

	tx_serial_data_3 <= phy_10gbaser_inst_tx_serial_data(3 downto 3);

	xgmii_rx_dc_2 <= phy_10gbaser_inst_xgmii_rx_dc(215 downto 144);

	tx_serial_data_2 <= phy_10gbaser_inst_tx_serial_data(2 downto 2);

	tx_serial_data_0 <= phy_10gbaser_inst_tx_serial_data(0 downto 0);

	xgmii_rx_dc_3 <= phy_10gbaser_inst_xgmii_rx_dc(287 downto 216);

	tx_serial_data_1 <= phy_10gbaser_inst_tx_serial_data(1 downto 1);

end architecture rtl; -- of phy_10gbaser
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2018 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_xcvr_10gbaser" version="16.1" >
-- Retrieval info: 	<generic name="device_family" value="Stratix V" />
-- Retrieval info: 	<generic name="num_channels" value="4" />
-- Retrieval info: 	<generic name="operation_mode" value="duplex" />
-- Retrieval info: 	<generic name="external_pma_ctrl_config" value="0" />
-- Retrieval info: 	<generic name="control_pin_out" value="1" />
-- Retrieval info: 	<generic name="recovered_clk_out" value="0" />
-- Retrieval info: 	<generic name="pll_locked_out" value="0" />
-- Retrieval info: 	<generic name="gui_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="ref_clk_freq" value="322.265625 MHz" />
-- Retrieval info: 	<generic name="pma_mode" value="40" />
-- Retrieval info: 	<generic name="starting_channel_number" value="0" />
-- Retrieval info: 	<generic name="sys_clk_in_hz" value="150000000" />
-- Retrieval info: 	<generic name="rx_use_coreclk" value="0" />
-- Retrieval info: 	<generic name="gui_embedded_reset" value="1" />
-- Retrieval info: 	<generic name="latadj" value="0" />
-- Retrieval info: 	<generic name="high_precision_latadj" value="1" />
-- Retrieval info: 	<generic name="tx_termination" value="OCT_100_OHMS" />
-- Retrieval info: 	<generic name="tx_vod_selection" value="7" />
-- Retrieval info: 	<generic name="tx_preemp_pretap" value="0" />
-- Retrieval info: 	<generic name="tx_preemp_pretap_inv" value="0" />
-- Retrieval info: 	<generic name="tx_preemp_tap_1" value="15" />
-- Retrieval info: 	<generic name="tx_preemp_tap_2" value="0" />
-- Retrieval info: 	<generic name="tx_preemp_tap_2_inv" value="0" />
-- Retrieval info: 	<generic name="rx_common_mode" value="0.82v" />
-- Retrieval info: 	<generic name="rx_termination" value="OCT_100_OHMS" />
-- Retrieval info: 	<generic name="rx_eq_dc_gain" value="0" />
-- Retrieval info: 	<generic name="rx_eq_ctrl" value="0" />
-- Retrieval info: 	<generic name="mgmt_clk_in_hz" value="150000000" />
-- Retrieval info: </instance>
-- IPFS_FILES : phy_10gbaser.vho
-- RELATED_FILES: phy_10gbaser.vhd, altera_xcvr_functions.sv, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_10gbaser_phy_clock_crosser.v, altera_10gbaser_phy_pipeline_stage.sv, altera_10gbaser_phy_pipeline_base.v, altera_std_synchronizer_nocut.v, csr_pcs10gbaser_h.sv, csr_pcs10gbaser.sv, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, sv_hssi_10g_rx_pcs_rbc.sv, sv_hssi_10g_tx_pcs_rbc.sv, sv_hssi_8g_rx_pcs_rbc.sv, sv_hssi_8g_tx_pcs_rbc.sv, sv_hssi_8g_pcs_aggregate_rbc.sv, sv_hssi_common_pcs_pma_interface_rbc.sv, sv_hssi_common_pld_pcs_interface_rbc.sv, sv_hssi_pipe_gen1_2_rbc.sv, sv_hssi_pipe_gen3_rbc.sv, sv_hssi_rx_pcs_pma_interface_rbc.sv, sv_hssi_rx_pld_pcs_interface_rbc.sv, sv_hssi_tx_pcs_pma_interface_rbc.sv, sv_hssi_tx_pld_pcs_interface_rbc.sv, sv_xcvr_10gbaser_nr.sv, sv_xcvr_10gbaser_native.sv, altera_xcvr_10gbaser.sv, altera_xcvr_reset_control.sv, alt_xcvr_reset_counter.sv, alt_xcvr_arbiter.sv, alt_xcvr_m2s.sv
