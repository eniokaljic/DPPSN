// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h66agBFVuDjQfqH+Yc47ZdK0ZtRvyU6pcVqggbj95FN60xlhRtDAwVue0ymApwBO
rX3xR1Ghraa8v6Mu9GaeIflPv7AQta8GgYT9BK5bgGD8BqevFPJMcNKuNa0Qvwkt
0Wsha9xglnNwQbkqyergMCA5eXYaOlqiktm+Wy0DroE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10256)
r08mrmBzO6vNAYlPbpSZZmefkYBPzVx2vOm3pi7Aqon6iqrFxj37J9i48nyW1nob
pagowzHtI+VrjsoIUPkleUfpH9epXcwTimTIYUjkjALR0PHrDjIJXo5ElaYQ3PpF
exMjJK0wQZFhQKEwvuDfC0h7/UEZu2zK5ThHs2lWC3VZMJ5KG/BcS1P6caLPRBxs
B5yyd4MStLznNN66RlfxIk0GMOTBoD98ZnKtmDMwMHR+hmjr6o/uHs+27Bt0nU6r
gh1Pfb/6WvpYmjQ1g/ybmCQkWiMjeJpYih1R3FE+FNK0S4LFGRxtESUQGrz0cgAd
7p+nMQP+uvnHIHz6i05uvVpmJj+L02RmLheszeldRaV1RM9YH5q+En9JllHE7t7u
U1BUMrWxDOfSjDqDG+jvtoevZJxP83RZa9s2PH5yFg0yLvPD2MaOtKykHnDNCjZC
csECC8FxPcTKK9xGUYFpMsMQ+4HMvj2VUC5ysdKPUZUTRuS6P9LTnyBwQABcoVMw
URiDHoDWQLuox3Etd6g9Xa1FuWCYFkJaFjObTitK+tyr+zgwLqNAK6Zs9X3ubuBP
9NIbMjt8wtm3KSY4H9RdE1qooiRcmvd5xEFt16ceXLZm/Toz5vDkg/zaBrjy2E20
jSeykJVlCJMdGv3MApqvm3+BLkVDbp2Vz2GcuXCLh1k0vE+28o3s5MkVQPF7rjGs
6IKZuRYHzStqwpyCfWVnGtIP1YrA0AB7y/+X248kYhxz6q4l/5GMYuh0ggbVwFDb
U2QEVvSIIl363jLMJgQN+rxKF/C0nxHWIY9v/jh7Tj0uQ0UG60eySH51dPIbtiF4
LFFXl7q3LIqeMOvfi4OVW1Tj5AwZ6XJuudph8Wi93VIzv5FBU3lWHjmCBfQY9/NA
d7NKVV501qTHPX/NAz94IbjYnyRFirU7RAWnnHmHg3ZifDp/LtE6dolPsrOFedyS
J2kIlSMFm6qhrocDLJDCO1j48WDIu7Q3OVtmxnVBep5lF81w/a9h9ZpwaRz58bBl
95fH27au6qpMcUUbDSg48b82o/M45dBjVSsq32PWSmaQD8bMKLsP09UFGvzy46LW
uC7NyCzRjpFYqmAyidmHOlPpPg5NHveI8/BlVpXqxa/dPZ6MyAEKIPPVmQHbEcN8
m5QKBgxhzmfvMK4iGkgtQObpVGmmKZqrR4ZE31miZ2nZb/RSuBcOCvwou4NEHx++
Gy8iiwd22l7FfG8vbM9M040rZmFvq63gokbOVNA7lKhRlTJOH0hW81FreymYhKvM
SrkJAcSCY6iVdaGJ7G6bibtfvz3FD5Jp68ZSQGy1+/dpbT0saRkbs/kWwFJbX3a2
zCQjSOqfzUPPZXEKUlLiKT31yQFint3MiJK0uFTKXaRJjr1P4r+E/FdJSZ9D8bT6
rhKNGpg69cpKNasBmD0U+MyCexPd5gXdSnz8HRLkK6D9bbD7z5GDMcJ2WIwSHR56
/gmKhKsVQwoahmZkwPPbYqYfEutuaVIx/8JIg6dBXbPn527UApg/Set4dJMq/iFg
9vkI3P2N/sh9Q10ZIkl11Bk3wi9MnUVMoVc+iw9DzRK8DubXu6UK4jstJRPVSkRp
s0UNQW5fTe6WBGeGMYqZma/x1MtEAYMkA/4qs8TwMtFAXtHqHHhne11bmie+QyJj
1EroHxJmKgjMjs6YRBoSFnq7BecUvBYlIhXkfJXIHhkGSBpSCYCSbpsdB9Rwy4Uf
51wd3Z2z57eFEHbi3ccM5PAIlc03sGXH5ueI7jUGFElww/U3ki93AEIBTlSQ+kH9
hODtprfqjVGb5munFzRIMYKxDZOIDQBN9bTrAU5kRfN5AhQBBvOFQlxMbF1sKoNj
i9qvJu3B5/dugmMVKMqWNXT8GII2g8OCRXiHH877LjkkDANc5fFuOvAqyFBHoz1a
NY+341abAMU/79oZ0IIrKRfT53wIKSh7AFqaPKODdMiYPSGuULZSabdxt3GImlgY
LcFLFQA0Ayf5/YKz6sGpKLbU9pGhxp0EI1lYT859GbF5bDacaWtQopkHcUw/6ahp
DpTQ9us1fIo+59HtFQdOf8AToCb/zZsMCkRO84FnFNlZ5iMmnUtf/gYJ1+Ur1Iif
DAx4Xey5Ue7qaVo9t4ML8pNUwgDOjNXzIBLjZZtNjg2jj1zU2bjo7wj7HztdZnkQ
ac53tA7dch+SfDOvR1M4TmRDNiKQDrWSjGPun5ibAiCfUgFnR/j7E+a4MBAGQBbH
O615Xri/SxZjo1cQUT1LuwE8AHdMuzG6UNf1Y77mNnbaqvyEdzsYuCJPkYfh25wK
j8WFJRxbYTm/Vjl6jhFpCL0kykFt9DosVotw+opxEmAH+ZnbYOyQJSV8iuf8GIhW
JdhR+EOuSZOMv2TEAxiyxBwRubE9VhqjCoqYHsyu3QhDunhwGsDCBoT+5t3gtuJB
LxNDWSUVaHLAhWhN7QuVTFWeWfhb2I3ppUWL2DwC1GGSyesU0qS4IDsqMHgPiTpN
zETPX2XaF9A5tu1wD8rPhZZtD0sYT4WqBp/zM/nYUjM0I7ZSERLnzjuFp6BYn0Mr
fN9/WFcKDHeV77Ti6ZfgBd3AsfjEXTjR6MGjcVkbkl0lfzpc9z31gyModcxqz/ll
iZw3BnObm3D+OaDc7rMGC54Ggh5kTaqox3JHkhXbJbExg1mpmqRQq3+nCqKYqZHI
0f7GRrskimVM8zL2R8TE4l3ZUkdIPsPxw3tcYVooVOiIeL1lo3hn0MPY1/XDpjoV
FlNMSRp2p6S6uIzSLeYpw7eBW+4fCeDSGsqOd1BiIm+266vK058V0ApZwcwbCyr8
i7436GrChyg9rAZQAqNVJJqw/aWUveK3mmmceeBlCjkvk5PfQUmQ292oM0+Mss2q
BziMf79Af/XF7X6d8IiIOzuPP98aLqHZ+jMnzl/ayqg0wuoFZ7In0MqAyIpYjQv8
jo6F5nSb6gpkxLp4VgwQ07WmEEOb8QIkLAmnopoW04E3FazO0nzOZgJnLZlJViqO
HT7P+dRckRbkQ2lvzX7ByHNWCvFXLIN0MtCQLdlK2d0bcR98G2kYWijKuIYNahf8
G/FJ5620LhBRr7F/wbYwK6PE08Bz9EHMr0JzAClRBulWNLdE6j1u6x3WTHGTI072
PpEui5H6bSaPve373SxfZvlIeXzAQ9k0m1adRjCopnIOxchzoylndMDWHdJHnl4L
yttsT7igwfNGhw8Bv7RB3TxWGK33FRymz1ZpbbNnMC5lBgUs5mq/IeH2Zz4L74/9
khkUKXDJ3rJo6nRL4rzcVgJhlbVw3N3oKoINxNjzqBTFG6pqbTVM543U8pZ75vER
1qmnm2FTDfn8kF2gEoyqFewEuCSiT6ar/WoW1px+UT4r46mnwpQXrsKg97Ut0kqQ
7jBeAWXKbCoyMN7eu4PIXVw8E80gAz1kPEsCwlNI8i0/Y94XrwY1ubgZa3/CJXtb
c1SxaNmcZ494u/Vo6ZEKAZ8NFc+cCZlEqOqrrLH0gEaCyQhYL1yti6KzeEF5fb9O
X/IJAr2np1MrZjoe0jqhgIxV8+RtKuKRQ/NMXVcwHlho9WxvmkdZSMXlo1/sSHcE
XGA4PQJwRRI7KAv+pfCWojLd+eT0xUzhf4D+QJ+oaySvmWR4S9EBxk6FIV5fmJr7
wzDGTBuUXdtfqtDesWytfXDcs9ByEwJhDHqG/9ffzjerj3H5fi3CE9OccIWDaiC/
uo6MghchiNxc71GfMRxXzIi6kTyn8fBQ68fYrbttfss+gLehQXoPqH3XUhbOVIC5
0OY57Z4+KlTJBqlKhsd9OiSV6NF5tutlyeqYkRvODUqnUAE2KVKCnB97oMOfB7Cy
DcU3RIkb91yB7eXZ8wc2HH3dnCNkECr7bjpflZlo896mZ/EmUyfxMrQKEZchwl3E
eWDR30Yb5BxZkhD7nmnnwNP59gYOxK34WfhWVY3FwGSzDxZLTMj+MEvfUPxekj9T
ZZVfI1A3Z9HfAYNjxxVXE1F4PtVFswjmytQJ/AvRcBvw8LjKjBoZE699qilm1NXj
EaJ8dYdT8umr83UutASalAo6iwP2JFGGYUHYrvb+muSb6moq+0w2hpm90vQKEx97
f4GMn1eaASh8L5Xn6+LcikbUHkrXM8keHnspkEj1+eVlHLZVS+iIeS7Z1ltwiEId
T2vFnlHoFAbG29fRmfFrZ+/qu3+CW08JMv7J9AFVpr8QbglRsZXxuxPzaLl6vP0g
YKwOpPHupoUtsVW7YUOmW4Hmxz00MVvcNv53MHXlxkDMqk7cv3rzl7awnhKLZ0G8
7Aslj/5olQbzI0ISO6yD13SZZGuwyExbiUkX1WFlEvvr3der3y3+3OSw+XmWn2ei
g/BlvbVey6YSwobek+hZh5g3XkhH/oWmcsBAtCJK1cK4AU0NuJSO3HQdk4tB7bUT
krwArmrqf9jCyEOH6tcRSP0nLp/R3vxbU5oHNCxXqmfOyJFQqknWq8o4m3wkTNum
/IxpvyeDbblzXIlQP+kAbBKmgm+vKzbFq4hFOpdS6Hsm1pRncGNA25lghdxjsUGs
js1QB20wDw8zyjX/BznZNfs1Uap2JgmwU+GoMs54iccfnBxDFjzCgU2GGPsv1IDs
uJvrzzuf2Ti5QqNNNeLxP/b8KIJE6FjsQhbIiRWzF3Gysy4eR9P6EzHVkt1ZDrTM
hZnIhE9zga3TAG9ckaUJi3RF/pnM05Z03TNk72zXaZ+mJ6r3ywEsNaSc6PO0qSEW
q5mz/haqGmlCxdOdN4uJm6y9CR+1FbI7t9/bJvjmZfZjD1RHDoL2fEk1Tm/xgg/o
lSUI7QbaNfmWpAx6TxmzSnyCqmJzbMzWVZJmQ7Fh9fikLtzbTm5+uarI8d/pU2ZP
O0ZYkioaKH4hwpfQU8aXK0y9tmHzx0NvRtD8YJOSdvpfYjsIEL9kq2QOmZ0rfje4
Wdh94LJFiA8IVmp+OQIKQ+p88OFS5hFLDIK4zhk3bS88+H+DE31SXEFdy6MmIgIf
mBBpcR+4iqjfnffaXpmuGIhgdIaycDsXTnDdJMbjuoRjDNVhWzsBE3YhkjqupgPQ
yRuyRfAWpTeNmaQ/n28dVj8/G3UsIFyU8VEQ5vC2G9xcE26n5/8R9crdF0VGrNn/
lX8ukC5+t0hCQXnbp0/PQz5nHCLJd7ekISNVSyS56YHiyvrGC7kBtTnSiSpNprLe
niR61hdyTsDlvuMlx7kkZoRaIGC90+Bmj1csPQUCxzkwk3zxpxFEL9Yuvw3CeJdM
nALejfsd/GGATeJ0/xp8WLzH58/9y9NtKVbG3t9z0NkB+/Mkemy1qHgMzkwelyxH
F22BXDpLZQrEyanuBHuaGy60c7YOVO3QbSaM1JOnBGiUMNsDNIvXwER6S4MqZ/d0
Lhe/WOKczLjxhKgCgp6RD9GqpN1Kehm8+9BoiB47xhzc3ZARcMm87J+vo0CKd1cu
o/y200qzm/PeAv1i+4juAbQYpcfxT4BXYoY+zIQd88fa2BnAFOLsgG3iGqS82b8G
fSjhOMxSk10OEDFuB5Ndk5f0zBXw/kynsTHODvNDMVGk2aGCdnSQHWOUhku3JwZ5
fr+PCVVb2FBkM30LchZboqXsUaicHib1pUSzEufruf+s9XDxTQYeXwIzeJDpVsZ4
bNOVhudSR95pgolc+jFP5agQfrPuwYlALDE2CtMoKbqqgN5vMpQ7mrKnVCmPSHSN
oAKeOu3iFO8rtq4w2Ho2jInHNlSWP9AeZ7fiHS5jOZhd86TajComh5mlQuWieRI7
hwL6bN+BamSWNG0c7DPxrqLDFzwXgYru99wkYaUuYEitId7CLNdsEERsKCK2hBDA
XAiWSuf50CX132ZXcTQYQNq6uvWR5No/9ecwMuV6L3Mf8yvL/5uWGwz5fdgUbmA9
y+XArPhQ6ml5qo4Dh9gEJ2xE0YtLum4zbOHaLjlhNWQt2qvuSW530zj5qadHvb+E
0PAyMcat3+S9RjJVb4SGpqwdzxhTpXOVBRF0g+HKAwWXfKexyBtvc7X0C0H2PdNc
k7c/P9zljNM8gA6wokqY4pp/Cq67+Fi3Y+TvgtlOFbsMfZfmtqCxd2l2P61F+Cz8
T0LhYBE+g1dm9df6+D6c+Ml0/Z4V53lU/6VK9gJOSSFw1AvZ64ZexjIM/naM4nN7
xR3XZECGKEIQ1O8re9CWBjQysUv0IiGLuoSDsYn28/vyLSUcpSEY4DSukS+Kda/6
FMli6kqCvQ6gfqIbF4WPVz6Sw5V29LarFPyinoLTglKCTfBFn+i38InrFnoQ9/9j
fir8fcj4/l0KfcSkJa98A+7cggYy/u+Fagzhe1jL7H28qPUcLj/8Rqc1VlOqb2fE
Xc5ZATJ8H2xAXIOJIq0PTNxkHgs2ZpSC1euSmTo6/fkrVGZdgq7fRJzHSqkAulQQ
6ze082G09c3yIv/KP5qN0KqY9z9KM5tdgKYiBqVYHmQQcXZRr5QhvwnrvHHjasxU
jgoQsjS/1NDEEhY/Pl9IvivzxxVUCzFnp8EYX+f7PWcWBv6VwEnCF30SUsq1OKbI
VsZ3kvqi6KTLke3/OQr5Qqy8oUO3jTegK5Ax3PfoaCju2a3+roRPVjR+Bl8bKd33
b3zhUqJ77RUxzW5QU2PNlg2F9wIuR0UBSqA0qVDwDC09SnFetq+hmi97fxinlVVi
O3R5euSqKLSIHOCuC4V3fBaCJE1VyTzuZDHsm8xPF2huVVBUvauRctLWO9zZMg+Q
x2prKxw0AnYyqFVuxNFlk9YjECzoLyig4ZkHl5Si0C3+WlGuXOpePXpWc82lsk8e
an9qHfTZ8Wp8+vx8J1JjxIPBbBe+Ak+B4kW4hU9n7CmRjCx+bYLNLyTnUXWE2f6b
rkLhstQG/tblk/voiDvvEvu+MRNnjrmbSWBe7Si6bDCXdzZaHDpnD+Y/XmEZQ82V
wwFdp81srjZglAUgnspC/oa4rymxyQai6LtLEZ6i4Jz6IaIWSfFx8mlTv98ahBjr
7dMnp1KIZAlEPlnqrzN5ATuXmoak579GQ2dVIDh0dIU3REM+lEMvRy6WXKVTOcYf
dDnpzyGyGoZmbVmN4KWatwK0SG1gTRpdc7CCl4vuUXr6HptXXGkZso3Nn1rznJ0A
mlc55XGv6W7aB7TmsGLE45LnVBeLyjQjNDDlqMVaYnr/Rmtv8qDd/JCc48gLmfoF
lP6AtCcbmFSuKEmJGYFdVIyPknwTHlIqhJY6BB3tvEFIOZ62/Sg5aaWzKW2B7wr6
D3O3HI2+j4dRWwjzP/xCPFReHVOopbMfSUkZVHz6E5sr9yNbvaQ/gNUigAsIMbPR
bzJDVjt2NjOmhh3xTlGRtP8sgdy8t+myWEgFaUVZgiQkzjJtuLYOCKAH17/ywTP6
WNJ0zp2V4te4P6Ky3mxnuyuW7gW8p/VXtm7FaUFEuleYswTiO+78/Gm9fwHHaxHI
swLlr3rV+nc7O7y9kfJNHCnpcg7lHm1vp4zbZuIMi8YwKOtlXTswq4sopvUDtNyB
EPN2MJ1T6WHHn2qOq7xAu2fhdpLeiW5OlV/zh7nApCD6rmKSdQc0o2fuzFeUnF+w
4IrYdrARhiNxsjeXR3jChH1PTtc9Jc/mSqCIieeavgy0iTEkSYRKpEekykNzmEDc
WZWacPe0eS5VrRMJ+ZwPJ5pmOuZB2wWnJXt8HpdumR383OSP2R9bhkuQNdofnZSf
9ai9NnO/ZGQ5501hFnPrNGCo6F80Cqe89LN9fWtLiFNg6M8OOTQH7CTPhDiu4l9u
6fdN+VHEgQNqtI+Qo3bPtEVykPccmkN15GYXpza3TAPwlLNLAfJKabhj5fZculRw
AREfQ0k6HibhJ+LuMSRoZ93A5MkmqYwCn02lZMlDNmuVhubPm5ytJC6cQLhQ/tyO
EFRCLBpeYIf9PNWBURXlR0fpAu2LVDKhV/yGOD95yp+TmxqCBnAPOC9adPOsXkZr
GZeV2E5MJbFOLMuMgLB+Rd19lFBFaEyIxiVYU6zoK+ulu4hje4LQyQTazfVCJLdc
MHTDBjQNInz5QK7Kpr2WVDK30JzIYLvo5qrSQfD57ZoPdRgaI60VEt0AwoQuIST0
FJYGKJu7Flys9PiRUZdAZ8ViRbYw48ADgYbB1P+C8x+WI9c65eHxEUkBVfjm9Eo/
gS33f5WX4yttX6kPwxS6EFTsjrCxdj1ZBo0bJisBjbiLGGlWLDfrSZLIe3w8/cLn
lcwjpqcjwheRQa54UFSew24KyI98V0ElTAbNU+hZE3Fp2bOs6aP+tkZqmj64qKMF
beK4DpEcSnl6mPzGKkFNL6UERoMNrj0D5hvw2GnvoO7eiz2ZIZc8+UtsIFH+E6oz
6ggdLLzfUxyURmBMlJBLb7f4Y6JpxIwvwVW1zLPSrhInrjDDBCy7gcA4VUggsdPq
2aW7G1FNXEeA5+Ov1sATniOTsd/PYYeHz9l2EgklFwvBF4mXKcU4NERtPP2mKOqj
vrVTKc8QdSdNelQQfP8rKmNwmvqypAnydP+zyhzBM5RsTA/ZKt5sCgGg7x3AEXAj
Vs0xBmYZg/xoyGN9FIaNiBAnpXVyUHYG0sDSTX2QC8fFsbp4xCDgqasnik2Aw2d4
sfHK7wzbK4ZKl0EzHOeAeNdGBCQ+ECyQlbD0OXaM3g8gOmPHFQLojBMe9ydfnRhp
W8jvhTUpOmgbcgW6n7QXUM3OKZtfvJh/Rs8dIHAyeP2rFJwGT0W2lBPH/iDKhvJj
KzwJmwMu6X2uAaVa1lhAuNuEWvpgcYZI+PuAKnxZQD2JcLuvRLJhZSwiEZZNFeim
biC6oglCzm8LcJ9emTVvVzQ0p6CcG+TM3TsDH2zSY7vPs3AziMAFRcjCjUlA3Oaf
okq0ZgfgQSkbmTlQsz2xnUYVaWzqqCbG+zV/XU5e9pxCWVhZnMgJpU+MYTHseeFe
Q4Xu265utpRM0Uw3Il1nGAvxSERqvYacoWgSSTX9gVQaixig/FlgsaYufQKT7OmA
kg7lgwnXuerfaSa0K/oektnFkLBDksAptdmnBVLr23s2TO4oQ0U54XE+knxHEG8T
tZBJ4rl6x8PcCIlDVfw7tRtEYT/v5GlHMlZPCgluAc5FPF/sWl/PS1X19PsCRZHx
AC5d6Au78lqO44X/cUjvY58wOZ5dV3SnDtOaeUrnqL9mkh1gyj6oD1v/rxJMTEYH
GFsfU5kZnHhtRrLMyTPxBOhwqYBbR7oseFJiyd2O74Pi878n7uLeIuaVsTtUFGhP
v7wvA1wN2dTgSCd8V5faDqvO0fa7Do7MgOAS4jdJw5R9zPCjnYr+CD4fb0CpKSdi
43CrgX9ne5YK385PyQfWhOMCFXuNi6HOZvqRDE30sOyX/tGxJB5O+JYbF817I4dX
v/fOTl6aieJM+n1GVLsG7Ideg+OqyjcLoB+W5gREyQGAD20axJKClsEuQJO7LAoQ
hRHtmFs6N3Go0z20Nlcl/u4gOvD653Fgg1j/dGZOxF1mEkBS573gM0vP8c+TVQ92
GeezJNBVCvc8b0BSu3/mMhSrPwSj+D9Y9JqI671rpCm+Fuv4a6WiHvKiNUN2gvNg
2Wguw+XvmbZhseRDPgleg/BGiR6YsGCDs5bJLCH/GmK50edsUtS3BKQO3k0SPm7W
1NFcvyY14ezDkQnFWnTYuGYzhSh7qBm6hq3wBp/4Lcl/Pjtw6iy4A+bSlluhIEML
HhCGOsTAIDz1PBoD8o4opq/iyRpPQx+EBCEvGeLtGCY6F/m77NIba0WXHRJp1Dko
KTr4a/EoH985IUuHl7w6x4jEVyF4GAUWEWr1eJvppE2AR7WaVAsG6ozlzk27dlcb
F3bzakJChDtnKxNINxWCWZzI8++BpHRipYXWDEtedQLNRAniWi7+GpR1p9ZCPZG+
qQtkgftDmDqtCsj9S9qx3b23BgQtmxGN3UmLhidjg+ve36ghZQyN6iJi9AmGl5Cc
q/zd1aN3e3aHAVlkgAUQcSCblhEWxUJCQOIsUezT4EdCgvrOVWRsg7K2JFFT9PzZ
5Q2QAn3L+YjKIY/UX8JV60OhXJoJrvMcK8IA3v6enlp5LqGsN+V9b54NlPYlvS6q
B4u3XGPiW3sm74m9yEzELH5UIqcOBuBeNUQRzjAHY4h+CO77yA4syzPTw7yJ0qtS
ZtTezo4rqDdPNSlCCMYSEgPPJm8RFSMKqSfWEgVK/vfR6ngRaqrKhVwXxHbVDALs
oTW9p0IT4m2Zvjg6zKm0gKkhISYpqPOo1eTPW1hqE86OUoO87DV92G2Ublmqjm8U
Sdi8kpBvnnh76vjc3d8LCLcOxeZ8OudDK/dwIf8+8XwqzbMHgvjGRmrkTqLvCZcZ
aCJaAllutuQDO+/zcWe7YWrD7AtoeokKawQ9RLGD2R6smHXcIXGCW5MoJzcyMcwz
Lm2u4qSriP7n8WcqVZONX148dAzkUP8wF4rze5CjVkXYT5tCTM5JXmQppDUjda5g
SwA3Bz3Q5DehGK7ke54lYcgUCLZSha9kQBC0+1SMuTyFv3e41ydMRDj8fJidcC7t
9euIIH0Z1ATpCRVlN9Mlop7VPqNkhv6uqoQYydGvwfT2Ih4tCc8EIKxlMuFH53zP
po9yUBF5YXMgl4EWYyj+xoC+tFN+kFMo5YJ1G4jYQlOHDpUdgRHUuFoBg8Zlf9kj
3iBcs2i0EfkBOXhlDTlMxu2XrvTQWd/6QUbyw10acdalJh193hdzxA/y1iPXmGvp
SlytJcknlh2YRJE7oE19of7+4+ADwqVKw8GTLbiASeGFy690rL+lCOTqnrSL/edY
KfrWiPcG00cDBfJrO1Y6doHrjjqNJZEQf3ANRikdAPxvMvUdkuIeNcXgDWPVlZ9/
c210xqOivWQskf26UsrgiNCv+J5gxAQ0ue240Tupi2Qa+A9eJBSUqClywDaPU+hd
aGyCdQnM/fDHhEAZxLUJZwgX50ci9DM2xDKrhJmfQpTEzFoiy6oGxIN+ZbA9ceSF
N2qSDrnoQAo5Xv4jH0GTdjE+glB2LsPqlW+6/lBwUWs5y9l8Q1LNLCf3A+sv6oc3
DP4BoLy5jmckecS4x3lrD+crvqrXS/C8DjWLzaDZ9tfEi0SsbE1/Tg6bjjaPT6tK
NuEC9N2RsPAyZH3noOASAFQfPRzb2/T1zvGC35TWLc67WklMxwgjgz9fr9bQs0Fj
i4ND1D3bePlzCpuYr9IMnkvOGR6CS5gTXjfNZKiyoz/N8UrOzvPDrMYdeckOoBgM
+nFLJfLpjG/sKeSy/depKWJ4Pas9U8kvpRoIA40/wvWX6Cak3Pe0zi1dOkkiSBhB
tVppnL4NhDnhV9kuQF0DYZoVRveqJkFw3VYcthZV/HZ1PbYKvee1WLMQV7ZXCsNw
ibOF3D3RlkMGEO9siKZ1X+oW0YR5mr623qEn12/8JPGRq6C+2X9lcT3nabmo2XlK
x/kOVfQgt4EjPFqaMJZ4cLUHmELd2FnnFz717EgJnSXYysB1oqqb+VRqjkZH8SAf
DyHx0MfI8C5iKjeBTxAX295UkozHCY/Cvmv8C7uqDj1pzJBgJMagmVpCfiM7mB3r
FsTtaYjmVZ4CcR+D2wREpZnLReSc31DYSSvmGIEkNGsVCOKM7C8m7j/X8G/MVymS
h/2mBU7wE27pZNDdyBhEFtZEJy9RHTB12rbZCQS+HUx7fYV0hasKdLPb6xORbsye
k6jBaX1Z/h/ZYbiHZ4EvdtyJ/URqV7hhmJmLJdYTCss9K5b+ea3f26xBGVEg+S7p
215nkjlAJ3FDCMwV3+LsWk3oK2+Rt2DiGJiOhXX3zbVx+4viuh3z2qTAqeAqLr2z
RK15XBhM/htcA3U+KM1u38Zadk/rhJQ9xkJQBAE8iKK27nvdMfi/mU3xBmLAq0PD
qZmAab5HKuMHtLZkfRwYh/lLhwPmOiSQfl5qIB0e55Fu7YoOlcOZl//gZDt8CKX4
fq0Nzm/j5fZH2ncdDIhzXGqse/F3MCjgzNfUYxVNxgE5i2yG5lYdXbikizyuY0Dt
slNXjd44rX8qGj0Z5l6zwS8hxoQVypoLI1ZQZetnzgWOd+Whfw8loNlX6Q18Fi4G
x4d631Eu7Q3x36oiNwHaie9kDuX7LofRAZfLoTF523op89hkncpdBYjBuWCjyFGu
hg8e1IvCmRE800sz73+14TMA6h1RAn6vs5lGZUtlXX1kFwZJlqL6qN+ZgvlXKHcn
wnaTeyc8D00u+zYqGyXiBm6DTcci9KEUn3/0a+ZodAmsFu7kEZLrzBqGS9yTLDim
naie4cA8xh26TllJDILh6skOK1hkwAjWMoVITVDMRc96iqfO2J8StIep4jCilMpE
Re7vrjVNsfP6MtnD4WFOG+BOtEAvKGjGgnxG97RV0Gtqk+NhZOdZ1M2FN5nx8JM6
0DyNZ9xtZP81osA4MZwf4fwhMzyVfBY41uBjN705JLLfeREVCm9HSQnoJnEivGhE
Zdfizvvc6OXwjriFyblSuzXoJmX8kgkBqtcL/HtAbxy/4cGx6tQ6fbVv2/J+SjdJ
AHW3j3G5PHrU4JySZfCNfcPloc8xu2Bn4ebpmxEbChVpCmeRFcjJl3cGG2PPsP2D
Ajs4O8ooWKR2oW8UsKCwHsEXbH5JLkb2hC3rgu5NTy45EOtrYaSt5PyMKnhYhu39
32bEb72S7/wNrt/nFEkG5oWcMadplFXAxLJgbiRFGU0goMX697BXkKqPkm0M/kFp
9CjR9GeNW6UjJlwAWqrwP4VGq9GxkJ8oesPER2r4K3wZSPg9qWxAQB3fBDgTEOTx
ZNXvEI6Gl5kRljEKvljOqTU4vw55hwH9wNJodtk6yXS5ViCBRJFoU9boSXGUIuoh
W4NPxV4Enx44eFlweMI2eKeeuZYcAi0TdtoZ5KoyGpPincFDQ0Vedlc4nnRJFcCM
KTxJ5TB9OM17DvCPYJsBN769g9Jig8tveOlkwAYrkHJRm/yVFFqZag3MqzumHvmP
l1lS9j1Sdajuftgt9CSEphruLsmXbR/YtstLJcrd+zfSeDmwzDUk5g7S7eSPZrcd
G86NKIxh6Gm8VNnXpljcm56b+O2M7wWITrRluKAqlLt29W/18u3b+7EBH+RdwNVz
Oq01ibawRqo5Lcx7L+qOec8eAp5h9TSRYNJDrAlGEAbGOsEIRSjG/90ycyyl3NOv
0cnkzHXNQlS8xhdiiqMnbhaDQWa/R25I1EHJBQGAP1pfGQyobGjbZXMPcTpuY+vA
HRTCJjCRs70Jopjh7+i0iCmeVQ2p8hLMdD+1xMmKH8r4nLMoHt+oDPGXf0H9DRxU
Sw5TdwS//g0rqxjwvDGQRRsslIWBuoOqZcxdtCACkEnsO+n+sfD6f8vOv5i41L0e
3ab/De/DbgSmnN/5sfejW7CsYSF8vOwN/J2RWmg9Qtx22evLcn9VT5snd3i7WqVV
OblDCUQD8aLTQFdh0S0TZj12FRt0WCxVsxnwSSxmtAcSHr1jM5FMkGkpKJxDMSNF
Z4kj+KRYjpG7SibmU0k4XjL1p8rfaYsm8KUP5XZXoh9Vu71flg8iG2hdPJc7dUOm
Fr1SgQI5LzMLh9/dt/cuqB6rRk/PUMgPgbe2XzyIIa+tpOgN5dQNE03FaNJpHHzG
X+FAumbDkeSF59sLYuzoqS5ekjx25/vtzGqHXo4nzqWFs0mpz0QK1OoffV3bH+3M
AoFCKaHv5vnfpWYZ0UMrY0+2fTcDJK2PBchYGCnB8Mo=
`pragma protect end_protected
