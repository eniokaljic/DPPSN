// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:50:45 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b12w8dTGHyR/RlK/1MSDTOey1CJG2/JIiyzH2M36EU8T2IsV/NOYhfvBp/jinrrp
BqPYyveNN1WKKh7rAZhtp/Xu9YaROKJE9E9AHcat++rMNEXLsMQPw/vIyTQDy5pA
T5CPg7p2f01JJI8V145J9xysY8i6nm7+RscIcaeunZI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21920)
dvovLQEJ3cRR+8XnP3KeMpycvor/o0DcGc+qLYTOn6N+dULupM9V7bpUEh9OlW1d
oHk6sNJw1OosG+0AJ4GFANNCpuQRS52ONKXkwm+uPGfdf+Y+dVr2oQkfbvQyOOtA
ORx1vTpSU/tKmLUnGQf7Gup0zlkj0cyLoZQFluifycVkuyWauXiMGqI500cpeUMw
VuAvu33Dbvi6takn+AZQxH9rvel8d71KcyxudzGYFvS/HgwZa8/6dlT5q2Or8oP4
Jp2tklMPM6r9O7y4mHWtY1+TVzOdfaixSI3VMDGbxrKAYNIGAuS+qNlFY8AECXar
LEEqmhT2eJNVUOgAiN1AxEuF21sQXa6vP7mj/8QpVt6hb6lOZqzoub9BBLi9cyBP
a9qOWai8CZNJAu1VpWBNoDMaKiu2bK7GCnSDGwtZcDz0nR2Dfx46oMHlYG89jJtZ
UxWtu/Si2tzWS+YS5k83t8EMFjrRYJn8tG5lCxBEFviN/xCYInazgmf1wD5GOgdT
gjj9iyLlYpk5nyN1J6Mf1PKPMswRMNWkOdo1aDTncX2tbg4oI1eOwGvX2ug0s4o2
jUE29NCF+QX/bbSWu739aNwtWDc3ZDIwGdxyHL9cyJoou4Em3AYHvDVnTLHR57Li
TRg3WwCBGpS5xZzUUxCpkWgSk4W3TafH8LiOLkcv9Fp0RgL//MNSFKWcT+wEEUG4
HlcH20ZF+JO1gp4GcsHdC8j62Z/iRUhi3jeccexdLak4SENirIYoPXDJIMvHMwqM
dfUtvDo9nmCTCG4Fw4DFzevD4AdPUq+qBSHQfPUhgM5sx2A2Q2aFgSqc23xzY03x
G56B55jOOb8p4XlGnD2W1sVMtn0By9vjIyvtes1PKkzI5wzv6bw7qprSWi8+uk09
OnH2Ap/lC/zmrKoYiX2gGDHUBvmhRb+c6tJFxbFWCFKX4JMOA7ay2cNc4w8SqCPI
XW194tdErdh3kDaPCRojUm+47Lw9j/fqJJiL7om2jV2tUQQZnfg5NdlUFyhabyIj
tavzSWaPQiiYCusTERSu4T0n6c2F2RqeDDfGB33nvFC5QjlKZNIGy3Bn504EJpxm
Z+5lG6GcJTxzvDTnxp0FgAdSpy7/bPHYQ0trmU2tP61DbhO/pwwH6YDK+lMDMess
vLoRtzAkjKYpLscvMJZiqgVvnO++eCAKV8n0N7c9CgR2Ky8eM03mj/c+vqg2dxjk
UJE0dlDm/wU5Ul+9xzey5uiIpZrWYv72+BWKVR1C6ZyrcxHWvHPCxg4naAbKgtn1
4zKYzBi9NCg4stY9N10EEW3+13HnwqK1J6+2esvzgf6GHZ3SRTXlMAECEa//btgD
Uaj4JCuX39Hh0hLYvdBNJ18B5ag52s7IHCC5cZKiLzhVxzyH31rYIgRfAUHKJ1Xe
iHQ/zNX7AgG1FMFsaB0pc43Brz+I7jLIu1mSOD7v4mYCa760GyhTWds8N+6nLEwC
nsOlC7U6Kp+rfrJO7+nKvmJJlKHV8KEJ5BnM+C+ZM03OZhi3DTV4pnif954z69YW
2See9U4N8WPM4iFh7G47xhLzJdR2db8PEfxwRgGTkjWeocmPvo22+LVRyk1iUBUD
GwUPjO0+UyoMpIEACSj+0Tj+hvfCDDjLso0i4x9Lc15r9P2oSMgRza2Jaa6ap+fM
TJ8LFWqQUodGcvDUNziEDSEWUt9P/kJknSuBCb4KaXYHN9Ai964Fb84ANyg+h820
uQiQCWjEjh81l8zw3gv1WfG+GzXkjc0QvvXFFHCAHxLadYobxcsRv/F0gaF0kRJ9
VH3VW/sbthX6wI5OiBPt2amXb1Kpy4iZMV86sZFJWe4wxh3BwD2o4VD8XWW7h2SQ
Wt4X8kUwM3MEsFN293jLEiX9MJAxvkvMSzs/7f3/qz55QoQ3fr8jpm0O6xisZMD9
mJwVBUQWcOSEZZGdBSlHHQpA8/e3uhJL7V+KzsXoY7SKtlIr3p7wzgWp1A3UkDNL
KBXIGIlFMMtdP9yluR05SMeg4Wn+4pIEyLdHgaK0SIGZBnNSIr/R4PTBKucS31pc
6qGdQhlIJ9rMFFDDVqvHjB2CvcGUlE7OhKKcP1kwH9Ew38/aQluL7DkB87x34hLg
H5QXbxrVtRQ7Ch/N9M+VP3scneCWbLMnX8x8MpJSSt/3E2E002B3h9aYCqcXqzBy
O4Gfy3hRI8gOE83erhxnTjoekB8V2LwXZlBVMNsTidUAz4sLzWNI3dnjb6T7jrjD
OvrZLsB5C0Oqd5pLHmtv+8zZF+qON+VOMIqnwc88Vk3/TXeIH4XCTnYIkav4zSi+
pJk/TMlHlzVZyhrHUoUVS3AXqOnuvM2nGdOcfohqdfmCRTtulXJ069dMmHCrgdfY
Ge3G0qKQlrjrl4sdrD0v4Dg4dr/NxKOPgTPfgi/7O8VpT2ERdbQiXOZj3OJ1XyFS
kM2h1K/W/wrQxzccOe3IKxKwZzatzFX7KQpLd0ucVuJtE/8VWGkRFw+GRSBOiCxI
ZF5opupjjs+EsjYLrMN7PzBIfnC0dagaNM+C6vdbcm2j6Mp+M3Ivpu429zUTXAGW
HWNhuASdW5zhVqgyqGNNm2vA31K5DNb6udmXq6eqJkjlD4ZGZj5xw+nF+uJ4NPNe
3s9e/BPQ5GKuX2QpT6t+P1d8rkudTvognodEcR35yGlW8WqK6KGbZpDTQR7dShqI
ZnnPwzzIjXIQHoc5lmD05If4yrGnbvUrJLX1lM+utA8pIwSkla2Z1aXQDAhepoha
FMytr6OStjE3QwX+w8YcBN6IwivhwJvlILBeE5OnPbDK5bK+co4nwS8k59rzvTJD
nVxywDkxYR/ngz1MdZbrQo7a1jRj4dxhPxvVAEwHkYPlvkgpGCtAnZ+Z6L6Bu0rS
ghgZrMljF54Pv7WjEqAEXyyTdrZhsTxuNLJ7/c9Z33Fzbb6ublnOu+JBWzbT9iEA
8ijArTCY8A184s1tXdJMcA+0VtWDdQWsqM/scehtsRvpLAkGYPnW3RClQsDVI40G
JVc1PPTUVhu5YUeH0/puywacYTJe1e8oNHSBqlfr+N0sQelPdRK24xEtNeom1pwy
82225ZKTeWZFrBSpWHETWaBVdRqdn568vBEu/Y1dA8YeQ0AVa+qdOo5ahKDjYrFK
QDo++Zt7a2mef0T5SXx9qlivec4UDoSNaRfnYE0T5WIKtV4LQjMW08eW0AYzTcr1
yM3gtNOZFQy8HhQf05anKqS/PenhNVo2X0iUtxBX53Lyhcz3Hq0HioSVAKV5PpiL
YyZOYcu88l0UjfPp8qMPYz9CqSln0fTIrNE20y3KYiNMD+sEZzGOqnt1y39gGVpF
e004+GHxAUTqb8JicudY0wwSIh7HzaAVyWElFQyt5rM/yzTchKxVPOSInvLJj7Fp
15DzUa3wjBzeN+rnMuqQqspqxLejw/mGDIsktxxG9Ak3qssgEx6BjKnUU3f5wDGl
W81ql2BMwDmLvqeFZ1MA9V0KtkWe2rTHoGRgnEsSd/+SkSgohNEO+OPAf1uuRKm6
PmHY4jqMD6UmvQqoHKBEN/Xh/Ne/MV5WTkB0nwdqRevfnUmNghmmJpPoGRk0fp6m
/hmASh0qYJ+IxKRMpxhkkEJw4F71ZU6JoINEcTlJ+BnhvoJaIkj0VzKy/Ti9Olel
mMbGAGn0KG859lrq2ny1P1i/Z+T7e2GgudnGVpwfqWDyhWXfAWj4wbQN/xhuFHUA
jd64AGxzmooghZYh2pTaI83ru+Y3m1qLbwlZ6T9kmN+bQvciA/x0Xs1eV+oURYvp
XBe4jpnAdmzqwI3I6vSEUGgtx9SkT4ShgF7zwPSHSUcgT34eOMN2pv4OR3zVs5+i
sZ43Wtofrn299vgmAFGO7CcnR/MxqfE0eflLc19uWZv0CvmquprAPM/j3515oqT5
TmVQHlN0SUXsy8foi8yI8iqME/RoNFMwh9tsLrUM48OLoFn1oa7MvHoKUDkyVcgx
qaN5a0afLU6o0giT8sfSyiM+iAkcygfNP4UKcNNX9W5QjwLGu+Eik9Iw5yyRrzmf
1xXp27PdvD/SYaeog3Fy8ZrYLCeDjFCbHB9ukoB/OFjQQUWEeY6qPGIH0XHfzUlj
h7hCCcrMn4K6KhN4Ow7N56qytQTrP/kqWPGfxrFohYCkSaqsQ07iYPQB+pGDtQQt
bg1w14TB/txhjsz2zrjGcPIYKTFBb1OYz8JO3myIu5nl6QQTyV1GM+O8jDA7Fdvq
WMtM/EVmeKP9WdW6y+SuAK5Y7rJkH9FTFW2z461ZKjxLLuCC1AaBY1CkDId0hhTM
2YPiLiEifPLBuzgnYMMPm/VtXmANOmjp0fJj8Dq4tAzvTJCHRdJxb/oiypEnoeId
p/3pRtW52zwyGTj8fbKsvMgFsVSvvDYIhmKEHBgWqpyplsjAQ9mOCyUqGydcBRfR
Gk3EFGlrLXELc1/0fT8+f+lMqWHxz71d4lrERysTyYYlwRKy9y0zUiHim0TDRiTj
CYJlAswsV/T0wDxxZ9cDouaVvM9ce4aMpepR4B5babq+rzXAEprgbWcaiQ7skA7q
gWHhItLq3sIKAYUYYHWWW7ef2NuLrOomYilneeTA9xtVF1aTv24zsIorOd5l3o2E
MX00XT/gxBuZ21ht1vlczL5850Swhu/i2aQy3x2SlnS9ugh5I8wq1q2oJps9p4k8
Gu0KzSmsHEFSRH+bb6QX2jlpN6IHGjWHOczrvbyf/dt3Cb1Wej7xcene9A9DrQ0n
9n00skyswN1H+ghEZovROptyFISp6k7ta8nuO+PS9Yez2/gWzy0MfpqqbKbIZJlO
zlKzEWOwk3o2zmqs7g5T9bN+0UIkRfGqqTlTu5r/N1LkyFyTB8t9g+uGq6kXLHlp
tIyHZ8Wz30X1jfCwOklQ0e+xG05QNFnZFNtVF8E1CtYw/HUgOZJllJ6WQh6gppSz
twXkt4zc0NwNHp/LrYI0NerXvMxeqm2Oq8A7VtXkzm10FZrty1sEnUb0P1l8izu/
+UDQIXjm1Ebd3MscBS0AzyLOiIxMM4PMl2EnCRIVdmyp1Mgx85Pdc0AVxVc29CZL
t8sOXgL9WNrljnqOFTDXChzvHNUe+Nb0TIa5rp0Xvt8e6gIFl2BJxjD36EGQIzJK
n88ihu80yrb3nv5hzgnILcBJmbYvjrxYjbiqHB4J6rCDvzaVzE9AhYRvoLqsztEV
X0Z8EeBeT287c02bfD2y8RWmydWikUoGKEI/XhPmZHB7u2S8uEPZPLLm+CP3eE0J
SZgMxusH8ZsOKZXATizha0JBIKI2yEazuYxJ5bTU3s2Sf8ydhIZUPo+IN7ucyQdT
tq4mLs72GMlLlXFNEQokmp2C74n6JwWpVqGvhdq0KVzf1g4Mg+abIjCWT99o/5GX
xS8bPY2pcDR+fu8db2LX3FmyDca+19warGRsIi6nuMeunlZg65OV1iSARXbzOVHo
sIOsR0ZzYGZTqhR8H4KZ2Nel6q6W4YxT4bz/g/ooTt/xf4ux2Gfsl+t2RJdbCmEo
v8xS21vByHhGpsOLpJUcEgoT7EnOLFZUHFmFsIVOOl0fBYCUyi7nqqz6taWl8Ofv
eYVtkyQSFYNRH2vYLC8jjYKBpT+bY1eRh2Lis0xSQ4gKR1s5fOkxEk7T3m5aFvUv
2yTqEQwWn3n4plygXDUzupS8m9iMBmkz5983Ej2ldXVjxriFcCKw5UHTJwpaLNi8
LDejLHTNGCaSvbfWDQ1HjZut6383PTFNbYkKBOImpNTxEgSWj6QdOcYwd8upkild
qz30Q6SSBPR906m3+ClWxNJS8wfatQHjrht3y7CI3ng/UXLerrCmCyw3t5keXsPT
1BbC4jdnnnLxiGPg7W7ge8a6JXw6th7qbL54gqCQ7I3PXa85o5FFrpEQlJQDvWkx
y7CSTfaqQxpd85rpCzjbufpDR4MoBLRGGhAZ0YcvEBicj2MzfhA3F3i3kJaNPgWK
5fSqReX1rvVk1EsPHXG0BwV/0ytmwYi3q0rShXJvwSevDJ6qjKC+SgiuMY7k2ZqV
heto+15QSgLEu44JduKS9tLI+du4k24kFhWG1JeKM6vATM/Ve5l64ibGPyuR2gxN
su29apQ0SAjBGIzi+BHMSWOet/k4SVFsLolqv4Lm5qWv2vf+iznlTgHgaJO2wUQU
Qk7SCc/mySbe6nc6VIXAR9DJ2VsYiFpyo5INDcIxF4QxhaKW9uoczC93a+qrIISV
0Xyz3zPEnSlvgAHGUgUb8jg72r+jdeFwFJePBjuvAJPYaYo/WacChil/oyQqyYZH
xY5ESLB7XBmDC71EmfmqoETBpobZagNFdLI5ToNJHB2IUy3vdd9GBywUOOu/dakC
LYeOwrp1jankJ5OpzB6aSoLJIMP/SMKezCEykC0HW8Vkgv7Rg2Ub3BAQMn9cf1Gh
BMFu5iKGJWkwC1WVsdXJvEyJgnPJXuA6LmfI2jhLdL60/IhCJ1YmJFq9CSpSfejI
giJ1rvj7pl+qY82uh6kCZ3xdYDjSPcbGJY4tda7Cb1oO/B7f0XH11STaZz9gb0B1
uuVhVabnWOpB9vsrDlGuvl1k2a5fvfftecSO9QLS4fMzDCcxJPZmEZlrkJCXv3nc
XVqL7dYvSy+U3QtlwK1w22xntwJ8NXhO5Le6F3o8yOOyvk3sYM2nOcnQKRgbTjlN
82hJLhb79EKHjyAphrkBjBBXfowrTd5A9xxt34SdpP4eaikWgP3GJjDYGWLAG40O
hB6XNwnwop88c1u5w0uo8Lprb0G2II0XZQ/++U20uo16WRWRllUxtyt6QMacEosD
5hw6lc7alNDkCOnMUBEUaLbo/yviT0PElqxb7P5hQa+pKbDqnHtfoyjkvsvVf2NO
eF2pcaBLouAAzmy4/qnMiXIVA7iZhRxm+HOj0MBmM0hRUWRzf/gsvl5jgsPxMy2k
U0ZWk0Xqp3+vJycohA5MXoOPdVweKYInFKpgYHzYFQKc+vYfKOaPFj5Y06v8fe2C
V92/cKFspPeYUmU+8m5btSlkNYOWbhatEb6E/n4NUG4qvpt3jNMmq5dIGozttqvK
+xpbw7l1XIgPsAVMEX4thfBFZYETqJSRStbztZxLfEVXCJ1/9o4Y7IHpfeM79dm3
QVmSc/IxEn5D3dXv87aHEMOS4CdDd2/7JeNB4AFTzqI9wtH13JEAfMgQenVzs480
nsi8aINw5RyfIj13tY8vnFr2uD/Au3rdzcIuERA4Rbn6TAJLDL7U5L9NJq2wvlJc
+X76sv2fASHagM8nJPnamK291yvYMQFWwLj3NDV8U58X9YJsvwQ6U77oq8CHBmoo
sL/xl71zxum18OB5yLkUZjaQbOR2+j80/tPpB2PRRsR8p+V4219lZkrFw19wd2pl
Rrzr3XjITdutOiPr78fzndpVuKpclo/GZN9AeEdkhbdj9VCoXHi26ZJHzXuaepf2
pqbSUB5trNXyL5yDhsMybKac4Xuye0NyIL+Ql6pMdVUBajm+UkWNqbF0lO+TXwvu
/fzWVHJ7wAwf6/bXtv+9Rm4Kqhe5bNFZC6ycgtF5JUm6bz4uWdj1N3WTqAmpP3ac
HKcJOp8YrEewutO/VggAcpmV+7ab2FqXbGADhiuAAZl8PuMrW7rkrOcLEBV+iUqe
clxyTkpYcT7TKqHJGO91wJwPS9c5dtMxPFefUZsW2XAVklk5va68YRbrKs7k7X4I
rDCrV2rM5kJOFl7CoTVuHqYZ5GfPISWT3NTuu18TIg0xI6+xb26CqQR8NQ9stJyL
cqGK2M6ancvjCYUMTwlLok9ChKpwTHFusDLIsTJLpSbMxW8sv5U347OePyMCOloH
4gpjuZZNhhvTgTyFX7C4Q+cMntYMASrSXr7FTcwb2g5bqeP7OtQ2R43w6gpxojL3
mcNimI046yiD6UYqYrWuslSXHW4ywKyhSAgIBt/nkE9HBgMmJWBglRwguUkfgsdS
G5cDNa/so/J8zKRSIR0KWIk7pJaaLNtesyrVn5AO/t9gsns+BjivWDwm822SGCQz
FiyURNHK1B49KTjdDvUqABy0rgugO5i7hW4Rz54l5mHlfx6PmVkg6BhL4z19Glrr
qmXX5qUzQB3yQl5UlEyolJCwot+rAWIO7s076jTjutJV2lPOoy15l97HJB9imz7B
CXVKlFJfpHtWYP/KhqTG8ez2HQszyKuPTapNmmZ57Y1RTmN3+m0Wpr32FBdqZAis
e+HXlh+cASwVYh4lrmTFMJ+gx4yK7s7MvyqAZmHOPUz2dA211FY+pIb9fqtFj/tc
44n7YD0BdVQYZNz4dAXiM770IJv0vQ8luRWtAVIpX47sk8tgQbMISl4PkWeUTcMT
OZQ57899nJ+GTbwU6NWji8SrlAAyHYGW0vTBEO46Z6GzF9flFgAx+fpRKPmefQ4G
o7rGEqHhuTLhkJjAAhTz9wK1+vxEA7jAlYYomtxIm1qAEMv7mZmmVbYuER84Ybzx
T4ZdN0V+00PhqMikGllqdc9m5iZ33GoSPb5uN3kjVNtKLgSqtaksNt5MbfkS89GX
0Ote9MNQRrXtprmMokwMyZ+qdKyOiySYqEDUCnjSIkOXDLDe2mCVwPiZqBGOMWBj
TtEUtmL7RXce1LDhQmrPtfkNGEOK3zgf1+XuoSzIZDHGKzw328KpFwBX6sZJYgBh
Cv+RohUYTBS7+2ZAfYKafFeH0piNsRSYivrQy/58gVcgY6cXy38rNaEqvqY5t1hl
oPMJPk9lGS2iUsNGkBeQSFNpbrUEzJAi7HE2XloNPC7Vo3XcIQJ4cK4BmRmSCQd8
g5P6t2ILpSHKupLWmTdDF5OamgnL+zKSi3LFdmZcxsrSXG+l4Wh2jfMXmRsMSssr
5ZklqrNWlV0aLs+RTaRbOYc4k8nKeFoMgqOi4n2z3ca2UEWrEJGa6oCiiVHZIGue
m9BykC1x+LYuyXObO3gqd4HKrY9tqrmsrrA3mk3CpLMtRqD656sDkPbk/obgwnJp
5Z2K0OGjf+eIu6TRhree/ba+O2ARWZO6m3J1mVyHoR5dYnt+bAv86VMA8cgUIkta
edo/bJVrT6tc2wtpjY6+FryqPdYvJw3dpBc2/6URF6bk13O8LVnWHYroiJQTsKqf
ehQeyfFwK1qidlRcEKo/FzTwEYGUdKaBeaNAmwtR+w9sNaxylLWxRzYYTB36Sa/q
fzKXKzcaDCr6srcDZ/lBgpImSF1N98toWBu/5LkAFnrzU1wJP/yo6qeZyNWmXqfO
+VSeK8a3d2dJhK3YsPCraGxxvj2a5TSJRi51dTM1KaIKLqJxAVg+mfu/XeRV0W3g
Xs4JfUBrE5bzPhpHkNtTG9Lya/F9DJXH+CevPZiZsPh8s637UFX20P58qP3vDtsi
mlpp/cjISlbVQUVLnWvIi2yRL4ltJMqwd9kzNHDF0HcOq8eRPHSDE4XkO2Jw2x42
5KsMq08ctv7S9YItiTS/BhWdvM6LQLxacFMGrUnZWjKHTWgV7e7cWzJePZrvzSl6
l3rnMYQWHUzchS/08suXR9KifUg6A666h9XAdMsvqqfaiA/MWo7/ZHdafL/x97GJ
7gn0a4SjifPJpEGOT755UJNAqrTa5j9EoVNqB43PTYdR5fHfY6maGNKKl5IkNXK/
KS8uibSERud7An+Lhfnoy9jZA6y/W1aLYHvzmlMmri4ALGFq71o6WE65pGtHAwkL
mUkSL1YNCd8XFLyY4C3pUQ7h+aoWuQob+zf41uBWisuyZD0Id2aO24QwER+s0mFB
QVGCNZe6HjIZD7Xh2sQWbK8fUj+mjUOeETdVuL1bVQyhOtba2VvN8adan1JzDyL6
oJHezpVDKJg2PfxJEH7ZqWFCIuzvGUKID2fVri2VUH5akedTVr9hS7ny2s+OKVtk
AfV5RO4jPncJUEcR+6E7Ra/7uP8V7ioNfbHt/x/fCPGqEN1mzzhBSGEzi3urC5OF
VFNkBxyQH4KoTv4kzjByJWIhme3AOOVfKHGTfBDR9OiTSOGgCqKWYeE6/gu2QiuJ
9Wy2pM4+ndk26laaL5PXMdeeZHLBCfhNRgp9Y7cvOuTr1TvRsLzuhfGCiWuwNx6r
YrRGNPVxbXDS8ptyNLaf+O8OtKs710Tqgj/VqG3Bvv1Kj0iw+rkRhGnM+uw4fw1C
P8lKiOd6rqEgn3O6FK0NH7OCT6Rs3mr+PU6EeeVz4ao9G+EN5gt2egP/LqwAFHcW
xQ/LVgtbCPbK4XyvFz3BM8yZ/K2kvjTi2238YJSzVA19iVgbSa40A5lMC+M1g84i
JKQfIzD5YD/OIISfYkTqnwWogYmOH5ip/lUSThUDjkbLyO8R31jIv292czhROsBr
mKvzhSkEbS94JL4+c7RRucIpZJQIepqdI7T0PNUjlW6oPFxpXv/F3MNu4MUlZsfb
W8Tg3/75Mm+4bHaPZz7xSqpTAUzf6ajpfR/1f5qf1EFwzfWmZI56bMF2+r0B8PX4
skLhBfXXZCONkovRsm2hZEC3hxPDAdzQ9vXvdzwrZREcaXVbQvHSwsLQ7GdFH8st
86Dff2P5itnU195g53swNSvIz46po57EW6a5CIg0FvLCzEqdYSnDiR5Usi/mw2V6
qCIqRi0feKtODYwM92ZmakxFqCK5oc4prUtMkJ8nMpdmaoSD9d8IXggbwLk913N0
CFTeDQdnidWaTz20/VjEJcHRfCsCu9eKxt11ns4ca7bjCVH9ZFn+Udb441V9ebeX
eb3GwUHlURZhle6GpieOiE1i/vHKaNg6ZinY4K/GtVwZofeV6hDbVEQEkr+r9cJw
vqRCYErlvOmwLKw6ARgwA0v/uBoKmQKYVV7RrzBEERYt8IHGKQ9MoPsZq6G0Ia48
Sp8WmpLEW/65Y10OOCpO66BE23snPeGSF4hj/VnayV1NvFIItJaQyxFJ+DFQD781
7no1wrqYGZglFZGBgAwjfd6My6sKMs1zzZTHBkcsF6CYvyLAplx5A51yBdQhj4Xf
qxaGPkJxc4ACBe3qIoLniDPGmjR+HHwOYYtLVkKuBmWQbnIM2sJ0xLzKn9cetHnT
1yM6Wg7EBF/1dJEAll20Ak0qC1yOFsVhZqGt3NOhO8ZRE/Ien7Eafj2jt17jYOZ9
SjAxMt2ZiuI5oBaP1EUj10Qal7w/dtrSRU45t8AoW3yPhkSXi/M2KTrDrJ6OOBaC
/OYga7sCzWDcYvnt5WZvF8axgm3pEh69XISlMVQC0iotnnlrUpWj1RMhQAVLLQEm
H8gHlitT81vtR1MlvOgayUr8j/XnrKjp9gUca2N5dGnv+QEKkJdNJe8v/SkxrTDk
gF2SyICIAiIOg7sqh25NOVsXplxSP3hrWRQCi1WVYNrFdp6iwlye7Ft5Ret91MlQ
Zhimlb6W0lzEOLc/ydC4vfP0z6z59tvRoHwXlmVCqIwza2TmQu7lPh+cgmgkCqrb
+0Nw7Fw6mFtN0wB974dnlDeMqbS5+6vyVz8Deqxf3+VBGQYggnK+q4/sPpIOsSZr
AFDozWuv0vgKQbQhuYj7vumj+O0f9uZdznxcFI74I08gmOQOOpFByNSPTVfXsPtH
skMIVqXjvK+XeFJuiC4aKvlzILaYIWTMKpx6UbQjHLi0pukBFhu+QcoSDJ0SxDhD
SPJt2pnvLY8sBslbWd5tXpK58LQqXF0yiB2PrKTSTehK/mGmSvvS19hh51QXSd8v
G/mHimyjk1srGJxmVoL7X1pKmyzFcfiC8S0nAh12VDJ3OAmkrACign+eUO/mVN6j
tem7GATrqOFX5nKk2eofGOpod5k8iTP0LR9DLOBTAQlKz3V7tZDzTZsNbywIn3j/
Tn8Re4vSRmxn+CLFVNOqyFNBQYH1As6KB8dgMyjFFIBuUgKO01F7V3lArGbZSU33
ShtExjxmLmUD5GMmQ+kwYwFfwKLDGrwkqQg4HWEhNI3KLt4QNZ9vgxw4sS8EFUX1
LR4hdD/ifc0GSSOdPZHPYFTcmz8zS24v53GebJXV2U1iDaw1j/7g5s4DSGeDqoeZ
5kzqNCtpVRlolXllQ+UJl1WCgZp7AaLjW06eazF4GtAWxecWIBs8piROlv2/hur3
ZiGKNjYPyNfZ6/ThsEHtWby9r7+nv6PCB60vXBqpx4URdZBKHh7ZkXKCQtPoWUzB
6WsCp1aND683hQFMIGinaub4NP+RkK2wfAC9fBTE4/QwamhsroCGJ4C2hPU8yNmY
OkSwXPDLKye3PbKI29WUaDppjxAPojiymKBf9Cr56dHUYhZyP80YzPedDOLjSlg7
5Ctu8Gx8soWHM2n26TwXXUeft579ajQVz8cFqcj2jXYhcB85FYcrXopDnuFFMvf9
xTL+HnJKAbDlCXQdRa/UB7w0fVWp6x/vEKiC9wKNKNmDcdd3tT1pGJyvMOzrZjd8
zuqc3h0qxXHCMYB62m4B9GKRxwkALdTBPwto/RudpD4BqGj7gBLy4sosWRmgUV4V
Kjix0voonMP1j6MFUBz1gKKal6lgtMh/MvOo1PJwM7cm0oBXyoPi45cTPYtly5/L
ba+e8/25QMygLxTkW4F0j3ywG/sOO4wJAVNvRDragnscnX/jC1/GaFykLc4J44rs
fnLpdcoMbHoC/zhNGhZMSWdx3a0CBWRzj/GSim8jlNWJL6XMYzFT9cYA3GLYdU0o
GAao3Fj3/l8r0JlDkRqKDkDIEozh0Ro1yggxYOSAxBEnKzbUDljtDFdidOLsWpP+
qZutEycGbHFz3nSX9hKkK7DVcKym2b6+S2e0WhzBWXZ9JM1DuHjVt57++R5HPz29
v+1f1PGIOdodXwX2BJ0YwYBMAjNjkJQllm0Fa+FMyXXPcE1y9uN956NRmzV9dRyh
TKOI3v8UlZVcZJxuuWfd7IndC5uVihIwRbCkIclV05F5M7fD4htqSKj7El1u8+0t
mrtNmatvsApDcpg4DwscBjxph72Lug7FqK5htOG7cpMeYnzWeyZbfG9wrqjHL93p
6weS1mw2HokBZcsiJaJX9uSWDCegrHYE9xbnyVWPIo9ZRq/WreLGUIuRWiUUvFTx
Zo2fnQJ8baTIkM0o0Kl0gTx4H//LdrYgirp5HVJ9P3R6PSCAVGxQcldy5PSUkD14
bBz2qXkM/r0o3Y4f+ln+QdaayWGXinfeHmI1jM+p6VQGek7cYQbb0w+dOoy1lSxx
+9X1PXsieF5RPzD2itLLfw1yQe9cVtknXA2+Ahhi8dQOx3MI98npgei8AMhfKvH1
5MQvfQR26NH1Gg5QyRxefWEWCld/Ad3EbNWWUYpAiD/jvEN16THUco9fUBCKwmLq
6SmQv+gqfpZvWwM3CJ+Fi88llXD0CrAfXzRpyM/HjNKGVi5D4uOLEWU0LacdbChj
UH+v2i6LWxhRTH1D8AtioW0qycl73jBlDjHNFdnOKPmGpopTBLNAvr+PCagq5VsJ
tR4jmSXAV9W6opndmWZem3ciSWplNTuIdcrRAvmzxju56aHg3fuUS3oJMvqnENER
uwCdBpyFsxI5q0KjLif9wv0HQ9seHmdUlTVjRHAofXbq2kCwqlwRH/ucyjl7ONCw
t87htRM26d+Iifz9ZItjq84cTfXb58611+Qs+vCnjXMXawfbr0glpTtehbNGGp4b
L1Yhsg7+IGRVEqoXskAwK3ilHE84WBihIsOvoiGV3V3O01Okls22RdBegC58eXSG
47jUdI8GWcY/xvYOMhxGNqikB18uel1Y8gC+Wj5GBHynGPWhPZR3mcCykqB8iif5
eOrbLk9XyXwXn/S1/z8sIv+B8Arct8NDJCBPDNAbu2NLiJKKyAScZslJx1eYJd+e
Y5RMztv78d73WFdC0MSo/cLEWMNotCBpHkkS3oZA2OZM/g/OvbBikWReoT7smxUB
BTHYoMe6ATbKN3V+dJJzUUmE7Y1VlmodgDKQOHSFfKH+s5Y5Rney+tg/Pqdraj97
47vGyBD4O5eqCrArkk/i3URkn1N6cre5OehDLcxga1wRodrpqYPd7AGUlizyVrLJ
b4Hhqq+U577vurnFWVMw4x+1E+fTuVKVIk9clOm8pIFPqRaCS1BrOs7B+7ozGluM
PV21A/FMdvQGsgVJu7N+A+6wVltaDS9okTCaomRvKtgg6DOv8ak7y8r8eWNHiPE6
4CVbG5YkfL+Hgzpk/K/DRnQqo9ENFSRjI+OjjcHhUOekz7YEBKdlSb2dKRJ1yhDj
t0fi6IAnai0+uuLYXkslF4B/pTTGqXC5niUb8MUtLhRhR3pUa18+2tYTOr30xp7U
GJNZaHk4AIq0nxnZgeZYcgyOPIGliENW8PNGFcJ9pYaArd9/vicZn75LdAsfMA8o
zf21ceA9j2JQxXcCPuNRDAuC1RurmlhiLgTqGPguEDbiVTXzhSunMKGRXYd+fDS6
3DkGsRKuDSV0doACrkdHWKMxJ91qEggkZWPybNlAAupPGgk1KES77GEaOzMzTKeQ
7AWtkk+xEkuA1uA2Vn+mmpXevVkmCTiCW9fMnO7xR5JcvJna0B3O7agPhdi1blBl
+PUQBzVaQWXF3wI7UMTAsQamErlUVEM/2+tDCyA/RWhI2W3IliOPqrEIg2SFb4Ve
KAgQqxjd8i6tWU3KM+aCUl8FC9VeCXXF3pp+s36wpl/ZCD0wEKyE5vIhEFdtIQJ9
fUDwoZef0mtHNhKiBB+UvDDipEYmyyuhALM5WXN86DD3QC7TjOPMvitsz3RednSC
4rR9AyIj2Y2WH1GX8wqU3ChNbDa9ZRWn8HECTj/e/ckYZrLjgp9hKwIJkGgokVKm
XmlucIAKrYtx7anP4Lm7zc7qzVqDf34WEU4CJEXDBo+680gAASpzygCJxQJOumo5
4n0LF3a5+m/kh69R2FsBpglykLMgjZjC8GMBWG46rQl/8Ej4zSqCzuhrn5NjqDd/
RHQdNXo6CORMGj1UGky/H0Cl7TJ5hT3QmH6GTL+SxyJV5btKjm5FVj/dL5CLkPXV
LfTwXYySa3ahTPV9bePJsvpnBNDiUF1Y0ZCNXfwc8M3n3ERDWZWrQLPlJ2EhHoR1
Xqdbhj9C6MoPoGkKVrbHLG4ih6zeC9tC6pZ9QnZMXIiT3r8OBBj/J5iQCC14hUGL
YTBvNFoyFmZpx9lCf9MqLtLeO6NQKK1w4Ja+CbpYYrjXOHEdKg6O2lIFTOjCPWk2
f/WTIxtYvEY5DYUj1J0OVlJFH8jaSpLAHrXl9nS3WhyH9J5s8cFuH6d0GSCns6Ql
QOockZnanGxxJg98tiuNO06cu2vvz2gYKCU6gH/IPXOF563AtLc362R45kQCuhOW
vm/NRBaZDvMbNsAKUo/KRLA0FL+NAMZlvzMnaNpyDyw9SmIgh37VhB4MrqMH97aF
2R4BRQJ6moWWkgm3/dZ9wRTbuENZddczb/kiwMv8w086BQpYqLOgQTBOTzu9b3Oj
IeAoGq70B1DlpIWvCFafvtYgnD2Z2EBj1kaG0PaDZmbaA8k21yNnpo/xeX02By37
FuQvlN0h5liH+f7SQ5mhM7L0PSRp3kUtIyGzNORJsVCrN8PexB1Oc6koJGsZ9GdH
a8VXykdrCtAJGWlprUKPr1tAHlrRwA1IgDCGW6Zb8n+bFO+gmXJJKNHVIq6a6dck
47yWPRz72Rci6UBq9F9dYIzRHm+9qLuSRpMw9sA6NKrDtYaSyRJ0PWwTlzE+xp5y
0oEF0co/vvp/8ll8Bxy5kyKw3RYf3UanM2GUp3qnYVL+/UirUoepCvmd6uPxVVG6
vt4cyUk0Mn5dRRyWDA1GxJ3sLnCPUEo+6tAHp5NsT8NMADUKDm2Qq8EZjAf2RrrX
nC7MCGWiEKosmLDlpn9mU1gvLdgPgeUcWmrLEnLgJlOBoLkRRs9ZAmr/0vU1PHb3
wRBF5cE/08fXX8tc6MBRnsfPDi7RaiYCwSLFoSBvTpOcu5JVzhq/+aQ7rMETGxSY
Ws6k70HJsFcIR0+ccsvWRfSe29VSUZ0EG+75NV5A1iMdzdkA/A4ZFY06Iqmy4PRx
VTvJOpTd8LaJGBFxWkca8iH7DP3qczHrhm1yZh/FL4mjII6SnCEI9BGpxWjZOux0
12pWD1ZIkbbdFq3EtDfQHd+Oj4OeJCm+CmL1q2U6T/DX67i9ND5lmyp9nuOfcKRQ
c5CRviNZD7LfmPyS3B1pgD5qWqQ5N/yVBjeP2C70ejsNV3q5+MYlXb85E37Qlo9U
dbyRbHXwbXO6MuE5+VsaDrOOcyK5aXBg8csP+1bbjRdTyvcF9jOqe7a5kqlBLf2D
w0BybRauUzphauzuInFugNPr7aNkBn43B8y57QeEiWZesDosDZAUK9ebhQ/C4WTz
u1dCGmWJUIuJJTOFdJn3iuqnOZnBY0oIDhPLu0EFjQiu1EyGIDrC2C3tcnF+9u/K
8bwVDZiIvwU6wxd1ZpkTgKti+CzXppBejE+NGbN3hX4wUhqZG2MgypU/0tP+jeAq
ewig7iZr9kiDvDlpRpP+Nhe6pdPUaCsrrfDLUfG76hlwDxS9Wx93QQfEMWj0gFbt
9zsscexdjXYiWPiJAPfougWKLPNPZJNFcsZC/1USptnVYGFYCBvOfK7VGBcOTnuM
dpbNTwrw7MkEUXnNnicPZbTFUHps8k5KXP3dNJhAbPoG13Dzmq3p6yGIBaovkywp
d+Z5FovzidCxT748MyiqJXC9kSeLeTGWs5m5lPv59ZlVfJqGu5lDSm/Df3WdaNdN
w2fE02HCA5Ztph8cJkRWQzl3TFsYKUKslDGPNENaTq43Pb3HYYFnKhbMmye0m6uz
TXdBcG1whHc8TNtlqpVu8ZU0dyKv3Ho+Xywr6r9FiEWUOT77pTZ4IBCBFnLfRc7H
YI3w9nIkTGrX881VP1B3YkMKbiqeIE3uK0K7BTlG9EyAXIOjSFpvkupNLob/JbF2
6xHf8rXs6678XynjNRES7H0XilncD32Nm1hFHxyXO+ykyC43NE/R9I70rRtW2IjN
6H6NSBo6Qc1uNRME3kskBc9Zt1vRPcORCvkT2ZY3yaUrMa8T/SoEcd9GTU1g2TUr
uzmeSdaPpGpMsaBuZgM/gbj4zeLINIsytR53b4wN3G+FUuYjrBLeuCLbA0AuRr8P
4XAj3ZrTXNS8tarUhIwV1bvrCq7l1Wlzd3GI9AkKDHj9lQ3g8QsMygVo4DYf9t/+
vV/PZdX57rfsGFpuwxs5sDbFXEjpteZIODH3elpNEpsriGRaTPbZZDIzvNpisI/3
a/QvUUkriQ2I5RdjOiBFtHmIrhVszDHnklvQ4AAcHW2rWptUnkvNOBK839p5hTYy
qyjEBK137zaiM73gI/KnXZP6ag54nrO0rLLBsZ7kyUhU5sjKOzTH8SqfyzAaOA5f
m5nAvbDvw4XleUQDKHnP42bW4RkKitMPLizbRoj/Scdb/nkY6yM4Bam+ROrZRRpZ
npoywL3h6L8N3TYubzY2eMok9Ye9qHYjrpG09hpmKT2pnjEiUcaoJkUjEEJjiHsc
v5tCWLkoV6FBkt+mSn76TnWcYNqZ+9O6fO+hZ26cOQIuCpsGL7muzLWgHBsGGTAG
gG04ZjqVn2LBHgP7/I/PcFGazw8Wg9Su0ypksExS74/4/Bzu7j/wQbajy7Jnly/U
zpMuopINPSNak+wutJfts0N0D4m0F4Z+d07vRrufWh4/Omtq7aMCza8U7TkmAQg5
tTok0/CWV9ZdmAGXZXhcv7is26n4t9rwWCjmUmCpLN0TX8goDCQLlXgIIP0PcMaX
7nFqxGOy1OUfwakTBaq7MlpdhOAH/zlorf/dHEUhVFcmChSRP5ChZKfw+WM/JVAS
PmwpOKoeMFQhoS8AHYbBcADQIw0/YfWlZ+rZ0sJmipPnGPIUXPlT2fLKSMb60fC3
6QtOqOq4/D0Kj3qr4oPtDgyg5s5jpu3ifZ+UY4EMz98B3Z4EfjmWZn1RX1MEyYxo
SSD2H0DyA8Vh/PDYfxXOGKSSWCV7XM1F4WVgvZ9zh/VxqubX/9cysEB7t/DSmHrW
hTMtHlDecm20m34GDYKCN+1h8cfSJNQXdqelDHsWul363S/TapBeTrP79u210e5j
4RSzmRg7uxXDrSK22xBtX6dSynpx7Aa1AJ0O/IZy9Yl1zKfWVO2wrhiaLFsK1909
1DnUfgvAtaFLf13XaJ1ClpVaQYx36NFWRQON1L4RH4LbIjuKqIxv9MM9h27ExR42
CbM+pfYvQZlLVY+6rkk02Qiloi5N/BtRo+eM/Mpc2DXFIFLBIzUsyfaaJ9OZcr7/
D7lppcNqu7kKopg5lnjXeOYAwjVAIT0Um18E6/81szmGzIvfhtfv5xwZAfHpBuUv
vRlN+8u7tc2NGDex482iQjosNAwujC+Pk9pvuOYUhIGhqzERIRcdfXXaw4JekrME
zbU9wlZTYFab1/ikdhqbCmppGRV8KMUCmC9kjcTWhtzso6jUtRbLV4W+QmFuFO25
J95Yykk8fOm5lAoVwYDKFDCAZ4cH9um30OpQdddieDGizvzHohUNWZm09FNd+jKz
7Flyb+muANHoQchMe2jzQ7W4v0ikXLkg7jnVSwmki3DoOg4ZJQJ+AozDUsEQYf3w
XkEPnbc+hX/JdO2v5bv5h01MWZ3ieERVitgT87PYt8uQkvqtyikvqSRUhBPPbrie
pbV3jBBHpBp5OIYXDjDACtxzZrFeYgxaqLrCCAaMIBzabdIDW6OYDOyLqW/AJ3xI
LGbxdm80XXL9eGVO37uOOt80cOYQaBIrtI+hfXTEySFG11cJJSgMZ97pG4PCxJqY
wA/NnU4lQGnzWaj0hPdPjymotSrnheUitBX1fvvKZrnmjuqcSZUpA2WNchpRPcll
uhStH5P1JNsnbVD8hTUyzDTdFtqf09dhLuCsIiN9bsZ82+GzCawhNEsnUrsSLv2+
xt1Ad30COUO3eCrI6w8wqHptogQOKMOMLxnIQRM7+JK60C2jUGjDZkLnH7zgJ81X
jctyqamnZWKMrveOOkTvwGOxpomEgU+l8R+LDotLbylT6j3V0cBBdPzKj0SP0uIO
qXCvBKdKR4e0E3NK9TjGQ6/YErqcLhinDaCh3hk027Lc1UA/go1unbsQtxZJS0yX
6dcK8TIxBeLxhrrz7fHDdQLiLXA1IIlBY+d9r0nKp19Jxye89++0VX3tI5rz9o2l
YKp69A0nYlZEwsEpvPwCKxizMwfdH5zbBGAVyYtqtcfwQfrId9+C87KY8BnyB9ED
VUrjGKFtphNVb+VeC6hgJ+deQqtWRAFnqWU03UXN6gO10J72PzcKJVELPcVhP7As
0ThW1q/PuCCLRoXI8uXXscVlsjOmsV3j/YYr58qqymojw2tfyYbTAGRWNCVaUWHD
UbpLSRcpRhJ60hFFkgWJXmLDIuhQRKCgiEAkqnpXoibNncBNiNWRcqwqAGnhVuW6
PpSX1H/rmL8rBxELq9oilOQyETWrayte3auuN7/I3MNyXlrHwh+uBL5qxbCNLnvh
f+snc7HDx63a5P7LKbdIUgptr3gvwSLPjMOb4ZMUykm8GzQgwrH2SxoetEd6F/Uv
BRPflyu79XadyWDXQhzXC6/lYJJgDUyL7iSuNSQA7a5kISQZ6COpVVRiasbVUrkc
+SoLIrprJ6H/ULY9A7XuVgJnBPcv5XvSFPh+7DEvkeL63zVwzScqWxI4IMmgTXSH
weyVDK9LtzmdSR9jehVpuRQJEj0FjCqxpeV+oVnEBZTMxtUadryXlADmnZFeq1dl
xrZVv8qSqt4nlaluZ+cL8/ghl6S2Kl7ySB+m1w4DALnHqmVxWrbeUet5RSCOqsVC
nxjVld2MmcIlvJOzch9TP+c+6bgR1hAmZDHq/rfTJSzMblpD9z/E/1NfKc5ldy/1
FZ7jIYd06rlbuQMzze1ijLSrpG3S+epztbaPSyijDmlgheDwtmULzEtFgx7ow6Zt
55S7u8LB1Dv9YwLVWcUG1rfSQc7Rf5CVzZP6t+JwJpIAdo/KpByaENrFEvV9z7xM
FUJim1lcrOkWAqtiqIGJvAb8b90RuSRCOyRXTpfvt1wl+w98Wv/duXx7v6cw1wGg
rujjdJawZP066Zaj/JZUcp0wzTSy6zkmVfurZv3jxWSoO1hoOwFV3YSAAZ8wL2Eh
4DgqJEfNjkkTKEva4k+ukZypz5cJRsBoiAs8pUXJOxjCQHck7RAc8TdvgFJR6w8k
eL89ZfH6BpHvWTE8sWw29+raMzOqE8l8Y6QhZtK3IZJFUy7QukGXio0I+K0PR3gV
2h7hZ6FGESAGZac9mu2iN8eP/SgQUFTkJP0qUcBE4R/eeODntQyxdT4cCJc9GKpb
+CKIuPH9IbWEB6ZPgO2tNNx4hYoA2L4BnZPiXBUO5bH/YKCCk2JUa5juNhK6qofr
d/yz+ncu8wJX6Utd9hOWOaw23zCkpkkXET1dq2ROIdDMhSvVN4OyxHEghadfT/8m
rcULeOwJ6nV6ra51B7ioKaivUTcTr8+R5d7KkdP7DuPiUAegNtxSo5TedT/BKC5w
weBgNTPkNBJvtp75RH++HXFXo0Qxg1oWaXltUw9cUAsRtIBRH39RMsJfPQ3oS0ia
b3PBtVgLPd2qj0tItkCahV8UcKi3t8Gq2oZyIVt8FErkdYdhLp/fQB2HNx56M415
R+bC+CCq8pMmgYBUH5lBGj50Q9sYhdBktClUEfb6z80IL876LC3SOQ0ZdIgEIAK9
SWd6cF/1TKRxiTpFgjBxQ77slK2/qWGXLzFdFNKizkFQ+x3fJhAq8CIFuxHd2O0M
4MOhnyHLL8RwJZpW41XTQaPamZe5bCvpvSJFwasHWDyrDv+12h9CXYeqtkHkBoM7
YUgfNd952JoRJEMJnOKbeVh3DjwLryVNfdHX7alzDUIjh63MRWRWygaUlM9pDT+4
mnOFMn9bN0bfDqLxrjCXScQF4HQTeVFI4qE5g/xOEHp8oeJdOoLgG/bMvTU5l0j1
Uoj8SIPtGSxNvtLJbaUk7fc2Dqv+Q4D06tZdBqQQSALhiP0PFKkX4gqIoOWhc0jN
mA/7kYKJN7dVb7mc2ShzvOpcrkBS/V4zXDL+Tk+NM5m35VWzbXjc/CUkl2TwrCfH
McnMnWsifZkRZJ8Kbgg8ofsKjyCELyp2OBmCF+5/GqitI9rUwmEZWGH1MQbT3O9L
8IYmt7O4k2t73Nhgp1d7zoZi6JnRhriQpa8xIcvcBOeprLIWm3N4cUpvx2Qr4Ufx
7hwzU7b9Fiv98RVnT5LEweg6azH21yRGNR7ZWLuDLqo1pQbmdvwJoCA2lZGkBxjO
I+VNLm6WUQCXMhGuqgBcxHDrVXFKMTitDxajKw05EVL8wr/hKTy5z/nYtqFjnIOK
ZmWks/0JKzg5FSHpMSh8pCKR0k8NmvptdvxO0/MNTFSauUuFuKaYd8Wq8rDBE52b
NQ2yik2ZzIZQMvlKGtrsFHRMLzcuAg8AwsGlCmXIRghvys60MSFIjNV6CX4YTm2V
EYpapBukbQwAWd+nMDBGwf/YoJaXxFSVn4SYXhLpSITjBCdu67EtDpbeAhYcE8W6
ji6yZVOmesyG23C2D64v0Fhm3n+YFVsoUY6j/Uabe/sh3s3v7YRbrzJ7YfEPHYn8
aRhbOLnPmRbIMG6fGKUsvYqROc86jkJKuwlKClVum1VvUu3tNCRGGTswxV67B21Y
nPWNnFgabaZ++jOr7Br643d6MnPHhZ0WCczrj1IUsFhaD/xVwHpFxybTgo6F1iuT
Cx6jzP+AuIJKpyHx/zlexcUj+Sh47pW7Pd8lGt28ave6MIcw7CJjNDyR4YOnvcK8
MuYibCJSOa/LoW2DaRBwPSOtiNBnmnGGIOMC5ihx/50iCkbHs6xq+0AGNLfmPiXQ
THjX1kd511RabrwK5pLu+G8sdspXxZWgf2pjTr6S0bG39YqZRdtrJs9S6JRwx2FL
hRUpzMVSTFfSpFX6LfZVfOo7pp1AMLnweqzj3cAUVaqkkdJkBAST/fg+Ht8xrhhN
dZhB95ImkBrMYzk9Px8sHaKgvjFmx33lHiLkiIOd8s7ztZA27XGT++uAapLVYzOy
VoS+4kM0CUB8iY6e/Ni+a5sK8XWTEPwtgCVg3+A12HYMyUOuC0VPIhw5WVRDI7Zy
uP42in76VbWRQT1uaMvRylHC2r9hpRK9GWeWr4Gti4N4I1903WnKTTiH4NynAbN7
e6GS+IxG3xY5Uu/sGGn4eCRNc+i3zkFKQS77GcmZKs4XTTB1AkdXRLQqvp4KGeXq
XrBlGQwnY5bY15vVlWAzWkMsITNOhK2SW8LrBbF09KaYauZmf8UTGoP6+j8+sBgm
MudL6r+q5DQpnOrGvsfvk0Mb82+vbf6xD4lFvk29iAWSg6Gc4GZ03Qez7QYRuogD
kOhhOLVjyWJoA4rlrJUXQkBHuo19SvJ+WU2fYa4qMcx31zY5fAkk4O8EgXOES63N
Xp0hk5xgfXHZuD7Y2kVJKIzDStMcpdXhi1bw6gkDATHjLOQ2DfPQ+hHeRXzS6LSG
3UeCWRHfd6GPllirGgwJKUb2q3VEnwJDVoOpOOrJmT6GYQxZyExTrmEY1rbhygU+
CLWg0/mAGSVH7LI5DDcA2GNTNaBbWhrQc+jTzgnPZQDMo1/KmfRx5+KtL9Oku/le
iDs3eZfUMVFZRxjYyr+8yZ4HZeQMuXDr48Di8thMLRMjqV1+xTWWc0lvsnjGnJMX
SnzkKcuCghoHFM3qMvFCdGDX3SzxglfC2z71lUYpdYTSJpzFQi44JEyjf1gOJTLL
Wf+MbEr9q+75txCRzJn98lV0/MozcCYa+LRep5zLJMsfiOeF1pz618VSk+rH6czF
ADwFrGavvAQKuIysNAT6W2ekXXOXt2IasyRH4iUu+nmP+NrOLs5rY1ltctYV0gLm
cxboTHTXP01yWWC2fNTRJpJgUnnYn7b5rD4ek6qIOuO2OTkW/I7vZAjORT7y4Lu4
SUGn/b2gMH6f5f0OPpYewRIyWDJYPaZggopeFYKiUj0SqTUmJsMVDzXg+F58z8Wo
9LCioSIXpzgpM8WvODSakphDOdqiXXaPoX+ftez4Dnh3VXOZbg+vHwZ6AK1FACmZ
6VIjU/s4bne/1+FEOFEqLbCjY8oWnwS8i9ns229Gf6tCnkle8NZpNR9s6CofLEfV
l8Xy+GFLRoOUJ/tG5BcWhp2F7bHlM8lAn1LkrJnMcorvcgvbm5FHuTqCpP7hy0nm
7+8nftna7LhFUni2kj8tfhejugSMhrH4UHJWyAJ2uL4Dyh5INTrvW5ewnXioiAdO
Jbqb/nGy+9rV7p+7qAIvrmNWGOjecdnEdSvmfBE/UwNDh6W8DZicFjbQjAdbmO+X
AxtJG2GlEndv9OcRrV/8tQ9ftnh5QrukXh82hhurDBxIr0TlF3ICpBxKl3X+0qV0
UfTs9FH4r4u0kpHe/TkIL0xbMoW/NPq5mqDWYjGPexUJPibq/b/SR7up9iKCYkzN
klk+hR2MiTKpG7PxLFoG/8ao9OOasBiSsBb8j7RHK4fggD7d8dVHkEup5vo2cKOU
EJOmwZ7P6UJe2xyjquN7TtWpPQfYWp1i1oFNf6HjFDLG6y3c5Yr1I7bXezpuy44H
hzjJCpDByatLJ0kSsquxEKmGaydpD82j4nIh/4SNfrgzPIgHdgPcDI7J/GPQM14F
3xhJXnpxFmHHnoKvijrVJ9qu5GZPZoSonssuSNApNa9M1NfSF1s0tLM1AJfxrzSk
KzNduNUSNimsCEUYdDLAnkWbpeIrPVAr59ZJXWIIMD3oeDBIQd/rHwO3nYvYbv+j
k3Hel+YV+3sYQpKDGNk16nwFyJ7Lu0/pIj9VFdCIVmtgm1pg+0jAKHHlSPnynCMc
HpE6L8kwew7onk5vkRK+DmmsZusU+FksrTxo4yxhUAzxgJwVM+1LBiqU3kZHuFd1
xnglTr/FeBzBFgq1iWo9xg3Tv7/vfrRx5tHv4+o3VDQbAX7KFy4XW02pBxp50bk3
EaQkcA+QMz8bwRaA7yGpRuYCsVRwbZkVUaZ7cWrNobxMCLPd7leN60cEbgiauH2c
wDF57QBB3fjF2qg7/JDutb66Ex0X2UKvxowBhEuBwVYgNkwgx9CRePtshdaBJuAc
l1xxZNXcizXQdGLDD+K/WqcxBU2d+H7YV649WoyQOBxbBXjOgB/LVHfqM9TSjfWL
kJy5hWVWLS08xC1XWPTKPOf8hJZcvd4IzbvaAjgbR5kDjzGiAGS4D+E+75aKJXm/
gOadpu382DM+HWWF0Htew44Qsxt+rHmiQQf8jr+hKGjyU9gA9wJg4fW1TV5wxdfg
k96dTnnBOBN74iIqQgHUm4+2GdRjc3IqI/r0dXML7HaV9lRhkH6v86Cq31s/Eq3o
h3V61tUlR0AUHxFsogGdWCdXqdOvsDOBtvcyorWnQBFumjoAQhQYRJO6oDzAcWDM
MgFnM54qPodQ2S9eoDLvGWVGw7uEL+y+CAwATzw9UJ8UeTcNBqXP/EwBXaVjqe9O
svr40nru4/kcOiU8BXdwBjlnJ+dM2ejb6pNV1cXwO6U5aEm2rPteo9EIFtTwQHUw
8fb1t/iE3s1sD0D1aVZXk+TCjIMneLH3lI5yd+aqDOtbDRPtaHLaSFR4+KZ6TBpf
QSpHIU14But+vvYWrRXRHh0748pkCW5C+BGc8m6nmn/daQWBTvmnikAgQkl8CJKu
8imO1xl2Qsv2xXKb4F5arCJUPiToCeySjoVrJVME14eWu99+GsmbiJpxZCvb2xha
5BBtqStwSp9vBFx9GE7K7Cr5f/ZeK1jlO41bF/CE3garN5SqS5mmtnAaRWmY4ZOE
49g231QS0AwarrhL/9cPwX++J9uh3QlLTYizlVvrhU53jURWnqvfB3pVdM4gvF71
a0w+CvYgIfpOJPlk0cceobZAlTKrggFws0K4N4dxIXLkB8lzEzKoO6uHAHorHSFb
zagQMYJwbuHKxmLEv9G9c8wsuqZvwUuKx3GYToOhvC02F9VRKq1Dl0ZmebJE0kKe
loZIOkrKx6fTMgoUMUR0dnZiIGj6ka82948B3lGgIbaPR8md5zgjK0OV5yA95wQU
s/dVXfasHTJdeLbVClfFiInRWgC4BR+8UnaBalATPk0NpOIckX8EfnB4yZd18aBq
TLB6Ry75Xh/zrRgX/wslYoy2eHi87r/fRzSskSpz+OK9HKJ9fmxh1N6vZGu9BL/W
RAzp+hAycWuv4pwBA56Qa0ScFCADIeER4DyH1ofiz9RHEOXBCR/pU/5vzqsk7P8B
R5b0CNQ0Qf3XiggnUXiogqH5ntctJMWuYkBjYpTJeqphTzKKnWZG/inzc7DgyApZ
p4Lxm4+jQU0mK+kl0U9pcvqYWZk4cVP+d2HL96CS7DkTug/JHOfc0mXPpDIWXk0I
8zW9LmT/fWv1Thv67CvB5ZgakXYYbDvwidu0sZk/yqoVAwpyRL5i6T7Dt/DpqMxc
P53jedMohhzASXBMICYvuVGPUKp6gB741mQXn7erNKWLlLbANJ6qfcQIIdAefFVl
haW7KkPOTqo+O8bZTukrXvWIoktk7lQI1sVj4vuqjF99ix70cQ5hrLIMqPzHBWlk
AKi81vnqn/PKc+VZsy01R93QjPgqELu//jdFwa2graUex8sAZxcVQb9DXC7BH8Sb
NBCw76oUoYLxaxezLrnygf+x+wgAQHiXcXov0j1z2sPqje4rX5DR5DBr/ZKbJgHk
2QD13VnVDnzlP5Gm6f84RVU27anOWhaDuJAvBbNfYw4jdqqm0DociyFoBOMCGrIR
OU9RdSuuzoYXdpTy6UVN5ONQttYetlDuMRriYT+sYXiXyGLbCjTWhEFEFvJcO6CA
pG7/cUT9FS83SU+iXVuw+cCrm6OHnOK5hSkdzhs/1kf1jYW/FufAHVKBPmJxK/b1
/c4Li8X6/+r8g3Mjk5Ayx/7oaJJRqvrNNAVf50goOWqXlkqtjGDlgeGrkXQWwBFH
TCu6j29Yt3CrKCnoVBQJiic8O6/txzmoXgOsWfzUDHGGvWGUBs/OXH3xVG2N8+og
+Yvc3JN34sqMDOJJgcxThiMBlRXLhps3wJ2Bp21pEwQsJcorQG75AADfhVB6FCAE
bUYfrh4bUh5AxdNldSnnWqnFowmVdCTXHYv+pCUXrFNUvTDIMytiERpHnKj7F34M
59C+8yBAVatEj4cZQso48Kh0kNK47R5cLc8hBUThSRlNeCNDzqZmeEkkHPtNNAcP
4GLOB5IDcp1766bXFeEGjwRvE1djDbNenaT4i7TLfXxLia5HXQXFy0HN+EcS4PLu
DCiKFm6aQOLaekY/CF78OTvdBW3kGJEZquTwvOk1TOouhqGveqpbEv7bsr3Okur1
veweyTfKyY8Z+zgY45k6fggBvzORmAp4gfOtQdQQ33QmxZYbAfpNRRgsQcczssFf
1X0sAegYHn88dcH2BuzmFHDuviGcZnTSUFHQDofzqPLovr+yBMc+4NjAp1KXdJaG
xVC/3bTW4cG3dMX1JWhg8vuionI8tYdinMkRsqO5tbBgrOwtOR9/AtM8iYqZ4xvM
vwhRnoaqLMcxLG/VYds9MQJgkUNaLNQz82pmFz9AJtMl0GBMtEHqfzLtVEHPa9Sv
F1Lkknb6M/oIuGK/+vcla4PN0zy6gaWJlk8UCoEr1R9a2j1wN1poYRmX/ZEyIUFP
2+qoWWrqu2EV1EzOHZ9wL3lrBGf0j75hopPsSAk5WUTCif/UVYsQq0p79ku+SPlx
7b8icVdjmD1qH7WBJ13ywm22nALcxu5xTjbrYpI8fcrVY/XAwzLnuVENX/Ti5KHb
P/TMCDrc+M6gwdC2/pka0S1DrvSyLy1XiM/Mgr9Z1nr5zaeoa+pM2sX1Xai9vzYx
/JGNAZ6HDumhENwfwDBSMgylKGn9DIwyqut18r4fHpBLcpRCAECJYmyaSMymu9ie
a0/7CJV9SHyugWOAQkMmfX6vSPB0DumFu553edbLczb6quD0jDpd87mERKs5D0vf
7ODGnSC9HgseK6tBO9SA9rGPpQkXkcVeHBigNIU8mwCmHF4LzuSDtjbeXzW31xWA
O/y45TPLdZjUr/+1NfE3ffVOk7UaUg2F7zcKaKu7PJY8FdxENkNHnacfeyN4ob9h
1+m+Aq8s/SMDf5/w4ylLvd85vT4p+CePQaMVVA3cPLUMkFGTgGl/L9SpkdOZyQVT
axlNALpSzSVK5Ugkm5Xzo/xoNgx7ef752reeJwL8ExE7ZkjTGMc1F+Au/n3cVDWj
hWxom+NsUImaBt1bnarkgGYWj+No+6OPMOqSk5c3BpmXCzM5Y+kISbOxpuhwxN8I
1B8bjP8LqY44/L1qRQryfB/6kwoLjLHjGEaPK5ECkSLSMdCX4ypw1/hFYh/79sSG
/wVbl0m0/cdfy5/zNVpNqj/edNF9fvSq8hrvFOwUXeLvvG19X3CE7Thn0Ac28mTP
BjkUW5tvOjlBwH56XJznsBvcg6g18dy4rydlhJ+9C3VxUUIYAq72nAl1e664IBxc
xcjgLi9L737LlhZmvU/8II+JemLaUJYLtFD7IZvEH1O+IridnHIYb79ca0ohohu+
p1BmKXly4y8SjVFPdFHAONXRRdYG575YeoIbyWofUU2PVKmuegEpe7UjDya5b7O7
JHkc5L2kAmfTJLhHVqRFXTAMCcra1ZpaOhcC1K3fp6WpIho4CR/Ue+lJuSXmo4kB
D/yBj/uI1v25I73mdK9QT0fnz4/IuNIdJpUtO8/OhFalGBEH4SCcn/YoljLhf0K2
VX4pKGJJEsXh2VlQVJ0g+rSFxDE35OIP1043THQz5FPPdW0wvgKaWmGUCdb6HL/i
0p06wWbVn7BUH2WCELljSUaNQQYVeR/oglrTEUok9jN+owuR2x0o/KokSXVJOs9y
7GsGvQP00npzla8ONRpkP2+1wakTuj8PEQMh+5GbQZDc3zzZIiG22XySCZ/OF+Yf
2pWPCayir04RiPSJFu4iKAkInGGsiTAA4bb0epQDZcAip61OW/x7ky018+PfUvxT
2IMdUo32WNEzNfGl7xCBmiYvKRBwylDQXfn28bJa3OCbMjioOMRVvR797hzZurkw
abqUcdqZdNafwhKGHwkSazNvqmgNHRwqBjW7i83tFgIWc8mNlRe/wFYfuqYNvUOg
tO0Jklwl5MwvV8aFwPCq7evsqXY6tlVkyUaQVH1Djh7p4lXCW2bDSM0QPQBo5K5R
LFQ4HW5SlofkLft8IM7k9YFrSNh5wunQrT+PZCkV64/eOe2cFxrTSsbpHGUO9yVG
CnL0g8m7UScgGiw9WHjpEs5ATARd1aeef8GjiXrz+ZtOr/DlSmar4olFP/bnG8pU
v82uA6A8SswpBaRo2lS7SIYnFS29wV8XAK68IfGphF7MWO7V94XIisR5US1KtxFV
tlf8agNygqcfDSF6CONP0PIhaVzp4UzQJw1HteslXIR+ymM1qyvJ9JD0qK7uDFEG
crdJee3AXahZFyoX0hc8e/IHMKa02pCa4RMhIq0qj5t62A2YcmwQx+oUjnEOB8/Q
HOkI16+LEyRRP5xQsYlJngCAsQmODM4vhvY9pHPWLjwoSyd8h0UjOhz1kwI0PFUX
RNDe0H4TfZDMJbw0e704jyqjjltA33zPXKHvd2zDcJ+dJtspvadrni9YqXOjnxko
T9lXciKOYsbQtPpwiqKg+pqiqorQ1pYDBTpHswzWtnQ//C1np/CdwrnCrERHAqVw
2BZ/qyFDME/HZ4MzOVwm8MzPtauYglk5+62R5DN/NfilpuvsJlIBwh2Lfq4TO9f7
8eYyvA8r+R/nEfhNfuxbckM8RTIfEozCdn229nnYFh8E8mY+aovoe9owbHh0cbRG
XTtfm0DKCeeAPMKKO6Kyiny6snr0K7laQjo3iyrqv+RXQLHpXXBnUWdrCTCQ6lMj
v3Idcoj4LmYDazQvRtBUXg6Yy+LcFeiDpFYns/ORQpZu7EmBZiATXua3v3eng1ui
XIxWu2Uid0X8F0q5cTRz0RG5X2DdCKbW2I8toQeloiSkvHDp9B+s7FUyhmNxBbNg
OvTS8qheean9cpqsr22QKVF0aQq/8hbi4unE2v4E0Ob+qPDvIc8bFz9mfrQd92TO
2mcT/HzyvHslHB0SGw27TmO4vYzlAhOnxwK9xIC0nfZiWYNJ3hxTjEgi0xd6VZz/
1tskaJmGV7OTPGjUzjIwqiwYIKgndmi8RrdYlDdA0lZb6QUm2yDu04/NeiSzGNpI
crraSMpyx+1VeM0XwBnqItiVMb4Fsgp9h9Ay/t6VcYxkCC1wTDVibX62SkLomgww
Q5L9+OAJ4NckM9MGVdEv0xl6660GejtGTVgZw7emKL4=
`pragma protect end_protected
