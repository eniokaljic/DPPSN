// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MnbJQx1nGqkHixAURqUkbYeUfVB3gMpRVIwqjORHgJhjokpAQ0TRwKsreb0bMpSg
AsoUbf4k29ak79cUkUtgHC0bGbVAQpq6a7FNvrnBAmRjvC47tT3kvneDqo6AGYBN
YKIe9H8EeuU20Is2WqUzt7NexLrn0wF9yV7rkQSu/eg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
LkCbG5mEtgoKPqTN9gF7xNStYexpwNZAlLMvSLumzKCyNfLJ/xvL1cmnRPfEc8yb
lBgqaTkUPaiQQ1WqdE/grCWCv9NDBrtSgh/kNu8dSD1LuoU3lDit2PgkrBdBfM6H
g0WU9Oxi76O6jGxqat0nk1IL8fo/VAxY/oN0uWC5JDZtjJOCuZHHn7op5EHhcGr1
kRMry0/SAK+FNo9F20GUnTABGKCdrx36UQ/w43EntFd1Fg8edQcveNesntrH7w/m
ekpMiZVFJ+65hoqlARfaIgj8/ZczhGpRM9q7Rlf3nfmh5R8jmWhazohocz+m52Ca
deG+kztIsb4sTaMZqlXOhQT8uNmMGsO8i2jyDAz6Bd0iQ/CpIBon19K/ZIyI+euG
zBpqKuT59kHYtNrSFpdGiOnlRt0f2jbAlWEbP+Oj/DkEqDALR+Q0FjcsOsjAEyFI
mToDiV5dLzJc/1RG1V/wapmgI9fCYzM4PQNn6oPRJGS/TPKEs3Myn7LtwGoi1bKU
cAsAKlXaMAo6brBxU+kqsvkN1rwXltX/7MtymSW9ZBFFIjqSNXaPK6uCuaQLL+e7
XGZPm/zXQuPUv32j9EURQW9/A68YOwqVFp0aSym0oQ3yGytwC1/rwoU9KEZUaE7S
UKDC1a/c5JqMFohN8aju5Rdd7A8MTkCb+PYmTR7Y78M36Z7EatKr85UiZUNNBwPo
3fWQVAfSA6pz2bMdLFo9R0BUR1+LC4/sBpYUmvRQiQu0uKHRn2FhhJHtbGgTDBBL
mIBW3Ya67AyB0jHK3cc/yL6sBT1rNYPcQk2HZPtVGSqIZqR/JrAnzmvRdXVHwYP9
o3Ual6v4LVrbHszT35uTdXdqkQYRYrLARboZ2ECNVRZHQ4e/6EffwD7a0HS5QWXd
K7XkyBbq14PjWeuQURBAh6sC3z743kHfjOG+lRlR5fNct+bqNLTj8b7cKt46Gnyr
Q4SeNDQSWWQvRGr41JZX86Fqb5W03G7an1CDG+m8T4+T5tQxOMQ+/yPW1PID3ago
anm8KRRxBaQEw5Oa1tEsCL92YlX6rIyp9icQZ1Q0VqqmHA7qqBifC5tg9i1/kRA3
4vnhhGNbS3h5M//BRJsiTCB5BB6kH1+ibGCoSIkHRiXGdXrHBFHTmxUebrvOCJil
NBWCW/tDLo5GVx9bj5k3nmePAKdY1lTvKh1pczhzBN3ec0YjbZwg+eKu27Tdky3i
faDXQAd7G4j6LskByXBTA4O2CcBf+uIIqXr0VaRlA1TQm2B9oVh9rxwuYHIhxxaJ
g2seF6rNsg/r0t49U2DDBDQG/Eqm6inqA6r6EkATuLuJMXqjgwhl1Z0YHRtr54dv
UPZfhUtRz6RhPyi0zq077BAeVKvzUetmZS3erpFkswz56GklHcNHMLmHXd3RjI+K
rWvPFKfNhJ+8cBQgYlvnbZZVbK3Ak4z0stuffQzOtr0q+gcoZU2Oz4/OvYIy7xYT
3hpKeBLNIe+3jfW84r71YHHTs5e52qbeYigmr6F9wYPoiEN/cSOix85ALXVF8UHr
G6EPQZuqrnNuJiISwbDArA5+DWnFaPUZpd6rwilwif0xTaKzWF3I7ZpY5rjazAvp
FzMy/wdmgu5GN/gcifowcAGK33w2XEb9yNqzqsZDlnJTTS19wcryFqU2BWQmOxnr
UuqnIPA48cmRjDe3keKiVo14/2tBf9F64lvByvZuFin8KWZyeu/mW9z67Sy86Fpc
aA687VGJ/b6lZOaXQLXiYy6TtM9mGSuaC+JHLYZhaGad6FWeysYnOFKmN42c8OPh
cjkhzYx5eXeYs3NrjjzJDiNAEQKLcgjAHt9pmzzZEpT9RZ4cm+5kUTe1um/xbFUk
yO/DNY02o+QlPRIhOeaJk5nscOgC6OlUmM39k9sD1YPNLgJQ+CE4anL1saILa4m1
WpP9EGdXDFmzPujnUPMAqZ35EmCcs1hP7sFR6n5jKeW0s3rXvF6uJbaGf/vPyQYb
vI1lurDNLh26rLCZob8Ys1beD4bTetKsFlhSjwCzz70+OVGW4LUteY9sCRJDPklh
Mhnebrt8h2IzBxeHbN/hNBv58yT4Oi8+mCVS+V/6QjzhG0BNizzt7zBLd/R5tOKi
pdGbWyBJhNcNpASJDH4uX5bYWsrFMrXcuNeWfnhBGdYrHoa7gYZu9RIsXjpqJ8p1
lWZe9Ys9vUqJra3XWnf3tsaL+EGDwjJlXnRU/0WYbiYn7WRaFWhwZ6VTvQAaVZUm
y78JElsnyqhkrEbdIMqyAIzsvDVCSEWFnqYkkiBfPXZnbSzGe3W1WLQjFY6NxvbK
i70zbuTn2Ry6hLmLac7Zmg+KcLAoQoZxCxp2F7h1QMzv8bx5Ho/X6tqtRCPTVkLk
sKAYLgr1K4kT2GOG4ZzvmpojTY+PKzYL6Lg23GwWb0fAIJEf+/T7LCQEDGSPAmQ2
JOTHgK02TYrZ17BumeWJSDSQfqSgVwAujlxx+CIF6gysaezMv0wxdMWwB/RM42jf
JMm0FyQ+NiNkA5I4seS3jzMj8Hf8A9R4Yu0q7s4EpEfV6cslxPNxj+yjWA9T9hXi
2Vfuw9vdKkRev+FZQkCrPKZn8fV7prX9H2wMKZEChh1aO3rlujr0A5MTk46rJMY9
cHBqR1LBgOIBXOcOOsX4c1+IVlMmuGHbd9h3+IzmgAIJVikD5VXkmXox82FFujMr
gj7e8ZannLOGqRyTQVkLMUTOJfFeP0qaEWBZ3vzkP3M4G2vnXZTR4qp8C4kR+Dhp
OiZVTkz8l7Qt7JAc5ilTydpPnZm82Klm395PsSBvFwEE+n48PFz/6GCvD2dagVZ4
Ptmyi0sFXieuhIL538MFMavCEXoxv6kqwV+1ygR7bNcFpd+jkc9qhGtUCqQIihlI
ZfQzQUNgJ7rCAMrCixHYIbwDlg5AovrqxLIxRWAqSlII1X3xTXLqDumCxEdKEmCm
8P1FT3WFRxqmsBblqA+A8zk9gzZIjQpJs7w4qdY4YIRZh46ABNFJYfVPYQ8I2z/E
ItagU9n6KM024fB8q7ADk4wCNEwKtx0AMWvECvGX21Cy9etiNaeaOoqAqBywpS0j
ewKuNSIzRfDg5KkzJOzoaVuuccoyeMD9XYC3xkitD7p7xBUtqSTPQHPGpX1JD/+T
kyOQegNUUwYyGkeKgMRnXX4u1oS6YKzIzb7HQgNlU4pN8NizxW5uod4QsXGICtQb
Q+PV0IlBZhZaT1B7momR40BiA0Y33nO2QxfkSOMpbqTlpBfv3j3HJQIVPgifQ/aW
6bMr78b5uKBu9l3UgifimlTloOEoEhY517IqtNYD5IRX3Tgsa4xgKCQ4kCrlRDnb
O6ikuyqTAG12xGXz2gCA052uyKp2BV4/dnrblahMZcA6oLbNm92CKZwA4qFwvZkZ
YjJ0KCBfhRVMen4SGEtEyZlo8/+GiwXKyZSLlx9RjQsbzIEhoTqUDS7ZtM7JJgLM
ckHAE+QcKP1996IgYpK0oNPhs3pbnMgvlmzofGwZDt3obSWRcRdbv9RIVZQAfgXt
yJcVOR6UZ7KUKpupCWXOmRkEZuJL763blR6/PyQkjLLEZ0jdCKvfAluA2m07GO4+
twSLoQ+KOC/xxEwhdfWWBcYyLKgcLRvc3ucfjWg1Di3mK83twPpo/kieh2VDsdix
1efZn7bUpKJD3uQ77Iy1jXhToGmS3X+77vnKbA20YTajrjGu7QAzu1LUjYG1S1/q
jCenzBXsUPN1Zwj9guAuYP+bo1lsjEbKQpZatkqMdWFW/C5YGSVtgJ2TvaRo4UG3
tBT/Ti4vNF7MwQRJHUqWlN7P3wwbayJWlTEY2wj6NapXu5KejOHW0dyKbNMTASTN
0Ixc5iVtJamQrYkfI+GKr+yPkAHu41/NxD1ik9FIs853YSsfIz8Mr0F3l947Z3CK
gL17+cVQh8ulWFnkwxe1+ddsE9IcpqLemAb9/IIcAVErhEnJuWQHDYB5G6pG6W+y
vKnx8SNb6g+yKzteyLDo8oW098MFP6/vAo2Wg7A5i+t18QrBO5tQF/OYjnpr2/Rb
pDuyBEldyoQPWThVldYQ9N7H16g7H+jel8s9UwaalcoAQS0kO/mWYz6qAaFSxFpL
sg+LZvx640Qax355FBVvNYbZ55b0s27HkreykWrA5qROu8JLvWdaL1YL2kwNVxEs
Jooi0Yvx415AH9wnehnqVfRZHFXOqxqaFnWPY+msoLM/rJcNqNTc9NHeonfeghXB
E+uHhQqz2ZI5qb+k1C7bF6DD8yu7gK/T0XEgz61qqyfZ8Bx5Hoiyx066Wtbggg2Z
74OGEwOw8cwBJjtbGExMkWSm7MXOZfnxOHqUdsLCFHOUY/NvLUMffYOZBn6aRH6K
dEhEx5Ywp4VpQC94IJp2qFYAHXQJgQTmsefIbz5PQKSikUJ/xTuMFTKXqaDrP3wy
ZL6O/c9EIHO889qRE+QP6Rn8Url/UF0a8MFdDF2oOUAm4wJsMRFK7YZpUo9W6Y0J
PPZ1W2rRyuKqsgbZTCMfQq3dPT2iogu9Towd6TAOLIDhNl9SRrNIfF/tWoiHo4nP
tZ41DOx9jdBFDEAGU56I0ZJsyt8rjz41bRow2zqzCA0vwr6w+NtbKNYnkt3MyZWe
wKOBYuQamExq8MgorhgnFKZJ4YEi2/kcg/65kYbcYeUswhSS3MTtgpkrMkbeCqxj
2da8km4kHV92z511p2czbjynRt2rWqY6iJ4gVSECz8lC15K3Iioc60HPis40U8aB
+2u+g/5YBTbEnpJdamuqjnxeANH/jaQOlPcmaD8gGP83MCc2zkiUzUPcndKTirHN
0+MpXeCFRSJ+bnmiHFYE6QLQLvYJl5mXD6J/OsR1ev/zm/V7zgnYUtpa54+oqNEa
A+X9/bhaJvhQdR+YUCopEVphi1oNGo1+/ZREPENYNmNtDGAQyMiI/sCHSo9UsUXz
IzKfp1lGv0Wlq9uGd/XHz9ssi8Ej+lXZ4wPkUg1/X6N5gSdkcOaDSVDdFsCVLT6p
agJkdp1tBLbDeUkPCLFkG4zTcyMbReqx0GFv+LpKjZF675s4If91/X+4/8Qwcvq7
8lDcvb+qh7TOCX8dhFVJ9vNASSAS2XelsR9SswbC39GD1RFVfEMm0HtfqXJbXEoN
Db/03qHvUlrUyO5ykfKLDjxYgK/YPqmOydgRtRhsgIGLr16X0sOSkR1hMHAzqx8q
U5amMybl3rDPiR2NX4tL8CK+eXkTnAs+TcxkuZVN+x58IQlBdmIY2EhGxdt3Dp6I
LO9Yqe//tLpif34hXMffT6Wna58pa88EioGUdATGo4RwNcGqg2URb7gIJpzBL/pb
8TaHQ/uqjdG7gY8iZoLT4gK/pVI2lMVVHBGxcWUEqVVZV15FSerkmEivWn7FWoVp
ITnXEHm/+h0dzmp4Gk07a3QLv/fV0ON2VyC1mMCGwjh+tVJFnjHMy+vvtxYxFZq/
dGF5G5k4s7i0d/P/CQMS1JJxvTMvj3uXCnVnlOOlI7zwJJrU87SSEukHwct2QHP9
4GTrYg3eDUYNg9YIZ+aO6L1Xauv67uWHY3kCtfwTDjPbV3fyfwr2MItslLwD4zgD
Nscz6m5/zaVRkQnWifl3/t1W+OPDh1nmeSBesOi2rfrbK6npdUyUIKfNB5yOYTOS
z7qToLJ8YO5l2U4+dPdjGj6y3/Ex8xAf4kuKKQzo4KJpkkJPBmP5unowXg67dnx5
iGtCNVRkXELvxuhAnyFir75Fo4BHCJm8vbOVf51mtRTyOL/S1sjse9mxG0dPoZ3C
YCX/GJRSUd6nCZetkDxDZ/dhmb/HWvjD6imtdsiPyQvjtWJ71zPkGYU6yQVOaQPO
HkGmWTNtA50nde/R6tinKwIr9ikqwl/kMKQizQLcdfNpCJWS7VjFHjs1g1Dtyoog
xLhm+5M+gppQeUaNQG46sL+YdwcZ1pH10pWlwE5KXzPNRl9YT4OSERzWzUdQ1dJR
D3nt8+svagpx3B3B0NiUAjehjPuj3fkPazsUOzfTHIzfjxP94mKgwP6IjJO49B0U
M3oZQpnGGej3CN7bVSKWh/IRNzsHtCqLIiYNcFcuYpd3QdHq55dtrG7CMyj++JF5
VZFNLsmTAv6K7zFTnd2flBn+gOnx5bgWDrSSRnuiFqo0ZkQ8407iQ4GNk4J8mXY0
kAf9YL2I21tLpGp6T45Jp+LX0+uCOtaKzW2UsCFFw6wc0LFbVOX4jNxUwJk9j833
uLkLVQ+Szx/Bjn2bTE2D2CH4o8DRgpU+4dRGjgc/vx+N6Iazp3lxbuMASNW5S/IZ
6bTp0hkyYOTGorcQ4nZ8aS9RCyC+AhxRS/Oss+PCf4Ca+LPpMRFmDz1NBJZ8CBRt
W0HoXE9qcs17fZqG9VNQlmI1+PnZv01+MUcMAsubN13locbgOHIfG+f9NFKgShDo
kbNGzkLbSASsiBwIN+CSOj1zq3l73Haf3hbsS5hI6aC1IfviMglHitfAMtuBWLUv
zJvNSsTF8y8RVcDsYcy3IZON04N26xnt1ibY8ltkwgnz1gMilmNzj+XsvRsA3EJH
oZ003HwxFo5Ncj2UQwVjhaG8rLcgp3CRiVDu0H41TMiJCI9Q8T3JQWlIZsEiQ4rW
WHNdnYVtDe9hQAVTPKI8+dQb9Q6ivYrTZsb5prAM8bB7+gMKoVTqI19aIQOMnMA5
wRK2X8q3g3mV+pq6nuxrEGgpQlH+xXAaUJMr1ECsmm6S5jbZHswx8+XuJSakt9Fy
VHhelOMdhKsQnabzCO3iO0WHgU/9nFTWGMbmZAWTihBINYToh4mIiJDZ1yxHOFPZ
QGjnx7x9pSC+tBxfaw3XApAcGsRClSfD4wnhg54UxoNro/IUHrNk6/tZr0XjQaQF
Ykyo+22aVzRjOrTgIlMtllx53+m9k5EYZ0ZJADINSCqbyTgRQv53S/pbTodMFM49
F4BYOOaZcnZJEzn3I2M8kystrvs/0fauVCschaIs0KvqSFcUSWbFlwV0p2mwSCE8
Ze0UuBqGBEPzO4jOODL3CkPXBIViMmhHH8jtuHTsaMIuYmNM+YhjKyzYhFwLoCYB
wkHFQgSETxDOtGPAZOliCHoQr6skiCfLGe6nzZ76ZWzBErUYBuCXnFRrobQ04Qkp
VVJpnRI1cJtylVUNrOd/nHYd5nL2JehiSzdXuHMvj7OkSUswqondyeVBB5N57d9P
nN8oYC7G0s7T5xHcsYDZ+y3akWGe5fN5ehvawlaqbDgaAEHCa0bvisvqGXfcvAb5
7gsbfBDJrBUQ5Swv1XbNtIaI/Qe1z1RPNsJH5cleMAZ2PUlcomQkmrw8i3DYRaNO
0lAVjGZwE2AVLH/t/zomMdrvvqyfznJWckgJNvFnlRnsnZQk42emznBzeHzpfMvs
LgebnwKTOCH8REHI3PZvNOqfwFeCSyGJ+TdrVxSN0JsYVFi9r5AJpVnfcxCKCnV5
8Ln2iL1ChqqDbRHM5AC8Wp+rbvkQJeXUtmvwxonWtEV2ZW+RkcOq3CkIjJRHMXzy
UCw68yZuELeGyUXIoAje/o93Tac0ehl8vcur9qfIuR1gpYYiajycYK67ExH5Cz1O
DxruMHj5dfhco+wEyS3fHN+XIvmIT2gGWHKPnXYlHh3LS8aDNQWCnwOv7ndalfH7
wPY+XWeH4CY/FGdombIki3T15MV60X2Ss8TsM+9gNgbl+fsnI8iZpIrKrOf3laF9
wJCnhiNFnfznw+Nw9aDREfxgx/LGE/5QPBYGaZ5kJ3n2sfC73lv7kymIndrv+3WZ
PE0SNL1C5uwYKvEew9phx6is8FiMqmzgh9R1v7LGxWQ=
`pragma protect end_protected
