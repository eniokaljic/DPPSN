// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L6nmlniYhi/22jQRXuNQztn9VmWOxpHIm08ry0/MWkciSjTFNvXh4QdiCBu5AJ+3
G4YYrjW5MCHKK7VjFzLfKAQCHUU+bUvbjlGCZyg/i4tb4Y6/EvsoTAMaklU+F1Uz
aJaasru2NG4EgAEDORQ5grKzJBO/3TAUxkr0GYmdYmg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
GwwmyNZVjZ8GdLl/zOhedLeJpNGreuRjAY8dx10bfPPEcLr7exYmGPba83bE6WPK
HW4/rF06kz4Wk3RewTc37BxRsj80pFclGTQqZGzJuqOEuGMvWPv7VfwzIZuCBFWM
QNH8T/HtEY+WTmuUqFsRTcg98i7j8zyx/mY6ff2KJN7IpYKpiWvOPOOk4ZArB6ZO
LEn+n+JfMsa+4chiHim/oVIgGNeAiF088L4UyTtIJWNUKIrW9BsqI+yGDwpC3E5o
c5TpC00fFzrRKw8UMXBB4r2kkmHK4Yq++XKuCljLJf+PDx4LSqOk0+xfK/fvlYmi
nobbXE7gDCJbyPKSYdksID6Rp5UtJHOyYKMA7iwQzd64P8xb+PXAAQdFcaIFtifX
wsTD8r+3noAxKU3a4rJgBNH8Sx2uXJZGPxUe6ukWfh2wQB2uEpZxWI3SqugIVwuW
8bIgHFkbkFNCr1X/7O8117qMOYfUNd/cOeRVpVYA6KRKjF+Ikk7n13pPNW0jgZHK
ny9QiqQ97Gx9YwdCqX05xG59woI5pzg9Bta/npFoc4d+iwMDxbDTHNqOfzYAH2d7
dCsgkK+BntKOV7hQqfQjI9zWc7qXWZ7y/cqpE7snYvAVrBdnQ7rlyIizz+4lnkqF
93rcH/1hHgelBd4FOzGYeDR2LU2abbLP+sorvji8mrGhQyP9ws8YBvQamVjpaWN3
FBGG6LM2yAX/ps7xmfzjjWQN3dhr/ojjWFVG3HTfADETuLLFVpVEtb4Hfvm+W+WX
BWRQsz5kEcJh6FSC4RgNizC+kodCwG8syGU4OYdU8pSNJwHNzrfX6reXHnuom9bw
PanJLL5S2XF9ZVxsjHMPB79JVQoHwoIWPWLgtEQ1d+rIUdjk8kDTRbXlOnOPr3QL
o4TjaZPQrIk6YiO/3agiyrMBy1alIEwcaq7bnqshzwcx4uttUuSIdJOWMeBBwlt1
h+T5DnInU5/geV+xjSuQ1cIcFqkBDM9M4N8CK4HNeubYZLKDS0rwsJdhJ5NJUMaA
9oxf4wezHRxkGfJDz3XTLTy1tk/s7/ayABr3fhHTcwVEQEHwWaBDGsriQyUj3jSZ
FYPqYOrkkkqsPeMqDiAs4UeZD37Qhge3ZqdhF4Za7lF09b5DsBCFEugZiAgl4wws
glHggq1fbHCpdVYXPS+3iW1pIuBRwCeDmpdP4znd5PZPcYTbvqghVCdPyKJNUdEk
B2Tun0Kqw1RGxsq7GNQbsFmgMdwcosx62jVIgDgu2GhAdyONZhKP/jkPvo7NJc8Q
eD1dMndKQIzhHP6Khpi0rQVdvfRmwiQc6dRBlReZWtkZ23vhhJYaAxUL/uEEUU5N
nMNFfrP6c5IJKJKuFSS8mTIT91Qk+AeMhuTsBoQyQJQLOUQmYOcJBLjGHuEIpIic
4777inmRTcr5orzY79dK0mPBPmXKixhfIzHOmnQmU+MhpHzmFwOPfAHIgcbjT/x4
Ul2ECZMtZ0yJXa+xKowstvVAMdWQftQbbDBpIFPGS+QwUrGEp6B8MIBrQ0ReNyWt
8IQXpfYTC5Yg2LpOQCWPdyZGAeFgmgEqeOetAwtVftccvYYELMK6rlZz1reoCDNp
kaLeT58+9hp0BXsd8BcrJvSf1OX4K5DNlY0MKtq2ydxFX7/kAdgmbDvAiYrODFvF
NI+CKQ2qHq0GGOSe7wjwTnXUlpt9VN7BQiddiVrwwnWGc9F8PSv7FSqNv/Lo50S+
kz4ipu6PYQZZm3Ew9ALXoVbtwGYhTvprLwMv5peqvpS1/C5FJN3jWJ5YBV/bqMZO
zGURwxAjMEl1x7WmPTkXrGZla6Kcf07C2sgrn069873fYaPXe7Xz8ra35eqhZ+2H
ylZx4bwRAW/p/pVcG7G1/vY9sUBVBud3jWhASiZHkMVYMCI6Ee5mNRv5CwjCBvz/
PB0w+sHoQdrBiWuNTnQyw+POiMPCjCp9KthltkMXA+jRjvdeHqOjUaOesVSGbvIo
GRoa8C+MSVTnZ0ASsRJZvwzModn+mwEutcxv13UhP9cARj0Le5xwnZqBC4+xm284
i1g43oxMYysiSdSMCZlohikjxcKbuaAQyudEraAa5ZSGuAwEsFM3YmNdPAGy6/s5
4w0fZFbPr/CYjvnw19RfQCQYmgb8BIrnGaEwso/ARxS8Pt9Nypyyu4N8oNBwS7n1
iV52lerbucA04yFoGUrFCUaDw3AejiH87zI4EkLqHtGiqBEXN5YoacgP33EAmYp/
hV5lJZ1MuYy7ZV9xSpOceLD+/S2bnqNpIjzde7fCr3eWZqR5cg26MRWRT0mMCwPW
PVja1i44zW//oP0hkQKKFNGmHRTeFy34OECVhfKYbAUa1xAsi9iE/uWo8LgQHoCM
1Q/WeIPTMDupMsYjwH66xE5UhfjZBQFyFvf62sMYyZIqyUvV+wx/9HgA21j6Y9dp
vleaW0pJAR0QCzGgkPgSNlKa2+rG1klk8HG5bKt/0qzu9FBKpsbim78cQwSCI5jq
yK1xvD9JXVbAZkhDV6cnSh+vZIrXEXjR8tLon6b3Z0c19s5O0rHgiSTxbdGPnKfe
5Rq9ZkJTzZ3q9Nm5KD0nBQ2frdeYBFDdnvxUAqVbuS7H29szf5K11PkCR6A79fBJ
J66X0ES3T2p5CcXfEYCgUZKyyirSkB+i+H4YPntuN/vMZjZQ5IYdMWsLVx8kvdu5
oD/dBN4Iuephb56deJ8HWEB2CzTKgaOd+v2rE/DMMm4gNyoSvA5AjV2CMl06T35K
X66TGbnd59KxX9uOcmLkHQ470FgZWTSOkQeEbcckVEPSBlem/bsFwy2c5ToT4GHi
R6ZISVDSm1ToLebTRz9ddYqnDha3wsIiaxSaXflfcVAHSlSufQROk9S70IOEkS9B
HU0n8LmKdXi/wS96hq+efGAZHDkV5YCWVqRVmoh5hV6OmHIMRoXx/iUQ8hRtq0Ov
Jurn8Z1gAwZY6OOAVJv7TKnKOTXfWb8I0m33pCZzb5DsjYWvRrx6DXpdsmInkVCx
kYpqWJuMHHzm8qZRV1sM68ZsFnl/Pol/CPmdZQ2BExzcgP5jEmpOYfOrtPn9ytpM
sv2JeTp3iVwXbJ+jh+cbq0ZKeVQ9hY0n11Sbuk5dizjE/RX27GEPPBzeBbPXss8u
93ldOJ1nR9uNTZHXrDqU7pXFh4e9ZWGWfvuPXT7jNWaTHcHEcU5bn5dFPGe+RAd1
DotMgsuQAV5h7cjh75kFBrz1JwYsIOperLBqcfKlsv91/7Salzrpodr+jbE1OKac
3tQ/f0/76gjuxG5TTOhgmVBED0vW72y75Wzuh49IX5NHyB9RhgZPrKBtw4z7kOsK
9Q9aXeuAaPOl3MGxPGQNArAKff8/nj/SS+liAwVVNgib9mSA/8JdCy74Wx4kAWhx
Zd9otcP9kuzxG4IgQKF+EYgtWS3O8VWPQv/zOI+sLQ7z+suIsFB7oQngoDSKH6a/
cewzCTLggCsVfICLw+AZLkMHj58ytZyz00NjcSaiqY8m9EbGpsGqS4Kew8ykOd/k
nXuwZ1mwiEK9+sCpPNh+QIbbbRQCtnxbfV0a+/0TkqujBXCUECc2qCuf6yfTHM58
6CJePr+Jn5aeHNk8gkvjWyt3RfcV4jX5PLLz/obNN1UYSZlwo9g6sEnq8OsA2WCP
QZmoYesdcBFvtqXXuNQZ0+x6piRIHHD/gX72YyjeBY/DedvbUTicuqjF231DumTT
DRyl1liCRJveG3UgFqALNQoeamwy3LlkEYC+BFZrdsohXOkMiKC2rnfwxu62ryUs
UV/YSTAbYwjhnItCSlBpSfISkToG+xeYoXI8Z+zP7nbfkmi32F5Lb00LBE31IRg/
/1MDKwrQtDIcky8IT+KLajTX2U59RDqkF5togT3Y6EJ1OaH29jfxLsvvWQ1hIi2e
1A3ibX/2xzIwE4GylXUNDa5IEson1981wZQyIU/eqRCkUmt7t6ZmKKIzjbA05xBu
ZP2JVSrCq8sqbeHUtPx+rd11rpBoBCPhLT28XfwKLv/a3Z9T+WzCyqqOew3YqXG4
zSncpyskAuOFZYrxwmv5Su+xj5YLD63+JJN/QkOeG5P+Lj7c/LdvWgVmC3vjUguM
wxgWRC16H6fDMfCqaNvA7MfMI8SSN6g99szZnX7UJNRc6TVIIebpClMBAgFBDcKd
5uVzRjFLiTrs0uSev9wpMjsRvIFkrkqMOkYqJ1lm2lbah2L1MJ+mk3dGAWA/wBmk
PgO3O5Eu9sqGIx4pP942XpvFtJhz9EVed5rRIYfTcwdsPb1L5AdKmKLEGy7eLdiT
lbFzzZiScnlIqUVOmI9/qXwGx1wxikGGtfN1M8p6bT09gUOi1JGPf0iBdmcol4i2
UeM/OX+HLnvjS3bDBOu0SoH5pKMnAwVsdjhDFp1VG4SpwqzAxgeWU2z+CaoWD9Wd
Ock72g6T7uYIJ2Kyy8YyLheEI8GM1xT9jxsWE9K+E70HqdF4/HB9U1c8c/kcQZFJ
hcAUW2Dh02XFi7hQE/bq9fUtM84DdnysKvus8JmRMHJleEwuKpu3j/jtKuMJD2zc
9/NVARQPzDeGJ3jBK+nBRvsWo6JrXgi2r+aF5maFcSQSvEd0sTuqh/b57ubnbxSR
LzaTRw7aiUm5wfYrd5rJWilL+X3epRWOg4Rvl/tJxmHFVlByKThLonpSt0FP4iM7
b+u5gwrN5rGEadRj+L4NdDOMMAVgdndfFziNEIMWJXL9TzFELS/tPeVgjoj9i5eY
knxWmsSqR5af7MdtDRnFCn8x9mo9N3JTm6AhgfottE/yrNgsU8QPSAgxgBbJD1gP
PF1PB/EMQKDRYBuE7aD+sDS8j4pDRm/PtJXutWsIyDQcYj+tdMZl7PyRaWJitIJj
aRsOlpGXED96/ay9Sn8yqxvVOdUSqIIFreDkJIwIhXfXFLIxUehryGgvMepV4iMy
6j53OepxayNfJFHhBbWTYV0FjR1CbkqtRHS8NT9bx8HKRT3dEf4PUawKf4fkmM7Q
5wLYOio4OK3xJJvv+Fuiojo5m395eipaUBmC97uFse+muVxKMo89JQWtIiqG/Oof
cm4g441rR0U4Zwe2STa3XTIJDJznUbwJIDWO4I1CwlDEValA0Rd1kzK8sGc1s8gA
N3yHcTu63GGNXeQt4gM56lZM8PwY1FZUDF42sVB8X3VaSSDFF0qy53VNDfyGDg2W
lCgX3UNesP7y5vnzExUvYuOYT0tUrY6Vyu1f6hwOh/EajY4oVi4jCJzBJksdqq+G
hePuJpffg6iY+8vY+niOUKyM4Iyo6mE8gzOTM9SKxUqIEJ6968ftz/p9YWIsfpGV
t7uvQTq5jh4Bt/B7XhwrZDeemTNo9e4V3IP+LQlwytJJglTJXoSVgGF0J95L3NWr
Ra3ULphE7VMYHO8np4TMTS+1MHVYZBl+YNxRAUmesA2cnuAXIhyzUbYOFl5Y6tPs
RPKT2aQn+qvByXs/91gfFsOuTtt7mJHbu/GYcFqNx1qiDDlS5Fg7e1LVzOZDamp+
rTFtdR0zgDWqbUYd3Zvmf0OeiI08KoMjHzql1AH7QMYnKONFz3zcpXi3HWdLmqWB
BNEZEHEFyxgZmE4E6NXintJZt9OJW8FOm/UBMvGtVf+oVV258Tx1MXyIJsdXhLEr
lCx1qrxciPCq7WYEOQpK6zNUZjSUa9J/9v1qAt91IZPg1h7qUWuT8IIGN+dc8B5x
vBHJbYcDDZa9Ngmvr/mbkGraxWtFMx7xRQv96b1Jj4M8IxPBPQ0dKlJYqXLiLFfM
NO6/8DGR81DGMr9jFuYLDGVEKmx10cL3pDMERe6ZrlWviFL2Ew5jEN6zsUX9OAtR
stMwQbNaYiDeyNSVJee6RAh9jbGFYXhm07eEuG6a0dRTzD8HhfyPc5BC2O7Apfwk
7oYAuVJxnKzTJoJ84QVDiKekoFP11meXEtZHNfL3djtWXkat9Ffq2xp6jWyNIUB2
g/GWEbrGU8Ca6RmWhsWUCIDxWY/ymG5cSXV47XyvgSWZ+RWVA321sscsAMyQihY8
Bj7um66fvyNzfBkWRxmWn99ZK7aHiRCYMBsj0eIm6nnWbbOyuWNLoGdAOafGubHQ
PXa4Nk8yUiHykn6szU9HR59KOZk/1JNAlNJAref0Cv5UfdfBLj5+PHCJMuni9LqK
+s1735bUfnOZ+KSu5hvfLQ5uNPGxDYJMeuEqVoMl9nfUvC7WwK29kmeUHDdtOi3C
FjcmbbAvCFpcKC5o7Kw9Err7mKBB3TAb4OIIMjKygzNOZfbrKDP+9PDD5B4tWmvc
TJ7bGvtgljg6RSyrgMB7wKo7r0vZdbOy3JncfeI8DXxZSJhe7ZGUl7FdnfIc/in1
gudbEH6g4R7xhfs9Jz2fNWJILWRDh8i2fogp9ZjEuyuPbcTHPhky+R/PNhq8kgQb
+rfKarmyA8QTV0dxKHPXtf+3eVejDCVB1H0eF3XOS0NoFs9X+YvEcmCBpoVnLgsp
7JiscksSmfVCJJ/uy9MRwWUhpzpowL0FMfX6sbQNcwLDm/20hE0c4mDgddyExxkD
S6M1aYAXBThbqSefUEXmw4VUZgSd0Kj6bANkESWOqGtp6aTUTDdYgAvqKD6IomHA
D8mRLiWh7cokwjIteJBpv82vxcmk/6dsJZeHPRCaDUz1SJ+2okGMQUdn7TIEjU4Q
5BK47Xr05plZjAq1e3fCUO6m6JzSJbK6u72zaO+MMaTeAPrRVVEjJfI4aX16G1Ys
xzYEYPz+oNM9MBSyVkUhMCb8K21f0bwok7DTnHYxEYDGO1Ydw+tzfAC0YRqyalof
qqxHEtkm5OR9U75Hf7xu/MRr3WtdLshsuCgYUxssyjQO5y6TidXHBKNv5PgpdENk
W75IrlYKHHe9xCDiuQK7qerBYX/CbT/QGVbGygeUubXzYW290cxWDE5KiPiqcA5D
c3ea9ic4FcPzjBCezL4JHKPTVsWsN1zr4XRpCW2SzYgXKsAzJeGo/2wfSf6/RmQZ
/aVYqi4akzPpDLkgcE1Nn9Js/rwku6J2xYhAOV+kIl/qY0n7q2ZqdkaAQRd5CSRE
Xh8qPnQm5s9QXXyHGyJYoBhzxkHSwBrjJOrA9P7R9ttnAVD0ulYJPbYUbpTs6o6b
ULKk4wgdlEuxjCCaH49HYENEa+Mo02da2uEPGJ+TtIT5xv6+eZr91UHvc/fMgfmo
esE5GKEPp5xGcvIJXj6h2wqeDGCHVM/INKnxcArtqIDx7k3seDZotxWrZm97a75I
o280XJfDX1ABCNqoZCjPvDcKtx5C+evg/5xYfJRrGBf9zZRRuu1pwFepMz2yknJ5
tGBcighV+SsfersXs7E7fQsqCFQ/UymDLGeX030X+dv68hjGmsyGVvNfU0D361bM
fhl/YcKIny/Rm6/y4p5pKq0j7rQcTjhvqmNak1WsHz8FzTqTPtjxL1bL7U78a5Vz
XNxAwdY1cK379YiuiKd2EIcJDAcUxbVcQEgPdXrNv/126ohUssTzPj1QNAf+XC8P
7F2OKc+kAfxg6Ny7s+A6YVHKZicIGYSmXEoUoHxfheMGNPyhdbHwITn9eU4UxfO1
1MWTSFbZf0qTCmGhjZZFmzW6hFK5fF93wiwaeFxa7l/0WAjWJXn2wYWYTvGSUG5z
MjdFnA4gZhfQ9Uy+XJ2j92eD2eTH3V9lKNMpWLxMjrLjnBGGHLNBfjGmdxp4EGpC
EMAs1hULXvA3Dz6SF//FBO1A1pd7xAOAsU9LemuhO99tYTcshOz2Px82nadMIbHP
3luoPML0lLV9oOA+ja5tQMTfLMUvezOf52xMOTY86AEu7gRLzY1exVXos4ggu9NM
KpxMneZ/+zSqYkoyUddtVDmYVg0ehDqgZ4cLVT453EVQLELXIxZL1ctzWzngzxu9
PMz/S2xwc0b6r2oH0WVSSxeLlGmvmx2zktqJ33e8BLsdoQ9zDP8yd33Ha1nzKDUj
68BYGdIcaj4oDwoccS3JFQEsunSpR2Av1MSRfZHzhbKym1Itc2oYZ4+tYHImrG9v
BSLgn+ef4n/b1ZnK4G7UFkl0kcpyiQIyMyiKWJZ3qm2Y/UJwoeFZ1S+uxVby5fiR
/dmuLpe2oQ1QGo4B09XbCHN8Et/fln+bLRNRVGLdDH6j1be1tDRAoaHqXozrkB2y
niji8Y/p8zKVWqgZvjuZYxDydWf64cUOF8kvaID+duh5bwKEG8J1QjLffrM2wmnA
PPkZsuqHO1un6hMrOTVB2kJDJFNOjBA/hHcl49ny1+8V54yLptF+tw5IWvBUNH6o
tCHMr+gaAxkNW+6yxH9GWu/+IPNS6W8f6vHhu0owxBYX6lod4kakbSwUVhEYu2L+
HetxxDwI4gHW7H4DICe/G9KFFtSddXmNhgeirG3VIXdCtz3Xvo8gezYtisjhJdDU
GEjsnd3EOWA7Zoa4aKxsip9FGjgsLxl9WRyahrsff/x3YIcFFHvOM7BeBPsXJyQP
WpEyB+w+0a5BRm7S4nTtj51A2sDzhorsCp9/gQCgv1a/UOeRDHadZH1rzqv9hPSe
sOseDJxQXQzNxljyXB5X/Y/W9JtZoG1+o29/eUFeA+yOMCGa6A4Of/L9E7bcRvvn
Pios13GelhU3gyLRs4YR4FCsqGMtOaEcj2+rE540JH7Cux4GQnNIJsE/sxB2PF2+
dIUCfi3ANHerWj0AJrl2ofuscfv2xNvjqzIxcys+Hs9poq5eR+WUY80jRT4SAI1K
jGf6PlBMEyxH0hlGg9AF/knE575i5l5LPmSfZ1pOHsp/PzgTFk5XIrcCGqC57IvA
6dC4lytYf8t/Uc8JNdCMI8wpLOxjzY6fH/UI1zQ28U89x39NrEGpgWmUmcw1Ufor
m2rwSATiVTF+ehWXs7N8lpmGOdcGOS68P7+VkN8aPmVpT6NqjFbFb+SgDdgInBd9
BGfOWZtgujbheZGKbycdXAceDb2dLG/2wkLx6Bz6770dv/XfRsNAOI95B3qIr/om
XDG/DihePG6dd7Ud1rY1KEPzDdx7mfjBlwnivU3zAd0BtmrC56+wnocw77P9bwvr
FyAkDsDf9ikkmbWNM2VJ2oSpqLPJsxaPhL1QTlhUYNTIOE8AZCMSQ8m0bqf6cTcz
/V5U+QAs2EUmPTdUXXd33JLVvoZuwCaeGhnTHTaEuGT/+RgLU6qc3DRGQl2ip/WF
kTBZ5jKPIbmXCfWkodXIKsl7/p+yXMdPjj7Ip42Uq80OYkjzlvbBWc3wVTUHQWmm
DxHH9y+/ZB1gOlCkiCZyvRC3Dc4hDmj99syoyW42oSTVJepN7k3skeHEZU5Oyvnt
hw16jh96lsPa/HoCuaCrb+A7DKPhOgc8RdVx/JxwgUk/gY+P7jZ95RVRXrMf4P/y
FGjGtwAixA1u/1xxf3sdG0dMxn1XneBjO6fee/G7ZvByD4mS85JlLI2kxx2fW21M
P3nT1M2spy914gjc6EDzw7FeRUWOgxcNQnPTqR0ws1UwjtU5bdW1UpNTkOYc0HJL
hZqcuFFulKo7xMWPPPeiA3P3c+d85gIQKF2bqhsvFEvAe28ktT5RqOh7JJTK1qqB
BaVfeSyvV4I5fGA/40ZQkS/4rUOh5KKrck1Jf7x4qv7LqjktIGoSj22Rii8AX519
ClD0pW0uEbB8Ij6MyAjCdIh37DZx2FHEcnP63oGR5G5kSoux2OtjDZSJ1h48Bs4w
bluYoPGC3BCpKRNgaN7xIjMz7FE+8qxt5eboBLI/PcTGF9F27IjMN/e/zumNDKkt
9+Pd/j9J4LD4m5UdgW433qYJ1BbmgRiUlgbqAnzWp4vgAUrVx/gkIArjm8b/y7MP
Pw9FbQfnzUOGZp1cB68vgcYV8PZ4WDYbwtVxumAm8O1NaQVb7gFCF1xfAmouSMPA
E+6/n6TKXYLbMkDIGx87q5GyLWVNV7dTSZGnlcpHZkeFCzuysMq/uFBkxhDcsC4D
Q5pNNEJQ+T68mfQrVOYM2m2saV/R8fXGT6gdCBXt1hHNZEDzN0RX8lBdm+Tpnw88
uf4u5HSVjRhZWNJlfps9VsyNDOCaaeVruBSPsUOYZUjElHDdEmuoSK0P2dD+AbYk
ZPvJcbJOCoz+p3hvO3rwp3SM32QKcP1gyoxOqJu8EFDocuWuoVxfKxAl3wU7Y4Vk
7MY7Xrz0Oss+e8hcO5j+6hmf8SWZQRliWWobY+fNd7niUQwDSTavxw5AKHcEQEib
UiHofm7KTxYtEWLvKazRVFJ1UzgMeU/9vBOIJPdDxKDKGrCNKC3aeC/fKex44Do6
lgssZwmnlWAHbWwioFG806NF+VuQdkz81n3FlN+KsDLZ8r9Tz4yuAyOPYHWTYX6g
K1xjCkpRKAGb0fa5Wa6DL46eCsxizdyqzTGiYLcUyS3V1RiL1K1A3aBWJnZQ5XvD
YYrB3S24qe52a7Q08V7bm/sF/6bjoOlxpZcdcxzZsmkhXMs0q/OcMuU0h7GFd6gn
oUCneAyXdZ9j0DPdCr1F0edCvhTD0tKuTN2V+Pbp/caz/E2YrROrZXtqi2XA9hCC
rsFphjTLOANMLKBJ3M3D7kWmwQnrjV8bX6TDh43+wIvUa3b/jS34xdqvYsiQrDNI
JNrtP3FL1IXzx2B/6ka2/UOjZ4EwRXM92eBedp7kZa3pVHn7X2kV8AEreDDRT/LF
ZsUgV/ELSRJebHnQD4rWcCDrhCoqEebJ2vtSbIH6r77kEOpV2zyH8273tF4TIQ54
aVHrStpDM338PkBRFXWWr66jXq9JxCqe5nkFa+fHYwnq3fmb+2HICCLxPZqHByZK
rDpz7Rb+oqnAs8/yc4p6yB9HvAZIIGibb6fm7hOca2IWbFN2odG2h1RNSlXfKW4x
tC6TQ0r30YY9XfudZvmOT7h+yKt3UIvf5xe88DmOEg6Z7g18RxEItTiUpL53VlIz
lstnvjsHAbyrddNgzFwpLHpXIMH2rpsXenKxfMUij4aBLIpHL7fv45D706T5R970
5JrbbH0NvHtm8K7I/tIverRskkqvo7FD+BkGVdw1xYRZg2iZ2yDY4/D/5DdN5pWg
Q1q2dip4Jbbb9p04i66iimDZdBb6o6d2DQ6oUR9zbPTba21Wp3sZQIWLMhZ5ZpTh
HTrGfnshnZJxjpY0AM05UlyfI1wAqbFd+9P/prNxWiwXph289E6bd1/ZB5GHOJme
37vJDtAeghUDq1Dz4tEI++eTbVMLSOBApClf8YyPluosOHjJs20fYW53yqvfnAof
VMK5kHS69dwtvY3oA3eaK2BAIp/TK1ALA8PWd19450BKLXE026rDXYy5ntw++bZc
7jiBUQZTh5ZM66Rs5XYJMSx5O/Xaijb5htBy0Io3BB9MT73lCkd8+cN64mFQAXx5
Eh2SFGWNchMqMrUxULMn2CX06ezkXLnG+EisQa8kn59inZTEQ9MZveeTDcTxDZBw
i7Rcbz4LKn1DTH29hiHp4oNU7gYOATwGu0j2V5hdiyf3Ror2uTnRM3ivaAzxry4X
vk6/1amGoa8/IkowNpYsFg9QBo77v8ZmlNOz2PGeb7LudVwOkLqUaCcxyF4wYv3Q
JybsJyLhKuMm955xvbn5wvFU8sGBYcEC2mRXkiO56nGKaevnYQaPJP+3oWXWXAu9
40yO0CIpzNMYxjYcY0Cl24hfZKCTYgR84oOFcZi98Pyc5xnnUEGbzt+yTda6MUh4
qE2TsnAZ6a4iVtJTDn6KRBppxBDCPCdLrtz1M9FpmchEcs/GgApcnAqyIokPduyN
/SpVBoJlahA1atTB5NndBDyt3QeRsa9LbMAm3CV4hbFAEDlYx7c/YvZmkfFuid7O
qywRGFcjq6qjREqO/tSRbdfrafuViVvR3Zvy8X1jttzFRKqYOFwKTLPsze+LduVf
zDTJ12dGqY2m70v3VxvOV3X0SJGvKVfgWD1XK7idliVquziHfMQHQCYRsfYJppFA
5TJhZKdMeb3e6QrW+UtyS4o8+m2AmjfCkiYuE5tZJg6fhJTrsG2qZb2q64FnOIRC
oFvotdUej904zPd1rlWLh6jR9mDduBcaHruNAUqkO4//xMBPev/tgpdd5pUpxj9m
1vj/pKPwmnus+E78RVuyfMtC3zTHmG8EVtbpet9SA/nC7zcIyVkNCGFkFbnEOY/z
XSsE9P0LvgrUzFGG6eFUM9yJlco44UzBvf7NV0lpwk6WmmVtiAkCqNJNVefjbFkH
yumLDHoQ3CEA3fl91kjRardgNjPXLGfM7UTNErdoLbNTQOfEMCJR4Wz5jj8KSCXa
3PiiPJ/OOur61t3MhN/47y0spf4Htp+EzWWmBZ0cSyLtEy2aeiNFT+SGb9Vxftrp
hwB9ktPzrKwt4j8pNc7pyWlYrK19aLf/EXggvlqJLo8Teda7v9YLaW/2rv9vvjKz
GaICgYnetJrgH+vSpX6lJ1brbfRQwkjyI/OFxYmhm/OmhIBoNK5EcMqmd4mYpVId
kBHNk7dIo95Hz1zPAcMujAy1hwWgIDiDYROCc65Zwl3qt3e92WefZtLYR5ixTwAP
5bLg6lTav5OzRSfsrRyXPFbFTW77VBwTpBivZFrhiWaqt5DsQk0OisgIDGksHFw0
TZU2CzihF/b2TjEVYlD5PAU4gO7bNuMu96rdtg0O14NJBoVhDOxOrYpfcZrQOdqi
het9UmA9MoYUGDyyVL7AZ2rIFVV/sPDDbojFYqf2+ZRtMmqsfinc8BYztNJwA8TI
hY6K1nq9uebxUCWYxlFQmBYXt0Vmi4Sb/4vcoAa86qv2PScLwieyDLTCJ7BmsAmp
GCRTuYHGm+2BpF+ZwswlfbaGaRtqdetkJq/t/9CKFtkKOiaxs+GfK5U75lbdm0Sf
5A/dypr/7UFSC+k4+6hA28AKtHLXM9/UpaXlbnlLzCcrVoo+cA6uYpBVaKXyOAua
GSZeQ7sUa6JUy0c/uSneBDL46p4QKN77nL4UMIbRjkG7AnA38whZSXitYgdy0Jur
M5LFyzyvILGuXon3/SQSBy34XggX7GQ41vGdZZsdoB0/Drk3+maH6MOUTIN11jMQ
uT2VeH9JDk5I5a1mWNqEalFoAulLMtwRfVMm67Q70sZu0n+asj+mCfhLbarH/vdF
kHiAr2jSyNd9q0vFpjewr9VM+3rNxIi+yhbKS6q8LBo+uy92DghQHu633BAHHs2Y
SJjsSyYfiEbhlDXflv8urv735aK7iEAU2fOyhx45mMRA91d5rKxp2waTTtEG/5gZ
emWaCFIfFwY9/0/e/ttbJkKXZFdBnBZl0g4vHk2008LUOk9v7P9xpWUcadCauydv
AZFixzwYgLgtN85x6SzE+Sdd/Q6wuOdB74pSDVqQC/+DLtuBlvuw2ShoTCBykoz+
kuLmlM9TNUnihf/Ia+8z3DIeDCX3aSLKSTB7U8cwGX1R1EoE0W2FZrfe8ivgwDl2
Ok1az6Aaev3NXdFlQ5qISEMm+ld6FTj/yOK1UDTHHdw8xXCt0P97ANghv9cVrBNB
ry6Bj6In66K6mINRD5sqZsNpXDzTzggL7X9qAlIHiz9Pdyz1wBqvthEaaFv3X3Lv
yfYT7FHZEwGvP2a5c9sOIGYO+1BSmtE6wykAM1semA5mRuy8PK1nhJaKM41fZ50P
9j1P/DjBQdTexHe2dYukvLih93MJTtmzdUCoJ+gQpXp/NhRIZxdSsaIneeUSwchG
+Yg94AtYwemthFnKX72x3ZqmkxRGfpP5/S1vhhTdqxKzbTkD3mUnXpLDD5yOb6sh
V3QO6QQ/UKFxKYL66K1y1+VbhykgJ5QowrIhyQCJgCZmTKu2BxI6a8Qlt0V0R7tA
iiiZHPsEHyGY9C/Tba2Rx/C/+bcUnbHQvHi/UZOlKgwatfP8vA1t+exR2gO1n3S9
l+CKW2CB0O9m2KztDD5iiCvygFsbRWWIrULFSmtx8pV0sbgcWi4BAaHkzBPOe8fJ
D43SLl3MaNF0Iu4vCHrrjBWBvr8O2FEtkg2CVw82GbzCPokxkaIsHJPZ2Qd2REA4
xhcJOBx8ycMs3xzexTh8CvfD0AXZ8j/xlUG2atD8284WpXwsI89MYCFjdGkFSe76
r9xuwx7+70x8PCKGhNM3rtZMDyWpH0BncRtl/E2qFKv+4tfn3pZmB1sE1iH3klCE
l3j3g+wX4vvAb0dHIahQdrGAF27lQcsZAj6WCnxZtcDA/H+JyARnWVQu2OaJ/ZSF
qvaeYBwpmkoK38wCvJjVzqd6dWkAA+cjWoTNNbek5sT4VEegBiSa8caQbHxvEDxk
QgzPtziZtbsCbLYshPJmUaWgtylJ/91BUs0OfoyLdm7iS4SRxooRqcrWqtIfjq+R
a/cM3QXm0qkGMo/tVTQ/n1bzMcXH1Nq7ituJpQBSJFPYlxW5ABTQQTUWWIDqLXd2
ftEHgsSpjxL2DZNxGZcA7V64MKru2QL6wLqhYxi5RoZE0R12Rmxs/1+kkGW3TcjA
sbWzwr7PHG+SVWbF8YNjZ9zjDv0jzBOuwyLkbkYWASclUxmlEbbj2NC0V2hgK1gC
WUImyii0lYXgYwX/iX7Rz1ZMLrqWRabr4UQ9hjInazIeQWqA6KgdKiLOs3M+KcLJ
f60b7nY8HKDHItowiLzXr8mhoSMA8K/B9eQUNCjCI7jCBWmuaZgYs2RaPZBDJTLG
pUP4Y/6JwEovxZXE/J3Kco6BqPo4O6HLGQC8FSshbj3vUBkjlzFs7P1YIMjry0aW
4kYspM2FwoGj+gICjlgwkErR7GCcl+do7DLRkIus+WryjxvLt7iRqu9JJINqUXVR
5ZJsrs8lSCUzaI7ho+QM7JT5DzoYt83UnVjIT1tEJPfnPz5Dlyiy3//ZartQ/ixa
gTyG+VjnmZbeYhIll3sU7jxNOxzoR6q7PSGZ5Ub1+EpkKfACZapczL0d8qdrQcPr
olcc4pB4VV9W+SE4Mbum+Bj93xdXIIosGcbxuoBUe5x5zD2pFwBDKQa7eB8Zzjuh
sk5RQcWauydeZdegxpjJEVHAXQiqTGodzgaWex3QsFsjj75U/dCoJvDCUeZJPOV5
4cJWTmp3ssTNwKDx2kuSvc47TWZr/guzWQhQPNe5yCQqCrINz6RBoqS2HO/hjrgZ
Adh8c4JVKizB/bFG6zVV1X2W7OdnInfG9GDKu0IT68jKAsQ8va+SSqKjpAFB5lbz
euBLymMdRLuSTDdepx+mhXZi5iN/sbbDOa65iTa7qy66AoNfoVZeVekeXgl2P8Ao
QiCn6LHAl74L96O1RO/Et/TDuAaY1C0FAhaKoQ6ukDNRno7f8IScrnJvcz9uEAbM
j0Xhrz/rOINvGfALgw1AjY3a70ApmN5dieRk6uxK0adAqgjqBnVaPtxGU/T9m4Ax
dQjjTmBeEfRwl40oKOX/qgKp3Ha+meInJZNAZXwN/dRQDIjr42kRW45VrBip4xsh
A4p0Grl26z5m/layUhj+F6sqyEahb8IUGyRJ9n4+3f5cVWPeMUU18B2h3sVj/Nj1
BF5njFNtQIpNNFRVy1mdS6knr4mFaZTcQhofhFWU9rVguiXZLTjRYv9THYMtQGK/
4k/8BPl8ee4Rayu5Sv0YeCZk9GhfjziQ8oJSt+jz+0FTat9ImQO+wBBaGbHkPvnB
xIXXqNueljjkmVuW+7geRJsI5/VBFjZdP496mOyyLRb5dY4oE0fNM5AGV5Ebj4I+
eXuA4PkgExE/xWztHo5wOrFdk8hqGnPuxj/J4qUP3nAHnlxWvtnfD/KrZXWF9x11
S+AvmRtD641oIRPOdIhk6srYJAvo1clXYVNOvc+xykAarQZ7Bwy2p8Y9hG1XQcJO
aH1/hwfjTXSBtMNgfmS6ql9ZA1OPCwP+104yVNhSGpPHm1QfBH++SzdFY+yAooV4
p54oxm/8imnccJRuRJbaU7VwJpy+XWZj2Y+NkkFARg7p0CYiOAR4vllnWxcSEqC3
QfebH7kfPkTtwdir09BVoTOiLTF9ez5wfxKOfuPftQCKE4XKVqhGDeYDXCopc9bL
Sw1pyt9NPFrVz1XdM/XnujUcdYev4KLVo0A62dE6fP0+ZJJIfJl0gzUyMR5v1vo6
EvEqUDubNus9lr0Ip3uGBHArnDcmqeTn3mfmVmVZVCFVoE6QoPjrTPCPk6gi/mcv
2NBDl/NZDoZQMmz83laGel29sE3/VpCmHdaCkZialHNJijvzx+f7R2OGoxaz7k1Y
uy58d0AT0gHOC7J7094RqwMhn6TWEIbJqW3NooekwwbNTl9jbhoRcO6bBf/Zu283
U74r2HLzlLLUmankFuzyiTZpRJoujowKI0db2Tnn1+F8ElAukr011eR48Sc8kYwW
oeOyyUyxf0xUxzR99X/T48bCMcd4TAfJFpAMHXh5QTHnIydToFOhRVQWEgs0qDRk
XJiwsYRILkWvx2IOrUjwT/a93o2HRbLqcaL/Pg3YXKYlNsugPl5fRMd4pewQyjRy
rYSdNXsUhOXE1WHl9KoUuomGnvYxfS2KoLDLCkuBlTusz3Ip5g/F5oXEQsbLjFHg
F5FAfxNpW1tHbUUIbb6mK+TGKmkID92v/XX8EIyWnPk3VDPbhu8459a77GNNF0Uv
25pLGLNJBc2kJV+x6En4sZXPEH7VlkUX3NHeB7aWLVs8uT7EZzPbjaS+PZGaREOx
XlyEm8aaVIzHw5Ovc1a8U08gWLy8+7FA9FB8XCaX7EdzLbu36v/cSCUv6g4i4nt3
+uKvMQjeyyxeDloMDfPhFcWB3mXF5R6k8xoUh/GvMrOIxT0gNSIOntFANy78hwZ/
8XuSUxl8vUGih5UFvqLqFu10d2H/1fQi7Fh1VS/mCGnlQzWOEvpw0ItdejMslpCj
3bsgTEmgIgAIlEqTIAkv8I1obLh+HulmaYc/bbZoeoXIUBfL0YMOLZoA94OGhYhX
4DgPzZDPYnryU8oHG0oSWgm9ECl6QEKF0Z42eUzu4LBM/1ehPevPXDCRxJtckfL6
m6AstV5clst173VoWQ5DMJKO27hbvWqUXOEl0smy4RSUg82RqJDv4Oy4t92ECsH+
FIx/ZIUNZTbEcV0cGPRb7gvYa+gWqqLNKezK8dXuv8oUjzc6UFpZqbFQdkcgHUrg
RvoR4b4R5dIrcZfSU7BV8PNWQcBCHYQxqUCFpm45pzTzfrsVEEp1N6sj+CNwMxYu
ktbTsO8cREgxbyanHI2jU9Ow+8BJKmqNapZdmCMnLlMJiuCxBHet7OHlG1XvRjZ6
/t7XMBoIjmzjStl6vfIZsYLWykOtmNaAgdhDuyXE6/V+/fX0WSCkfDSMiBJqg3aN
hDCem2ry98Hq/I+1vPVP7uT2jYSdzvQw5AJgbusv15PI9N3VcM1Jhhjqo8wpOitp
cmu7kL2YPl5GT84Fvv757nIcSdxX0wr91hiRByRT5vlyXpwFwggUTHmIwZ9CIBsR
GBTyojt+0035KGF6yOWh2SaM0XI48QEu4z0FGcyRrfz1IBdjmzDzzyJ5RuYgXO25
2rPhomGQ51nxocWyhesjQoU2xPnxW73/ZU9CqnG9JU/9bQMrWqfow2m+buzef+p4
t+mwclau89dEhUUfTIL7eLm7ZEXg70hXxk2B8zclliXYyrsfBC51rOo0tdQuQuHK
lsaP5tyDkSBD/c0os7EA5OdYWCwrw7gZGaHBOdU8k3ABn8B69AUiMyKwCdtB9okl
ID/0jrbpvSda0SmHmpUEBp6Ma6yaXGskSU+n0Q5ajMNvG6LYC+4xjz89BfZOe8kd
mmkLp/4sYFp1fTL3gXoi2yAsbjpQE7rGoH/l3EAoT5ioZD5xnWw5aCgDoWHcfy3O
bqtCAuF5gk/1IfpOTqZrHefr4HMhwYc0Yv9Tt6agOoI3f0/KJbSORondnSe08L5k
`pragma protect end_protected
