// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JJxQ4I8sBVq29SmWHufr6GULgXUytVmniMm0JqR+o0StkR8VDYIB7i1n4jF3YUCv
XyfkQOfzOCm7WY3eDzVVrNAOjRPV8xYUsz8nxkKObxJA2qV1Z++RkSUItHWk1zyn
r9sId3WFFaog9N6DaRbXrlToONKc7ZiQ0N5AAAK+GsU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28784)
5R983Jim8CWG9Q9PrQjxxmopS6UAA/WMjfaGO8iE9tS209lhmt6gmVCl8WJFb5DE
BWN+gVqtTjDgpmlPOdZiIu3750p19qaNBLVthTyI7LMPrGz1C92Y0Goa+SFwXFmk
UY+ljWDmF+2ygsQu9CK2Z7aMbrXIMk8FlMMJCEFEzRIdS7oXsyg/6R6qqdMvzM9p
kgcr/ACMAkU6r9YalzOLrO6EsX9Vv73V0LH8M57DvkX9LPELm2oG9ADUPROq6jTA
xeh7pydK+9+htGSKuDyAH2qkIE2hFxWHizsp0x/6gyb2odEl6SPp6bO+pbtRmHW/
9hjhStmsb8h0iB8Yii5sMDZPPAOJG4otttE7uEI/+KWMm89cqSYH7Gt2tBSX2q67
8qUEVtOAP/A+uEz/zSiQ7ZC+E9b5q9UBeQNxRbReecQonUxxRJIUynqh3FyVBZvh
aS2Ibrwtnd17J63J4N9a8UWq8xLTaw8wUog6fBEMIVCYJ5lfZvc8YmkIc77oVwXK
H7doBcBG+r6aCVzmuWF7k546KNXx6+aRBrNV7jni5XJZJt+pS3oj3iKmYx2ltnYH
bddj+vWskI5TfgWe1kniWwLGkAZoTp34RRKBRtrjFBFrR/4x9KH040nqVIPsTRFN
AupMrVhcBHCb38XEJDbiyja3xeoh+cfBxjHedWHjLb0lxT4MbFdqFZU3ndkoyJ3u
supTrHXYYnY56dVFVN5dlXJV1782+4mSYjMsuSofcCQMvvNvvU49XQyYdsQv3TXs
WemtCyKytTrow6jgZlwC2iANPEF1RW3ia7a4DPBHLXnWdqwcMTZxqGUX3RLHMpU7
O78TEiuW3lZCQdqJzeBQVHwgkRVRI7K+npxP5DgczLxBcnq8tDpgQ8pZVC4GhN52
jz5eN3qAYjSiJc9mw2zWANoYEI750WbuMo6MGQLuaGIw6CQVTCQAiSa/lvaTyllL
1c7ULB589PVPApAB2f4GGSdfQ+VVcWrJ8hE/mRhU4cWXLpLzsRkmvEue3vfiSqh3
9ttiGpmpcPgZJ93cdOP4PffQOd6YDbu4+OfKnnNqv324S7a451iXJD5s+kGakLXD
VFJihHNywmJYQ5Pd1gKKV4a2jqKvdmQ/UzUSXtYVhHrCtz9fuBAeq3zKJiRkFrEG
M7RwZNGVYS0ItrlII3t8m5Q+tGRGcjQ+eraWGfWjcRnWBNdkMMwGAu4Z7thQExFM
HMtta7gz/9t/T8J4V276ndlfQs3lBXrLTjlMQIhO9T05zf15NcwL27tfdlSD5B/a
1HJhFAHTXpEfzXdjaxhBWn9dE3+vYrQ/SCyZRfcyqbLFORzPvOLDH8uWMszp1k7l
oPxOzqKiYA5fCiudDSHETjgZIRyCoZULRzwUSlvQXHysUq8HcEyT9NqZXUSfNmbf
nHNYPUqGG2MMSkHEggC6TpmaaId6XYfPLrAFaFoViHJsR7jqvzBH9hToPyfPTxcW
5oYDBMhvxLZLDZAWB3Dox/P54W/X5TNag1Z5iHtHYTH0aFhshagagIGT+PRXQ+6A
Xv/Hj1Ocr1nNMnuYJ0WJCVTaKZ4c/GnBiOQ+PPsd+1CgEFAHjhEaaWpDb39KIz5z
q88G4a3eG5mvSLGkTFCgns1V04jruIlPam1sbpKT8TvAuFk5wXKiAf4SFhL8+j3U
/6vcre5xYkS3PoOuJ6WJnryDG2iXthWJBxqetHE8tif080r3TmQegJ1hnNq7vugX
1X79MZHa9I5j8m7FllyBrfEXUOxy3bDj0WCHoDbDPCTkAEKjkCf3AYL5Hjj/E2MS
bXH3dN2wyP/5SITf6Ul+hkKrgJP+kOtvVYj6XIoVGtfmTQSEk5dat4dpIbu3XtFp
hM/IBnCWMyCdAvrIUUkXhz3EVK6YhMDTfvYbED69Q+Kq3RNAaYBab9GXSRASV1mC
grrNWVn+y4szrXSX1ClMTlcOknW91lJpdR8l+GP5M0QMG3KWD4dVTUwzLfNQfNOW
PUe1aT2cFOze9XkS+Hm5hxB+wb6HaUtHe7G5+HNsik8yiRj/r5UOlIOgHBf7HzcF
H3A0ejM7K0vdkwuDV2JwaLKFRrpTZMFQhUCyyUpzakCkq+zFUQXx2zySIVcuqvMR
g/CvFDBTI9j+h3Tc8TaKcBoTG/ie2TKpqKjL6M/7tbrKMbtZRaqlbz4SxlBnLnXE
V80VYTtFdSPK7eI66rJTWWzyCBrI6c2D4u3j+6X0tiL0hWyed/ieHj2ope05ajz6
01GC90ABgSTE4vaA0jFzv1SEzCnLHIplsOkIgilkXVS5FAvnfz7MZ2t4OPcnYwWh
ZaueHa9RrfS0eoi71LM63pGV5DNd7uWBTaGHD/fm+vIZEvIIxGZiuNUZbBWOdmxk
LbC9O6FUpSOMJiDgThmpkTI99MS7ClG5GNq4uNxFkYT9DqMF0f/e9WIVlWkuZqCr
vu7R6CX6GZ+EGLD8pBGdkEuJllxNtkKxJqUlYvmcGYbIjaNz0tgG2XovuShHCtJ5
sgkqcdNhKRsLcTtzjQGkvAQ0U2J3ffDu/nHXSJxdQCfYw+plTFeky1tnHNPh0Cut
w01NdMQwjhFNo3S+k4CyUde2ThER62R/Q1A0z+eJB0hfJFwK9tqHtdY+ePnX39LY
xalCsCHqnGxtfa4YLMGkSWjUBEB5dfFEO/F9s6KGKuQl9gyMdPnLRaOzY6gwj+ND
D0aD4krs/Ks9qrXIE1rcdGba0UGnIA7cKClAHO/PjXWWoztH3cNlkSoKqZztYxRM
CYxWIc73SLCewkOxtXnDdpXSbanEv8WAfNgannHqGMzmYGWBU2DvGtPy4lVVVK98
LcL7VxXcLTnj41H1AEdhXVFVqHOoTs3cQrZSXP6/a+F5ZtANXArr3E0Y11MNFLgh
QurOOn2Rp7acynLOvyq/hUzNhHjh8PSj7uG63rOuH4PzSBu+zJQVBgSBXWKkzp1c
82/+3wrXm/4vG472eKPyf+HDvLP/vj1KclASu0YoZ6m+2HBMQQ1ch53eaJPzzEIg
xU+8dNXmwqsBtPiAW0aExCrmVaaqphYN0L1F+tFmRA1jachtAEF+j77bKDlk1gQw
RLwtj9Jnqc38FFXmQspLWmloeo4eY1Z3ebWvGCPUZDqWfS6OEX0upW9vzdmO4rZs
o03VOxtH0WUwWHD/W+52ExkvaDeTzQIKoWp3ILrK2onZpqi1MyeQFeK0Nmw8Fztc
T0DjyGyYgeJgoOhTgyOMY1gzFJbHQ+5SfP6+5yZRjiQ4v4Wf+EbQN3Tg+8MaBwVt
wpCcJ8zbMUgSDW68zT6ECCleu4iDwdOuMzalnweytU+2c54RkioXnQtJ2/hTmDKz
8/dv3hENHzBLKod57K4APa4PTZGhScw8Qi/xfEtaocrl41D1/yqGoVGjkA9EUE7A
+AxtGnfbw/PGPu8XjEQjIs0xe1JBgeHuix0t6foLT2W4eyv+hmugCdaXM6C19eqR
Ehm6D38d2iZBQGSjR6nyGaGviGvY5xXuWeTZh5yFTQOkqW7X776HQj2/CMRTGWT3
pOLoK4DUftfwFroEbeL0JsOh3pojs89a44xdR+PUqjUiUQRAd52B8lQONQ01ut9F
+QpVgxDbMBcb/LRuGvtpnd3je+benRUmmte0M8r0R8HtdxWGdxr63rGMltrsGNLy
gUj3p9lLYyQMVKOhEYTd4PQe/NRFvGgMaT8Lf/E+Us1PdabgICer1oWGdP/Sj/c/
Ukr94wkm5rmSWWT/0N3KDswGYyuW/E6ZKKnldFphKMLut9FLlmAEN9rMQvBrfmVi
lBF1lt3sRWi05apQCvIYOx2y+8fF5WneuBdFWPzyCtdWn0m04xi5qgnaK250366b
JjOpGI9AkiolPGTnh/Z6Q2T8ueOh05iaE6GYsxh2jZr7vBe/bHlhyqKTipcBDLu7
k9Ojp68jpGNnGtegqiSSCye/oY2Jq6ReP6wgEbRQaVKuLJt99/HvUIkI4FCbLv0k
wi9zsaD/KMfRTOSEtLAjqE8ShasT3dGvxpq3U5fFKTHeZCxBZSV3bkMzJZLUcd9S
CIyygFku1lbl29Z2b8BJWmbi45Tfkvaen40cyhgSTwa96qoYF2EA6WRDDh69ATIs
WtHgPUqRJBkZZvJDcZv3OPYJjnfOVNGr1MUm/VQeZF9UxJB4LurSNXtYo8/SPB6M
l8YI5R7E9LtYDLiJinPbpNA1IeVKkNnrYQVh3OKNKvKC7mVn/L2smiqXURWDtWfw
h+x/pvct4QGaVoKiMO6E4q9g12xEsAyJkwsbHqzXwKkeoxEkQDn8P22dGnBrqMO+
zr99A7gQ29BkQ9FGGkj7eLsVpSP5X+b8L/wswvyI+KEvdb7lKhf+8iUk2a0gZh2p
Kv7IvTSI6P+I/hIYkILtOh4L+/kqTT8lfzl9uegubco2yfXNgd+9KVr7bT8xxRz/
YePEqmf8jeEbyzrJa/Mz0Md1KYyie+hZL9h008Yqmqx2fPTXmt2ZliNsPRiyumBT
pOdwDYnuyAmQMSA5WXuCV7DiemsRX4jYKHlcN0BuWyKp1cH9OPwtcuxasIy6tDdk
uH7kLNAVPhK9vDqw1Orx936N6omyGXywQQyEWaxkE6JJEQxri2PM6a42PZU9AQA1
thuYp0GD+iAL4/bt5eowV5eEKIwDdLvjUfEVd/1V2T4w3S1EjimmgAf1BV1kOLwY
J29Jpud8pSfTpnF3yxXoHIdvlW/8mY7B3axX3bhkBRH7Uf669ZaoWh2l7QbgzwBW
/0a3qn3x19csI/gHI8sKAjfv2+2c+2ScGLGKvkcFEkUg7Jl0/W3vKM2R3d0W0twO
QlXKwsKva5nf0veLt1iFNDo4WoLeKXGx/9enzOjX/95gZh2Yt5kob/ID5EFASciG
3OxKzVnHV00eUj6q4yxa7zAoAG89VEJPmHDq+bwpuuYEhrY2jRnzgXNfkzCa7HQh
c752J/fhRByDNOMrfeDhzMX2AWhV3fBW5KcVUvvwlvMFkpuchF709eN8QoNyC2mo
xbbu28zUGwGN9f2ju6kjBqpovFPkOLzHugShCaJ0xg/UjULy7Qs1zmtRIOX0LKwt
+UIyJuAf1wkXhIK005eDhPY7FcOHBb7fgcINeDNsKCohW0QLcqHecxmZBx2grBkw
Vg8cVVPSR71VKdzk8Qaonq6FLKQogfeJ6fP3riY2yBl/CbB5Bxc/57C8IJaRHr8V
KAayWq58l8jQk5g5Wof+33QmNcmD1jaI9lEFn5X7sJ/7GYVNv2VP+eat1YKDzMP3
EmCvwV+qBEFihpRidzo2Ma0nWPrVYS9mXoA6mlDMRhXZzYFvZnDLIdmVrRyjK660
RGj3dw9g955bmVEes60rZslGG68scg4UKcUaRYC8ep+Q6WiyyYC9/dcc1K+UYwKy
PEwKvF4TrJ60K4SBhCZ6iiGcf/pmkPt6PZEuJHXOWh+Y7bFUnUVcfWkYhCFU7Pn2
L66Thil3xCSV5LBr0s5QXgvZ1ZJkwtl+NSOPkakejLgbOVmI8qawf2cYdiyISqsm
qmYUma8Ftt3C45MTMM2YGvkO+lRELtfS2PpDbISbQcFo1QZS4zSn9s6NTKfZkfT8
FcjLdooh9jvpAH5uUKg26ADfb39hgsR4WNPpFSQgmR0twafOpp+jrCYxPYeMCjoG
1l6GaV9ECWEKscy5zPXyCzsXB5aQ9opfaSdIMJs7iKe/+vtsWI9QluW/B2DuAtr2
zbWNq+st+q/yADNRxfHXaTl7vDpcipS9A+x0NcUo3pq2k83n22LG9lr5NOFwvOx6
doykHFE/4FzynVBbmuNFH9ihYza+tIMXQ5w0S3M6ZnEf1eNDdaa11rHCZzax2L0f
miA+xTB+sNywgPgnfWZjFCfaDfKdZWIFcWcMUxDsK98Cw3PgUBS10Wo4PkClyvUV
oCfXiKLilNm9KPRt7M6qqfOZmSz1b59dNMjhBSfGh7WlR+WlRQfkDOxJoN7u/4bx
F5YCf4L/UktN+WN9ubzX2mfbu8mklN1XLi2qEAd4sxHax7FnonpxDoFYeudLmT87
EE9v8PtmqjoWDfGbsSTWTm5gEoji29Xjavy0LE49RZKN1IJp3ezdMDjBUVNIpoyz
VMKdRRKK4ysJmP3hEs8+p7W8mUrveBwReW4ScqDxE9R7la3mJgTzzO0qZoudKkhz
Psgr6/BrbCswN8cw4c4thzXhzPtOmYsvOZIyOdq7dIi161gh6St0HV7y076Iv0zg
Lr1FqvE/hbgoMas85KvTy438Etcaq/XPBKpcaLJWxTcCKZJ+s6UBNTurNbomeAMc
xFDAtv84vS9R7hUBohiBLIXEqo1DgcadX23Q6vTYEsqlxJ+sxxHi1vXL+oxuqW8I
/yfD0SddbwNsb9+8Ns7et6U0ZidLLW37y1rMVqhZrMZV4GUlRBd0T7H61PWxQ6DE
eWwDb9skG9mZ6LNaQXQdD4IsiYj0/Vq/LfoNdcFwjZ81kRnWkJTTD2GDjuQtH7hZ
GaUdgXCmupu0xJzBypVdq+M16PvFgXY49dg4/7JTa0b5sOj3njtcerzrc0BxSABv
j6lAe22qPRFtnhqTvtz2CtKsXvDDQZVZc0R8psat55IIGZ14XVdacU0vYPcTigUD
cj2OVGN6bizaCJ2mAxMJtTDMSwYOg/nz+4x3Uhl+83gzrSmILeWBpkiM9JjvsBvO
6VWaHh/YrBhu4mx67T9ZhazsFPronIvWwkV+zYV7Hj/zdZstCzl1KnYNMY1f36dI
CSQbFbj1AKgeLeR9dn2x4vk2DT/7OnLlGwrDB/cqBBMovDUgdMvFBeI/WKaR4wXn
o69ACCSJGkt+21M354IcTipSrSVPWA3AyQjIr5eko+PAhtOKkFUifzuP235q5dcF
SYYIuEGN6r5cQQEQdprqKhFOzEvjDqo/p1EDvG0b4EmihkyUZCZVNkq79//MTaGL
9DXx23HgTR8OzNbJ5PJD6ZFHHRWGw3KOLDasP4mLUPCzBY2cZO3vM/nwTJ1/cc5g
TloPJbKC1/W/gr20izBhbLK8ksr7C/XBwTKsKsm6LnZfgGfeoxY7jezDACe4tMAA
eWialiyK3JczODo+P+ejzeRQrowd/bOGCV+aruakmA4ln2GzJm3f7L/9OfeZXzSr
eZcI+gcqT3A3/EoMZiC2wSZ85W85DqgIXLpc+0CKApAUy61AeF7se8W3r+YCKUVY
ibOVkjkruu4HNAv11cv7fWDWXon+w7xQmS5s/nCZ9hSImjRverR/+vwZsFFAKPWP
XlQ3zVEfT1Pp5eQiVRuSZBAMXQ54RJVHiPNpmJRM2/r2UzoxPC5NdYmRYntsGh6m
OTwDK/mHxGJlWD3kptKdc4KiI8GCMBP7YagehBfFY+uTxOAHKBJDAoBuvK9B+sJO
W2uXeKM5Lfhy4HJ+BQHZ+uaPLbHCVJ4b7PdAlI5mpKB8bLNqyZ5EVmOenOpG0ptv
72pnE8DClCAFI1Czz8j0TEMocPDrZYOxjJYqimdQxypjN+VeJVzd0Plyq6cXUVFM
YjE034qW6Lq7vFHUUY4ahMXaNqk5ZrCY/bhpV5rm9EHHNbqXq+JVdZlIgAYSLLzl
DWpxcW4OUnStArzuaiK41jj8bajVe7ESoyuGpt7eo5f2iniyd2Hifi+5M8dbQVYQ
gW2g+BT0Il+hc/ViST9TWh4Iwua0CQDj9yiGXZSDsILW4xi0IN7fAsbxTrv5czAT
OZLONCauvze0zL2TIL2+G2M5sRXRjti6H2V8Y2fz4ALup0Id8mdYptfKzdqOR9On
6JJgfivCYQIlYNpS9bGaM+bt1+C3eslbioZq6tFCy5px5v58jdbQj2JcurRw6JRR
v5ut1sqQqf/ivfZJro++S3rJfFejqRLZiljWcfqjWy/dg73pqSqT5maxlJl1EyxV
WqfU2GuONr2EAShoaKfyUsy/eLnxbhZOxxYRN8eWgz1MqOhySNBCcmKRxnyjxcZ3
TY0bQTj6VEtBa5UDkAW4+u85Pt7cTraN5YNF14wAboT8cdZNmYtJ6AL9K5fJodEv
5xq3fKUnRt5N8mdvoyNdsoAnqh1vEHsRb31mZtm1XSypUa+LFEpr5bfuaUXIw74j
FjUyJWzNjbO3WqgLHyIcr1sWuuorTqZj8sAOw9YM6/PPAPmbUmxRZcdoHYLohXwx
pfl0g4N8dGG6mIRT3hjYN5SiPyBmQHM8M7Lx6FtOIORSwctg5MQ5A1luMQzaOD+3
BLwQmYvla06QHNJ5FFvZFKgpTe84ZIDiM1jhe8SrAS2Vef2f/0Riw+AwaKSN4rqm
AF/bKE1XAuCxxKgBqF+VgE5JxtFFf1k8LOPKzclquOR8c0SQkQAHQWsp1eJ9DEo4
l0DiKc16x8SDiTVbJK8ja7tcfcg5JWn8xrGf9T6v9JAzbLZcuXLHzQ52TuOF5EDE
Ri/D3y2z6ZqpvX3j2aYmiuhB8xcnauJ9yxQkgfDVwtbBJfht+W+m0PBIQ1Kg7aab
lNwlv88+cusXy2v5/zB8rKHsOZc1PO5xxP+Oorc0fFIiQDXiTkadSjantBfCGNws
cbV4Jm3szTELmBoaVvSAciwhPSKY+UfaLwKwKCEq1+FrQWnW13ssUucmWZWb1Sq4
2PwVb7Tf1WXHFgWk2948FE76Q9W0DA5Tnl94a0ZQA/C9T5utKzjpvJs/6BXdijK7
3O4IY+i/UDyELLYAHBSrZGwuBnhMs09MJNmVASZpEvcJdODpeznH+YGnka9Jvmf4
IApHWTEkCYz/0iexuxp6m8IxFDfkQpGm6VYIbpey55taeVRzJCSx8TkM8eC8CLet
/ntlbOyA4vdB/P63SYF3+BJ8C/y2lmqDlkqrpG8XhFeye/WPaa9jgBG2VPa+dK9x
P/H+0+8uGQtMENpwovu2McAA0Lx+2+Wz32HhOh+s6fIzuBYgTdBcHQb5B7RPftle
KfuRTbQk15t15u5SvimIWcO1nN0VGbcvhzYUFZc74ElDIubvq5AND478CT5ysRVf
cxdo5g6Bh/hGbkkNyBs2J5qCoOqq1vZzh1WM5OALrzM0hhOqb7yRlRb7W4/1NeTG
gDiszesQRfVwUMVTkFuIZcvfEVQm4C5iea2mAGDFR9x1bVO8VbBm1fdQur1j5f9y
T+Ypkk9zHjgRSGHJtQrefVwXsqzwhnvwmbgrvEzpanZsMFu+NyPgm4k2tTy+pg1D
N7yyBpp/ZtwmdGg2hyHxMUNr/W81el7tOlH8iBeh557p3HOzbiqMmFjsoTDyipoT
vI7hj7zEyzVpdqpwd27FkVPbj46AkLhRi3lLM3kq1l8I/8O/1yyHvYEtCBpT697z
FQXVqX8a1gWEM+K2FQqF8bkdLmBfWp88TY7/Z1ZiSXcOAzTElWual37Kw4gA8+n8
zEe1VjlO1nEGk28VT/ejNP7/yomPkktwp0rgm5vHtYEZxUwyYxYqHFhNTI27R6iR
kj62fuCg+R2JPkvZ88jjghbLofXQMdN7rnsQNMWTWCUnoWlJmaFqcdUKynBJ0bY5
wOoNuQyouotTzisCSmacdfRXNjo69G5BWjVlZTJkWEogODGn65xBk/Vr1EUxen9h
XU7D6gRwSCtHa8W8vLIC5alj10Haj2ZGdc2MMZSfF88yy2AMxwMU79TKaxnzZQ7G
AegdedXlXbf8u6YcEIGDqHdgvholZVHYd9wCJ2MCoH6b3De9+tlpEvD3wc8DjxM/
ZA2LcEiaZhKjOJEmqPAEnHHWb9iZWpeLIrnIAF9j2PV/cyq5mw8FW2aUHBxSQp67
vojujOV+hNR6uaClsVV8IFYw8nZWJ/WM+ZBF4mXuwcvyirldxqVAISQK+9I6/moI
L2cGq7gc00Z66ARauvmf0ntWx+Hcqxp6I0Yul/tAcLG9q40EPKIm4vpNAe4vttps
wCOtCLyelDxiwBdSPEdsaHyzm+vIuvOJzJ7oqA9VsoVpZh72Dmo4Z+B89Gxzd6dR
dv1cGFi2qQgLgwH+PdSFqPdbSX5FSJd8J0TsUOiQsN4KpGNr76UuBN1y2VWFaSmj
XQ0ak6y+fpQzGPHdt4r//lYfbwVE9mQoUHBjBAMkDFGxsccUTGdTUlrxX/SkZF/K
fNz5dXNGUWcNqG+fQalBsYRL8ZgYe1LXrTi85fp4gyOQQqfRVpNbOhsplEsAcXZh
/wpaIp7OY2J2L8S8UoqqWbPHB93A7ciJzxQgkTvGlTxgMhfJWOYh/pPzOKOwS5gQ
0tu0yFHABoi3pASxB8eAsDsSUf1eyF9LurBYQLLsVdfKf8y1g/OND4J773z0VsNZ
PzNKbhr+Fx4GVW4enw+HZA8EH0AhQ6nWQQe0B2QTDs83kkUPFrRqRVHbxYHXdqZx
N2iYHsko9Zdjl4IX6MEmrfQqPbckxKAFluge7tEYyD6vCGSZA9/6acOk89RKCS6q
m35BNn5KKU5EBMroFpS05fj2OtPglBGhvzKWQd2PRAqywwfcSRpOtiaksNDHqQg1
XSnrQ6Aaavao2858il9cLnE6gBl/oqIwVDJoUgQU/eWnHvJlwhf50kMdMfX9jUGq
Z3vpCBJZGi0tNtc+6FdB/QKVeMH3ozVIbqWhKhUlLhtoVi3TzAL7H56SR+CEoYyS
1nBcRtURBNdINNUGR7O6SZx0oz7l3Qnld4lsWaWQjKDR3YAw/lZesNBHKgpQT5ki
Tzk6ywJdKHQjxAEfhp41HPzgWkA2yvgmEMdqDIS8skVaTgNhJO50fBXgI0nzfPFw
MLlDszYFRIULSfSNTmTkmSdvpvVNv8DP1o3uYvG0vI/u/QrmwfsD8ac7F73OB3MF
lVIiX/JQTgVHGPDf7LfvN9MePx8+gmskZlCyxKG9oxtXrIi81V0wAknI2Yeas6d8
iNpXpWHsMWgUOajs5h/yB7DwcfLHu098t2dyxs6hBCe35Z8OuGDVM/hXHGJjsmJF
qoddimQ0Af0BZOL3weYT3wKRdB05LMCFt0mnGRVcmX1ZRLXUHRAfXIctDAp7klrL
hked/P/RXjPCz3ezboiXMzcaZ1ttQenc0Tw0vB4GmmpVhpkD+XFlTJCYtt4lHCV9
8ren/R0oi9uxEN0utXHRIZuqWku1jM10PHcpmItQeHy2xwgqvNXBXabGHe1eQdkJ
He89N79y4DdYF/bDaRRtZ7ZZtic35RrIu45ra9NhRXy9Pve/AC9M7AgnSe58qf8v
oZ4EFuj7LLFd7UGMmBrDvPHoRYpmytU1pJJ0R/Gw7LX2FOyhrXS1F3YwonIll4fG
r+h9pnTAQVeVS93UvFHYDZ+Z7+MsWfIbIaIyzzHS4anYcFPb9sFcRPd76n1om5Si
V9pcKxN93QNDSzr+CviON7ILhFaUtbzNPXXvJOLVywK4DbUS6GpKSesMLF0qf44O
ys1gqhBBz4e35yTmNZc7ATjGVN7kE0NLlTcJ5g+CC0U8/yt/mxsweFG7HvKKQYv/
V1tUuHELST6owQlz/YubP0iWTFOfV4PG2qGLh2ogyq1QJDBSfS2p2PbVbleDTrd8
4O1sYbQKFpdB0JKrn7K5EHb/ziusIIwW8x9pf156I0FsaK0gIpZ/3CgyxZksx6Sy
y81bTTe2lSk5RLzUxLlnFqPm+HOx3WBGu9lnhhTwe39a1h3ZYKAo4lhLyRBv6b43
dZRfHMOG9lEQYwsyH+s+Bh/D5tm82hkBUFHmDQsOK/yRDvUTSzcvJAMEWtbHTInu
rTFszENB+3EQ+BgkYsYVkQHzziy1B3tRHXv2EPQh0hZ6o+vUHb7CylLh3kAB2svW
Vt1aCIOs6h9xx0KAJ/edbTUPkjrpTShQqCjBDsWZ1OU3UM2yrryFa/Wk7dggpfil
eOFGvD4rguZ9toPjt3jP1mS2+AzP4IDPowsqYCIc/pITZw17/Zx1xn/9mXNsMsrs
JdyztWckymeSyDl7YzK4tAGMSfgL+X9rSQMjnTVeP211/kfXLzO5L5ClfwrhKT2c
XeFf9capBjiMDH24uKUU5arG92wTT1Fei2SAqkkz3IkYjq90mrvCtMJi8nmzF3n9
ygyq6s8rXqQBG95k1nR72UvYnSQSbUfSp2+cTWwE9fUueNFoNIVywrDH9aWnU9yV
8clB/fygX+NFYFBD1tUmM99lb9RXWKKNTdnrtv4+WoLtKHbA4KA3aP5H+yKEQNON
BYRJ/1utNwxvEfGbz5FQp4wt9cJJNPtU0MAmyE6B9tMwUBFqOL0FYmbQAioq3/d0
dWzYr+4hQZPJylcPoiC1dhJWJKP3ITYRpvXQ2nqpIj103no8fQxX84oH6ylychBa
M1lLERfWpOMuNWGLc8qbkZq+DIL0ld6rsp6OYC0FyEmtIFRTGV2HID2zwobqfGvm
WfB4pbKuP/bxW5YpKsugVhHaBPEwD7bMqc8rUfJTcctLkMHkBXrLP0nqgRi9hQs3
4zt0K/6K3TYtNVuXWPhowFw0dZ0A4ONl7MyB0duBaFd2L7Z0pdHhgnEhTaDFxnCS
H7/qv9ZhAdjLengBHkSC4C0Nqdzj7QB0/VDIO5eYueer523czSHAtdJfcQ8ekH7P
5qk14j6fJt3MU7muBA9FsDXGw6KORxm51e7lNIZW9rUoj4zXt6iYlKu8why8ayrx
cvYDG0i+DYTSCJcNZ/YZjpc/qgjw7jL29Kpze9B6Dg0qd2aTwktOO8Yk1CCyONOy
LHKStEdjFhgKcsw6TgxuUkenJROsOOZQeN8osgx0tce9115EcVOvCBtKGDUnvvcR
2eUzTYGNN+cLhsO4Do0w+9RIzUdtpbwJU5kM24kyxtDpd/v4qsjyTaOUaEIP25o/
/87yTaF+euG/fzTDuR2bZ8WdfzOFaMQc7WGJaddbfcOm/X+cnh2oqILCyjDlQm9p
EKSQVJMyjUUFXaNvP9SOVy2Vj2SaBYU6SEB6BEv3gfvdZQi/yQQU95i4+jPTgL3I
QaxeYNd2YTE4KZ8z3idoVM2962QqXrsMbZlwM/8APC1NE9rLeLCGYUqu74Vjme5v
e6hveCKOTg+C711EXV0JqtLFsBgq9/lijE9f6Gtmt4TVUu9ObuTfOGvAcI4vUY1D
8P8fbYu90aIDyVIEoDTjOfpyw+hlPsVp7HBpQTlwdxUOlnZMHXiY8DokNWW2XgWB
Klv1NHbtHooDivtCBbK5Hm6by0ESHNUnKWLBdDV3fg6ehteh9aFa/Z66Tzeevidb
Xaa9Zqp6nj2LJdmkKFbzCVU5im0BCeNqLlYGIAVZweqyUId+Bkpkok6lukxSop0Y
Qm/JPd2rQ9KGlQ4K+5yczXhT0gXF0ku3jK9MqHuZUBCqoEJS8nXdnzCJ6SSklksJ
oE167EipSc0d9E+ISdm1OXjDhCvtp66+FYBSjBEObvOoZocZDZK8Wb1Mv2ubUaWG
GuhHEkehRGUERHL/Dw5hXF4rQU3SvDXkEHj4bvYvCCyiN7QoNW5eH4+EL8pBPybF
GOuyb4u6gsreL0kjk/Ga1j4fGZgMe5DPppcBBKg49VhBZmaNYu59DuQthj9P8LXv
EnUXL74sEl1czth0gvatuimbk2ge5euzWCI4hpLbxnssoU6WLa94L1Hdho3D9kDC
GU4+l/MhsGgj/hBYtHRY/FomVN7rb1PVdJNVVlEbmmkcR5VTvMbJWO64DEVTEbmb
MoSvO9z4aH88ESgDxt6nd7ZILlFnH7tnRG8zBnPMBdTpKsMUXdrOmIZkzb1uUvDa
ho0dPNEE+7cxbG/HRo1JoaRWFbHHgCmFOYi9LFrhIWilyxoDBlqwGqDr9CcQRre6
ADHyn4o8+kAhwjMEQzgZAWqIEwKKeh5M7fUiFI8PkOfeyr2k+OAtuBAOt56/bZ/w
CyXlFv02tADE3RyV59nu07PwA3WtW5iuY3hI69h+/KjuZoocnLbNtWkSulo/Rf2z
dziPcA/zJXqSz1ogOhFn6RqdcKlYKqcAJ2RItu7XhJYIG0L9cCrYO4udUvHmB1YE
PIm8GMTc0DX4bi6GX66MlaSgUJJIOlllNgSzP/4c4b1HA1pjoRQ2vaoYnRFS280G
pDWXwEi3N8R8O2WGrqA5Juy6spkna5LeaRs1nRf9A51p9KYUjSPMkwfz16SqAwV2
0IkxgoUE7MAPv8UxmCToOIHRUWoZIV2vBUW8QBURd9bfWk8urcWIYLakHkbYpPHW
NVdHMassK4EKwVjxjkkCPRLTnNx5YVI0uv4rSIrAv7f/JRSB42+PPOy8Lwgpr38P
oOZRD5qcLBCiapKnILEqhvDW9UZEfoCp5rTdOEouUwzL27dOBSdwJ9dF4z/0t6NF
1CeIWPcd3b3u3/+lbQN4mcYIJe9h4IYzlxjJ7xJkkiCbaYdXUggMxuTE12TLngBy
2v6Onni0rELVBjghWeYaacXZaxzcNtiiujEDQq+FnErVO3Tw0zy0uH/m1GQ4zlaK
RDcWHsM8dXKcsQdbx+s79RUJrElsXolzLwd1Vp6csexIVMfpTZzVaxXBFf9smZwP
pMieBAVUpybE6JaA7uk/xhm7n/bJjGehguiYineV6FF3isT70I4poh5ByjemzJgH
iUaHVJMyCdbzu+tVZ8hf5bedBUiXY1Ayh0PphSz6J2oMNONC+KxZZ8EfsSF5DS8g
rL/9aA2fEPzzsRXejD0aTPUf9wVtfQ8AAOQj9I95mj2qrc0uAFhThiR1pYlxDwAC
ri0OZjxllnlfOPAmjEuR4Y9SeRbGiN/A8qzX4cHOgGLVs4ToMYczfpas1QxAdOZd
qsjtlwCIqf8yBV/0lgoQkXntyhYdtXCZogcWbzDDlZpdDW2KqAvErpW864y9DleK
XRDillfVlZhb4W2Bw1ScubJwKeqS4IzkY5yma6WGszt8UgzTPav/kPnPIXGHcUap
dZVj3zaLrm0AFmc4sULif6e+LRdPmdA+PHpxM6CcuVxOOgwwIDaU63IahsbmzMZt
iXHk6jc41TPbQ4s6grcmqvwGJRxt58v3LcDoquUbTHbw1aoM19li3TLJGL5Go52J
UeutcPG2g1XIsE1COubB+YSrui6LoCoVOvF4WpJO8rxDer4vzbh3Hd6curLBFhrr
YbDJrJUHyvPpL95vHAnEa/8xAbokPKP5sf/izyDR8v23+X+bebAsaqYwh4Bz5+Qx
T/1bMNuo+VmA0tXWD+z2vfWzDsWFMqhzfciaI2ev1FLik4e17ieweKFjJrBWSRpD
hBt69tZMbaM/S5WUfjyylGHD37iE9MDkREAzLdzobAIUpOITCKG8V5kgX+7mGgiP
mljoGxWuSOUrt8s2sfrmw1NwQ9gI30L27pvGKwJtWPqFRY+BVO+DC8MFOTjmtqdw
wFs8BiqbiXqgtS/kQ79vxQyB5OI8Utlcml/CJDUN9yZDYaB9pxOhKuIV8tJ4A0Zf
G3EsInZoFpMHxMQRggh1HmEjwyYA1ByMTLo5FfCcHQUuXHP7DbD3HwP1f/xV6Xr9
G/kynNq3hyg0lAZyMCjVBL5YhIjLKcds9v384wzTVpGRWCunwxz0XzRPHzJgSkSx
ne9/Ivwakqw5+LKtoUEOUTUqNT0hM2wub1hopj7+tD1dWFjy+oC+jfmKyPWxp4Xk
UE3tydMflhVGjTG8s8f3mNFaHRHr8EoQjVy6YRkjXgh1CxYvKFYIwqh2+Il+sm57
he2Av9tEfV1kLjnNmXlR404qcGdJTmmv2UxK1LKoamoj8l1VgMDbfVmM1aFCW05X
H9bleS6flMftxvJQReRQSu/ecAWmbzVBiCb/VAQ2xtFAlmwbEQJ0Yqg621ZlqBNR
6h86/UhG6s3l4P5cGOoJ6G3LloneXH6geOhnk6iKZ7/U/PjZgTN/HNpFyFQ2T4Ev
q+p4lZxYBuSXuTr5oDhQXlfVrg46GA8JLd4siWWf4ItaseGcsEURVMggfBxNTZ0L
UGm6fReJnDGgAwtAJ9a4RoNzOIShTs9PV9LHxINHl7UZMuLTn1H/ycLZS1K/Q5Vi
Nglqv1B/KjS20paaQNaiizbRIhhSoU5cZNObBk0gw5oswmZhSgl/vR8v0dkFLvah
2t9NjGVcASvBWRbIE0h1nEOc6jy3aj0gpiMXT0fZdnjU3kZo1HUxCjFnpM8yI6Xr
5wttD0KFcM92w+SigbPUtoap0+yi4Mq2zR+s0SdNGPnqYzwr/fS2BHqPdCKR1opM
EYjoR/dz+/sPOgKKerSAFkht6b/W96IYLF0lEXOcpK/LRrFz9EIEVmUXQi4N3EmL
BjqQEY8GzqGjdicwr9lYS7+0TGHTTj2hhU4ASLGafsBiNgG0wlImadtZnyATQqhr
oxMIt98GrBaAE6hGZ79lCOQZJ8aDZgNJW/gn4p80A4Z3LS5DAeTDK8G1OB1Vtckq
syOlwwqVZLRqt7D2hgJWwDT7Jh7wRi+kbs0+rzSCf79nQdkAiUb2a6r66d1AgHwF
u1KcuQ3fiR2DjTJGwL+UBxD02yVk/SP1SNBLB2SHEaKyRsSkB3zF4PgPcqFpEs0d
RKKByy7q0Rj0aiDj8TGSnzeEzU8yYwUiK5TO/ZOE3SRw9SLYdnhpAKzZ8Adq9jy5
ZlhRR+vuanzw+TtPfLbzc3HCdV/2/ojZxhlifUbN/A1112fQXpid6mcO/C32VNtS
DJP+J197d8o6IheA3LSI4shXc6hh1BVKEX0oFrVDBXVNSDw7OeC1pN+Iig+nEPh9
Kg3ltQ+p0iOx1Rsr4WbnxIJfHo7m7RVseE7t0O9itJJjz18CfxBPlpB64xkBWO8A
VacIk4TgVozjENqPTYKCKYS7j1ZPmU/fnIhANL3p4GAQ7EDo8O7Y2A0nQh+vtJbE
BBA41Ic5KQzSlLnfZXReQ7HYY9XtzzjAI9ub8xFNwatuuHnjkk4EMsDxFWSRQoDm
HBA07BwgEpRaACbCBP/bvTkGZpeLianZS554d/mfQiHIIsgoACis1rGibOTKyd67
uwSKADmH08w8dB+JurqdBEB37yobHldt5XKKF8yZP95xB3cD5S/mi2WUtFE9zsFN
YxpGqWA2Jy5kTMJVTF6BYYN++dZdV0ehqGOjk0sjJACmnvtT7BbmWak02xII6F3U
NM6fvNGfD/iePbCQaCpnA6d3sWga/9hy80q9mlc2PNMFb6fXEbcNQd9JUtdt4Mxv
fOSfQVUk43YLw5QHsll31M3LMuZec440oWewcwvWKEj07ATZlkQ2QgooQeio7XA6
LNB169TrZ/XrgmjJW2s4VV4fR3hK/eSaFQcNSPj5Xd8Ny8w63IRHnNySByJdljcj
CWz6U3PVwg5dlTt39DIwHvKswufcXf66x+/2avPlqhosuxDWC4rGbPweCoXA05gi
0TrM3pKUn9nWs5fGWDabTJzWjHs8tN1KxsczyXvsnVOIww5sp06QleEuDoU/+qDw
PriF9b2A/VpvQx10AMHlG7Iu4rwY1Bb89ou2UjrpnXEfasPj1AS9L0n5CofQbNmf
Z0wEXlTOz2aU5GgYQPLuBLhjCHbQPgOkiCYWqT8I0nHeFayczY8A1jbLDHEWhdAx
bssMvLzKUtt/wPPp+M4aJuQ+ILtKw5QyttI3mRO4EPI/THlfRFQq6zixkC1tKdGL
lA4fgVOGomTtQaW4tmAucMgVYxgZ4uqxv4WvCt1HWHR0vWGHJMoP4aLt9nE3SlAU
+u80GJR+RfczLa6hAuOGgxS4qrB98iQSX2hoa9Pm4hiEB7aGrrYIUC7j+MaNi23k
IoR/GXAHSupjh/z7uYBFAADbgSaIk3GQlRgpnEyd68clW3h3OezfDIJMjfi9BmeL
qBy7NwKCW3YCXk1X+gcFpE4yVWWNVcHIKrILFkS4Tdb8v2Nd0JsTesUi4YtFDeZA
M5wVUvbiggkNaUv6NJ9iJs0OmkMqsAlxd2iF5xppLL1KTpVNRBNiTu634AfbrLBC
gl6+uTUFXtnZu/sHDGGoyqxh/nzWBhnbqrXVxKFXJaoJZWNJf6yIV02hIXuIrdXY
wdhps4tnHFYIJ7u+P2D4ptMfjKrIqblJXRbtA87sY3ewoo78guds6O6Z74URen8p
mBGimNR1fe/0mSH+iE+5Dm7HUfUyQ6wdNs7QcXOSeY3Qa7F3KzrXjJKYliM2zNSH
QvqKTb3sK4RJfBwzu4H5J7OtIqMOlSt/elx2UnW4fgMyEZezF4hpzJj3LVzkRwNz
OFbId3458iESONGqKEmB14jpmjOx+SXjvl4r+kjiCEtYIWRKZe+jlnddj0aLeD8t
PCCyE/Te92LBQ8yb2voXCyO77xQmc7o6hTmIQlg8qJ+iJ2S5KHoN2siM+dVSW952
tIX1bXFec7nyNk4AvLKf+V1q7b6I+678h9BhKmO4OGDXwvPt4L2SiTzMUoh8evTR
8urxs3p5A0ocd7wsW8alXuahLt3mtKXTm/P8cVYfF3Z7P1YBSOmJW9pgWvV6riP+
IooftAZ7Uxa07Zp7en78ulG7lLqXCKeX8CIDKBdJhEPQhr2SlqT6LkvGbUOyPqed
yh+KVDSD/zWGvURM746MDABoZGHcUZCAABZtDy+mrVrusH1evTkINttrljpeP2+E
ZkNfTd3/9zlNHvRa8NeUa3tjc61lR+nxE3ujw8QGW4rBw3l5WrHm1PqUJkz4F1Pk
0selE7NXwub9y/ol77KBuCo29pSEtMqZGPH0/kpyPdrbKJ0+xnx5kX0P4c+7VDyx
v7px56ZR+0T8TpU2EgpvpeyuNcCfVWxsNgXrxeBVpNAuZKGmgw2yxqcOBB51X9+H
wHsg/qK2SPB2qBc7nTnrW8RnVqeC2p83s+E4KSis26o3WPvqNAY4Gk6DGpnput6H
rvu5CvmYcJbR/CBNM9LB9ISOXbl1ZPy2kF7oIn3dGGdVHDM4aNJHdOA+Ca1LAmmV
oqjrJ+YSeiGp1DTcynDbp8fsCSZEm1yVWu1WPuloouotg1M4gPiPx5NwZo2BJ6WP
zUWjTI8A+HOf3FoME5C1UcV19EGe4i8WxCSBxgNaOt9KyS4qf4+/2uuKxNzRV8SB
c+gBdQYTiIHBYyHfW6Ba4X2eYy62AFvFp7IvbQCdLPnsxhlWmPQF9pg2uaRtDLY+
pAYDAvBZKJJjLOn0xJ4968wSRI1QBJ+IqVbVcVhHxhWgtnflQjsxhpfKNBOA4YUH
Y5Xu2/flPOUwSj3pjB4NBX2q6+OtAWU2MYaLDlFuWbQnzLq8o5dkQT5/ulmIgwD6
fU4O/qJEjBp+tBfaF+b789rVSilGoHAEAPvO/0TqQ+kaRq2ADIVVQDurrpou9Muw
LPrulRO/irX4wthtct2oYXQ47QFowkmxYzMWOr4b9UqBFpTAvivJPJclA38DWOLm
JVKfLPUQeKklEjZz5LyWc6+SiNUrZOtNlcz93EyV3wxiSZKYfysOKc/qnzCL6C3u
37UYBENxko18fwUPKFN9X/E8yfhPosX5u2ulbLu0MQAdpb4KnTjiTy/ZKJ80bv7Y
nTUq3rVQXgUYeLuxhPn0jpOWlrky84bmlBiJU8Ey8KsiKYjB/Zv6Q8TLzdts+lw+
8hkLYQl+AklFIr6l07TOQANC2lgrHkG8yIJxlyWPJ68giAtOKcv+IebHSBI3wZnk
2wlj2uvGGGq/T02JUgV1I4R61fVowbHeTkv7pNNtE3lXqPqtqgLjZBx3eO50f4M0
t3Wo2pom+hg7RTn1fjOIiWeDquS4xdh4dGPw/S6hhn6QUzdM22AmXG4RymPE/JhC
rK+PYUMtjkFSXOiYtCxizHTw5YIrovVHhgoPXNuZDlO4bpT4EHH7vlF+uSGzvN7+
hetZr3l4d99LnWzG58Od04jx8L2De16jGnO9pI458m77OKJC9fhUfaWdZufExP48
YYC6ShUH3r/wvMg91nWYt3E+xIug+ZiRYh0HgvUhSREyWC9FsUtvN+FJBgUAyELv
TtgjO+E134QKlETRA0W/yGGsJ7DQKu9yZqgTZybVV+NmjBEs5rgtFElhcrODAllE
7MeJTMfSGDMbMvZ1muAk9FpOJXjoyQVqD9RLDQpwchipWan6RJ+Om/bunkAM/FxU
B+szETvG4jcVjrLRR8AYGrZxOkYATXWKJRGlP78ZyOC8L1XgblYvZZ3yYK8y+qKn
Pgs+EXtL6W6LTderkk9TBHrUfZ2RwjkxVcr2PpbAbdVAh7T/rdTQd7xqq6Mnslxt
6oETs53fuIH0vWkvDrJOG91Yr0P9SnSVWw/4psjoyxlMR++tEFtHgd+/ruHZA84a
G055hi6sJ+Fderm7qT95zY838LIzzwDjNkc7y5fFWRCPkW0FkONt9qWukO8IwCKf
NPuipXU27I+0FNnW8EpDUdoGXVxDlbYiZprXpHcLRmA1uEpH/r/RzA7VpzyiTWSW
k9clE3KkJaw+uzapKkY6oEt+0x5uLxb1he+aGP/8OIEXKNjv3bAXPJhUBOFB7V9d
tdCc2hPuw0GGClVKgCZ9m0WHdKhCu+bZB9aZDR8lCuG1SSljxy0t7gTAdJyighjD
jIqFf2uqKDhsfHamcjocb5pENT5PkBYIu4E8enBNa18eSrIhc4CTq11OMASvRrqV
6As6zGDYJiS8af5TCPqbFOj5W6BfrXT4MbKZU+furi4u3AF9if0esfpyeSD8lC30
53C+QmJ21U8+hN3Tne0lkuhSRDzEfQQBrmXiTDIxuJnoW0jdHlhgei9If2Dl9CVd
FUtSv5a/jByVy4pSRjecJCC/xk5yB8+YjgVjYXHcupypvBTbv/8EoGmVVv+Nt8bT
fcuDcx7VmS3WeNITTR8tZPmGm03SWoFe1QNPi64ntlygbOJw4CBOVmcXBJrIiuup
Wk47RO3z4lO5OJtnz3anUwY7s6GNTOFugkXGCYQVgbl9dpMabntvoj/xm1NFQZ3E
AZi8ZryZJVCX0s5pdGUfJvwKvRI+FZfpWKU5uknBFWxr6+ohNdUmJccBfSde5ecX
TQVZQXs60M0tj2ProZf2R6nsmp3dJxU17/oq0JYFfHiGKODSaVLciw0k6X4bxvcu
vN+ooeWAfIG30Ty289VR7XLWGHTrB2O2ERpxAQrr8wwpYt3cnFHWKHp8LMrAMb5T
qFM5d/ACvgwp1J5g8KJWfzQxYJT9dczjNs+2wWCXNK8zjfEwxcLd6J1JdCIwrYwS
vul0RSv261xE+fditp04EPj5GaKgDkvS5FY/2yD4HNj5bYmbbxu7TlsLn0Ehvws2
wo7TMPT+Uv6LLBKwyIMrxHeh+2N6sJz5mPQnQkoLlKk/nydxJbZYQ6y+TsnJv4q8
WhVtCeFfUW+aA6QqnJ39MfKFncSmK/PxabXTk1nz+VVzGuhv+s5RFCRCGzcU5xqO
eV+7hnULtGW5zYQQ6ngpdAu58bKRcR4llz4z/8H5GiCMA9YyZLUnusAW2TiraItp
ycR2tGW9K29OflmkZUrumhOs/x+Z0enj/DahxR36iU8oPokakrlHL8jKgCIpDJBc
cuiVSMMiJOGpszSaXYBAyru3dFQQnPA0LjMxPZ6jHD6pSGMG5OLH0ELettKkIECL
WYQ3w67lb5LbeDIhQo0ZBV+VALdPzlvVtD8FfuBtR7jZX06s7tOkRw5xTP7KQfcL
M+Op1S0Aonhbtw9ijrcvEgi6K755253ejzQ6dhHQbIA7qrVwpUrz8B81Dat+52Wl
e6PEdV2onEEGjlo59ITfyNdV7H8QLb+3OqCQtTac1x3ncEHuEdd4Nvf4j8gq02tW
THuksY8ZMGaHx6lDRJzVXPXijrTELGjmyZVrw4zOjqSgLep08Ksj5E0v06wHgbWD
rOnLq2Z4lSEfskuvNlCyvzKSQuTi4GTQyvEc4THuqrTVLMdyvBd5OGTQbddoN2Ip
JyDrGFoxluCmd2I+hG+P6I4amD+Wq7TezzRb3j3kshoYk3Od1yQFyhJTOrSGNE7a
lBzzRWmOZHQcXdwrlDaoFpI/ieu+kFk8FpHhXFhx8juozLpXDZv34d39WBBiPOcx
yPTDH0npMLmcV5SVaI/jePmJRiT3EDwNxgNes5Lfa3J6Ogym6lQ8M1Eu/4/APiV4
jgIi05vLdj0P4jxzAkKi8epyDtEfVgtmq5rXjqte6+tOxYtJBxZKwe7OElwGCUBk
zYE4CdlZOyyDnmtSmLkP7eYYJPcPwXGsn7IVGGkff/iPE72MDEvdPENldqz2uS0l
e8STbRNq59O3VKIM+7Watg+MSq2/2fZLSmAFH9JSAGsgTaRBd41iJaRH4hmy8KOV
Ntmg/WavQhOTCOveU5JiWuQ6rI2ufdzXkGG6xRb++Gt35W8ORSormEEU/p/oETwO
fb+XpEZxMW150eBAk1JM70UGH286tyrrZ7vnCNbkqmW8JCiwlx8TjR0thnh6CzD5
A6ZwiStqb62bkreUsWdj1e7mZjA2JWlT0kF19Gog4ddwdn0aEiCyKYh6Dsq57YjQ
BbbZEpfCVTTonFl+R5OJHfit8ZLgPiCbu7kU722DjVLAkkJsfmXedeZfYRhNgeio
6CGyqti9rkkE6P06h2BAtgh3V0MDCHMQxF93E4uUWPHID/tkrydNhh2yddsUpzHh
mrfjzqMgoBhLAZxKU4tseb/qvyT4FWWI7k8FnBfSvvuoYOziVaJb1QhIFTmXLD80
K2ptssBdL+Hd2SS1uNEE3e8eQSmXrmzv5YG682dhU234binbGyVwoLBawjH1jx+B
sK5vgt8CnZfLrZXKRsnjylI+3j4dRdnDe6Gwa7fH+SOW/APClgLtwMLclnJSuL8x
XWS4a87Aauh01Y1z52SwecdbiVNxT96Z+o6JfUkPbQBvw4o4XIr0pWuOikIaxpha
ifepTiDiR/NdjYfSx5IGR48hrmdEEDHPLRCJefGOR3reJ8p0UVT1hi3KSm3mq717
fPS7CusXKfqW19kX382RlewF4MDQUIZqgkDRg1ciOrtbkXmXE9CzYlpS4vIjQHaC
rx1hx2weUEGPxZtJv6C+l04GKr3LAo4jeKCpE7ZT1gUPSpQg3hT/tzMbADc5pRfj
6KdP+e1QsC4b60goSxS2vTm/x8tHRIErhCNyv6+pE7tB4hkGveIEurzvw3i/CyZR
qCDivaIkQaHbpDdasl6+otJlr3hAO15T4gPNZC6YXb2iMdj8D88VGKI7Gj7rCl09
VgEtq3Cr4+tU6N2CAkRSiXusbhWtxC9MoNKW84pepuvmVZtPh9wBwklUFu7sPafe
DU6clrYTNyE5eUgD4NDxiFlZUR2YqSwn0NrR7Uj58SdQ+C7vsKxoMk+4haHUPjj1
z8ALSwKa0R1fMCC2uoB9q+MAvK7kL6Xrq5sWemE+WkRzKvydtrxCTKwHv+feNmiw
HrCs0BcwFaFO0BVstzztvkRdooVGHaWw0havaMs0S0fe8D6aX+n97o2gVHRCnv8k
a3f1WN9kZj8V8dhQbWvF/FRYM3cwxdwblBqPm2gAkLjBSmVXubgIKreQhgmlM1wz
gimTJjkeN8g2H+0U8/w6rl0WXR1b+lX7hDHnuo6stas/DxVa9Ul6vTuIz4f3rQRz
IG+XkVtpbmyT6HwLMuqWsRue9qwXSj21D0jY6MMypFjdTvk0oPLddDLc0xVAuRvP
ku93XNXaY7k3b54hRc/tps5T3Np8zU7YKZnsvNGnYkWj7TbL3nvWUh4D55RURA+S
4HdrATBa+FOqpurRCnfh0PzgoOAcgo1I5WYmK0NDQ/xgSogvKT7HcN3AKrvv+dwH
hBa04HgghaYKcab4rDY8t4V5SQt3W2UyIu4pefLpjE6yqKMLQ5nnxRNNaEQqQKDx
+/Y+93COwHhZgqZQvGgfUtMjr3DNfbVyoycc4buOgcE1wKK5HE+aWFrzFFiFZLzL
58LZtvHQJxk0LQV8M9wyBFuzvdoAhEr5cmXj1O0hMn66IOGqB9FVC9+wOjNPwJ43
ixvh1D2JhoHe/PchZCaLTrE7rG1qUtjlFz6t+AHOhQZVPePT10KYcFK/f3mnYC5J
cgCIcpUNSUDY0JwmO0imQOggbfS3aMK7VzzUMEzp/eHRnAtN+8dYVPrD869YJ6ZJ
K2zJNajda0KnX6bZ9lvV20qfZUYzPg/g3smDpbM6+L+yenW5zkmga5lPQ+/oIfjq
DNme7Ee+fJKdFvK8qQYTsbwa4HdU9c5AJUKZ0QKc/iMZ0Kc6ZQg9z3lZwjs8ZDaC
gQIwRIDtVD1khJ3SYMLsq6xomrKp5BMzeFquvGs2/EB5Z4krzFxv8kWUx+aYzJ2a
bxe9lYK2ii+E4HO/6R2b0QFcFhErbfrJSze3I5QbcrHBPyUYAUPSyerciTmr8QVm
ghkU9x6Cawl+NjkJlXkuW5/BLG+UzF7a5hCdWOWXby8ruIx6EtCryv9W1iFK+RfJ
mi9ZCA7efvb/Jkgry2PtDlKUXwJpvyA6iT9o4N+lsUYakFeXUYdCdgvOLpxYPsYc
Az+bz86pTGAHzlc4hnqrPnf0d65HB9R3cRqHLu5/gbl7O632KRwiwuCwcChXTVph
Kf8uNovX6GhMP1sRXZl6H7mNBgLCsyjgZMG/8frkTTNaoez+h5wTgU/7ZEBy8KQX
0iXz78FrugNv7wBO7IXeIXFnNi01zHyrgAsnWLm6k1FeZ1U26cIiMeeqXDXY1w5N
DjevEwDYyjdISLRrHEHQwN6I27uwyXa9D/bwn258UEDhYngOO+CQVaB0b6gl5c8F
nDHSzRgX0bpOHf/iXz88HFIwQLDp6zwPclHzyxZisLLd1FoZlmIM5X3a4FX8kwXb
fiSfmlSr4g7Mv6RCaZnItTJ+7FRpwYvVsBiBWXboiTy6sJ1uwBPsop75uQ3uw88C
q6J2+VyTULkIkrwfdqWAyEKMDCYbLPgejIo3iRZ5eaTXM9SwmRsrxlJkdEFWWMuY
73RICihRd1HSu5pyL/AuTeruPaxEyGgQe9HrAQHf0WFnA9TGc5deLGIXbxmU7iCx
O7Kesnz8azq8fzNnAJTjxpVSiXdpHFyTMVpw8Cb0iifVx4Yr5XjiQ02RWwS2oJXW
NBsQcQRNBPpHMHpviZs3hTudo+rhLMca1chZfXu0S3CY6LV2evqLzPJ6TBvcO8bd
PLc1i7mqP3wnA8pbFja9YRIm1ja//BvyElmTVfjJwaldvb/rBfc84RyNZSFfE/QV
KCqB+llqLifSBgfWUraBam4FPXGOcfNLAfhkeCWycPRK79brIDQyYnbTZ/n2A2Qu
GAHUmD/fRRGkoT9fgs8sS7m2tRadBKu0CRYdms1a51kDY0vFnPsZkkawqyNO2fGH
z+vKhR1B/wC9Ck0jP6ds5A1Lkm1BmrtNos6YwgmA2EKl4gGwoHJyHQoKTPdplVAE
ZDm1KBctBgQZSrwktwvJ6K6b260+P+NxQH/AA/7SrjPH9z+K7wQt6OR43D2+lEca
+E+O8dC9zXedu2jIA1OI2MRzA7u7S/HTDrrT5Gx8wHKi7k9N2PFZgHcSQw1ciVyI
3tVQkIyXe7Ka/t4kXBoTwpee4ljyLSs2piZTnyqyVJ86izYtNwnzc6ft5V1h/oQx
X9msJvpoxBdGl/xyzTPUiZKcoYThGD2C46tijmW9/GmyQk2GJL+4IHPt9KPvNfhl
EC1wbNnZziPqBKhyqxsCjHVhkK1m4OnHfE7mP4tj+Snalo0BPG1/CEZhqbd18KlQ
qhjSnA3fg8HqfIHfg9DRM5oq2kxO2+oi6kKQSpUamA/p1+q8P9akhuiOUqVl599E
TdTaKN84s5Qrtmh+110Cx0Hss6WBKMC2+AtACfEbMZPQE10qshljWf0zy3qQF+8y
YYH9DUuBQO/+gThBco7BPaZqFcsgff/2W/9LwJ7pNIKc1B5MKXh+OBj9CSv1FDLr
fEU8+qa3og/dTKWaVicrevoSwxHpcKyVWGlDXdHNZ6Z7pnu1G2+ff1l+fFw1p7Td
LEDCLM4SjUJspeH0pqxsY0pdRbD76KiQtuNodR7cug08cjehcmU7thX5JuHJ6+lA
/PX/nDYMIBpVPxVMze8W+rakjnD3yjjB1NUB2uLEhs8iaJe9R51dza/EcdQuMSrf
4t+Wv+8Fo3+nZ5tQZ86sYlfnu+qwgZgHCBgBlqWIhKRtVOheG0rcdcBELxqypHLf
h1wwOrKuneSg9GbWfoqkPsNTW8dwxsiG6C59gs6QZ0NxdIGUeUy5FoG1QUR9LghW
aDQHrgK/9I0z1tcwkMOcw0D5jLvxQsEwMxc6NCjk917glm9nH00SlI5nqFjII5mM
QJdJFBtpu9U4Vn/2OqxRmBZYRN/DbBxVCSWr4NXPHX1sCVLK4uEqvdRT6kSzpbUi
uj9sStQettgJlkKIfU+3kb1fcBvIH/f2QxECfAKK9J9vYgMWZQzSUqVbRb0bhyB0
X3f/Ugkt9M9KRCFNJpYaMuAF81T/Bo+HHX6b2Q5Llj9r74qdSkkN0OYZqBG2L+zC
BCS9bZihVRs5vyOyXNANoMX+bcHf34UiDLUy4pWALGvf6M6THRKl2AuAOQrHRb+M
1OFvw8nipard4VcwYf8DOR+K7k05c1Z799EfJF2MjlSGuH+yBgWDUiPQgrpsxJDk
aUtnq4CZGMayQnkWOJNqn9IkqZA8lgfw07pE6ZlgpzPzmJbrcEgDtIWCNjXMVscK
bJQY7fe/c7RvUFMD58+y/m5x8MjTS05CLwYm8oDceW/mMh8qEpYeXk05AQtHFeXr
b5Xk33nUShPa/VCGwh6rrwgLHwk2P1WMk0Sz8vhdzGyliBdozMT9iQEPab5WQ1Ls
haVUyEz7tQPJqOGf1LeRyMIG129OKSVA2D6meKp5Ey3OEj1N4qDWsT72kiHo+a2D
DjEvMf8d1oT/mfyJnohw8JAUocQ/a9HbW3oBXRqEbRtfUCqdW8IEOe4jCAmuCY7Q
j2PiDQIu+94mRmdDzv/tLBFKnKM7KeogbpYL7EX7bVd6rrdySV4tuRLlxkWHfdIQ
CK33Lg5pNuTpZG0l3HMnTF0fu8CcTTFOH7wxglvqsmX/Z3OX6VFCNxFexGU7+mC4
gd4kRD+T6XtnrmGHVXucbRESP5abCQmfKrNtaPqiHmLOUk3wvOT1LwW/b6Ahm7G/
s85P6bJlSovxlRtCyiqbBBt1dxsQAP1vqWJYsp5/mWFRAPhzl+rTdyroRyH0vfse
gPTkR79y3WVCd8CwNCtfJYrB/MYlNicYO9ybSuIysGkw/xCQLYmLQ6yRRZ1pq/be
cIggmi39Un1CLEpqag64yemCkhi9uehIUEc/13h277ZPS6P6uBBuZR3dE4H5q8te
qYi6KIPwuAv7s39o3gi9jMfDLSNnqs5DFJbqEF6TRoEh9mr562scPpP9yGMyAFqQ
2P/2sLpd9rORwDoHhSGLcpJft7eBYK3D0TZy2utW4Qfr78imKSIhyCeMhRG10Ob+
HvkVlSi8/D2tqDWEoGnqZFLqjq8Ng5uteDH5CKgQUSmZSS2r7GqbuPI40lUjaQ2V
o8E6UD5nBEUY6b4nnLpBpvdKKMfcSAtrMZNep2LXacoNcyti2HsUZ2Qdf0onWke4
B/Sv/+mwZNs9rzLPlWQ7WMmR2DHoXy5GAhbc43erLHAchwYGGNeYBDU5AtLkcUrO
xPCitwMNM3NcymBTGrwa1o7CCyKUS/HbmNzjfEChe5+X0le91Puk83A01VWRr0WO
/Ldjb5PvBw/OP+T4uukkjlO0Fcxym24d2TCeet3zvQENpjbup3YYg5uVAFJ49ASp
UelLxpTXnkuEbb2ZN+5yro83+uTkw5ptjN0HEuVAJWtpCmrCqoUie8o9LG7RMH8u
zvEiMCvOb7dowgEXbpRSRfoCIq9oU07bWurCQc6JueQXGf7hrYyvwPwpXZh9v7x0
EpiSNnpfY3WpxFDpTGX74O5oRgepSoo9YHy5v5IxJvxgBXvzUH5hU8aQE1R5kOiC
NYdpEGqrfEnQJ3LZrQ+pVeEydBcMfZ5YaLWNK2Nhhk2IVx7p0VtJv/u1d0o3GFz1
OOtTvnzIAABCUL/bfKuP1OYfQz2O9YnZackaPDkzfXs4M7ln4/y9vEsaXz6IV75T
3izY7+j8pySNFTjOi/g04kAq5706ZpQW4xy6m9POYEBpdRmMr5PwypMtgvQbMhzq
rIq70ItMYBS7TnWh+XmUuQGWW4N5quG7AeSkeJfnLZeFZFcfNqayZAXUNymKfQwI
fXZpgDw7k2ZNxKQpNVbUm2oV7fSe/nIwq+rg+ja7PmPz6DY/LEpVEad1os7/t5nb
La/qjNfAieoGz3o7Xgg245czrUy6hMPeXQyh0hzkzzHEQ4jGR8IEAdlPEb5mkTUM
BD+GY+6/UNzmV5I2ecoMVThPj/GgBOP1jH8iVAUOYH2vqacLKS7KVDikz8qOEmn/
vMjl59SoJ0iQcsPPdZ15cloKLpPfM9zsQXLJtRhy+zM4HMQZNKWSAXjLY7ZFU4gB
w/UQ6D3n3F4M3Rh4KXgTXA4XHS29HNVE+oZHvd8JTCZgdW9UEkXCIH3cJglkk69i
Dut6vXbbP+rHaKoQj6MRqFtaG6t+t+xtRObRbk/8LVsr/CCoMr9fzFw+yU7JnnCJ
VRpYKnUPORez+95y6ufhhM1eQTrR4tYJAqEMo4q+8Lbex5qoOsa3Xy4Ns1uFg78e
zCg8Fyhl06e7q10stJDNWH/LuoS1Hj7VvIqG6T73oyhl0ypEzRD4bKOJHWF2+HQ4
x3NjSGt0gElrTnvVQ8vKdXVM4NzBvoVIxKlRc5FVPiZ2X756FHKbTOSrLkVK9Lg4
UcV5ChX1XSny0AFwicaop4cXNnbKOWfF3UNdwVzssSzkmTDZhkkL5tJCp0W9SaPk
k+48abM9OQfFhMR9YXtb9QuIkHyndBJ+fYq9c22Fe2r3jCa81Pi/hi/gI2S0PixK
tTRagYo2ym4EP6U1O40hc/BmqPNeoTUr81uaCIH2i8NOyIbRYsJ8GroipUMgO2HW
XV/62fINNc/vIL9D7IbdEE51D3HcssdWMmOYNtHMCIMWb/Qd02RQF3kk+En8Xn+F
3UdNOBUYhznc1O8PuSB+tHLC/xQmx4416I2Qct2cErdqjEgaxoPH2gFJC4A9LSki
bK/nOaefADcf4yY634cEsz6M6b/sGJkomHqUroXVp3JW7Pa4MHrN6B6mSJ5q9aqv
u0eJQNnRsz+I3c9935BxjW2BzKqs35/oEOua4IrjiOVrw8NXlFtH8angl+O0mBnr
qWVF+LOOMOwCYNoUxmDjZ6cFZyk/7C2FXDWB/gTzh36ge93lelMN2rEjjWLqnaqA
NwRyj1qQZ4bmIy+gf9QbQXnnTloODCviIGAdNK456sesid+DAeIUuOcz1aIEhK9s
iarGoWnH+iTTRBU0Mgn7zKcTeIDTTDiEZEEc0uyclxAExYpHWpKq8Ug8PxIP7UGF
MJxSHtMQ2f86OvTGBkHPzFgjayxCKK2tWFUUpnwiHiFyPdl6NLuzzK1i3Y9Hf0Jx
e45AEnTiJQ04RnwB7RH6VvMGdD1GNeFs7q7i7Nzm1JZZ1NjIl7Zbs9wyemY+UGiO
osb0dQaDTD3iTSwH8xOd5gEleB2h/uHAEqJvY2ZgdyJ3MAvPu+a9AX2YV2r6fzVC
4pZeFra1yLVWQ8+xD2ckJX1HFE1sv9I0EDvlS58C0yOlKtKAqAH1DVO0pvWuvPOn
2A58YhVOzH2kW6pqgoFd0+f3IMvcDUw/P7kEyDFLYMuQx0mP37ZuyK+brMDeUaQ7
Z1eT68fcjTww+uBuRpaoKeRQTSJbO/Ze5MsRaNtnrt2AgW+mwKDvpn+eaivVuJQ9
xIVRJKr+7KMoZGvLnOfAD/bOLYI9v/XutXdaOpfpWKLTPMpyjiENtEE6mplZMvFw
nJNpAMGo6z1noMpsuJnqxEqva16h34AVYA+yfgrF4KdDWMtXJm8HpNxhQzVkdGnA
fqnd2rwD4bViCjujR/0PdXCImNQbd1F/cwF7U5cUCGt4XBRzwQ9ySGz8xRSKgg/R
zIKeynJYMYpxmu5a7RerZGr8FZF22pkcPdmUzmf0wE2dOeiJE2C6e+hQUlXvpgj0
j9bi0G8LI5ZPHeUGUSEuE4hDEA/ZSrXKMM907s7tInXTIgB/ea0xfwxl5FwpcW7k
oK6Erq44XVeL4um8ra6ZpSnaJlV16P8OPDfb1vQLqqo9BUZOAQdVKykWoVcfQwNX
QIMzDigwGfin0yAnneTd8ehqWVV5ErYDcJSdrs8W+JhTHp4tcsB2O0sGFiBOsCWR
EMUCsSzK2dn6wRrfQElAZzhWBj46QAIdU0jmpFMyX3KsR7ZU7cHpHQBTgLp/zz2G
PlzXQ9Tfn+dEkEDz7ZrVOVT4AQTwlBxuOC9173WQIAMROnnmT5963kM+wnLXukGY
v2PYByCNqJbcD7N7V/YZTJb52nEll7gZZuF891CryUS8EHQNM7npxXSdghJi8PUi
pHBkaNYjOlfSRh0MUbpxWmEIyptYWWHXzcKjV/8+y/yVGrOPAn+IFEgGfsUWhDDO
+/RllUz+A9Ocn3XIxdUv29TLSC2n1asU53pti60pzKZhlVTkF1bKCJxt0M8mFymJ
RMhPIETiod5iUibv18/0x9V9bLslUvoWcKx9rDvEGL9brBpQQ+SitXohps8PHLrB
wA0WHMeYi6h76MKjIN6asP4CJK94i19tI1wJ50U6Pb705uIxvqV8VFmqL1uYimjY
y0fHgaUrLLBf2mWVO4vjSlNeeDAURjmuuMJqvMVcNz8WzgrE75I3NIsPqRKEFfxs
f2NyQVsi0xjRAmUpr1NuD6z56opFfLOffHcrMSaqq2yTNedEMlIjNhv5XmGMhxUS
0A72kKljVlxyNVQjurCdUzO81mwthL0hY9srGYGTtRPdPZpRnkjstKTLpaqaDDPh
uMxtDXNvjaFqIck0k9epW6t1j4ejPR42t6lgQk0OD7NhIOjS5HTI55L8l8HDP1o/
dQgCJIBsaNFWeBxGWPAQctkczf1cd92IXpmf0qiiFWYFLEIuT3LUqZ11jvdhCai7
/XqJvyt8wQjcUB2xwJYkzavzz5tAx5ifcjRZcbDNzR4yx67W3oKHYO4u3oIB6GtF
1TfnIK9oYMdPSVFP0C0jeWLmSyMqhSiL50Btbs62d3/ABQNHI2ympPS5Qj3YwHJR
fLOD4Sc6iae4yHt7VfJPik/ZAEAwVPUX4R3Ufy5n4y1QsnUWWDh1LGDp4+jg+WXh
GTi3gxa7GJ9Zz2Jg1o77FPKyELGrkSxbSmh2uz6qRXkakPOae57/b7hJdDlbZyU+
51b3PEhwtwi5Xg3YBtP8kFWKfMS1F3PN61bP96v2m77UchMGxUDhr/bws7lljd58
4zs3SpJzQXeu+60xVXjXVGRY9J9IgDszY/W/r7Zc6JMHfgpDNI9WUdT0KzgCfR0t
AApSdlhR1kJZifkhtplfbs0ALNA3p26ZNHCbHZsyNQYIBhEDhTnBIG+xr/yh9gIJ
AgX0JtXPU8cNTk/+x7Ji0FL6877NuwiPyDrFtVP/03KsXi4FtzrhiyrSdNsZLZzI
rBbWLlOhe8D/DoodlMc2SnRrCwjNunDaCXRKNNvlyyzA/4qrLOQG0+E1Wx8O+MpF
uvoUo2649pTPCMqro5xeuIN5/mXlbhldygsJGv8RKGH9z/qVPScflUjsqfl+AQNf
z74QHDw3xWGZUK1efZasB8n1Ggkv2AEjp4NItlghXPFfx75dU/gdvZsHeGNsskW/
U1ptDyVb3/KVwhvcOJg0bizxX1GsYdqGTv679e0Ktjg9RmIH4X/maw87Bz1I1pls
EwwTNJTg4tj9xK2EgdqAG2A9iPblMpVIctWq1Y17XNYInFw5DBjH0BKzS+K7xL4o
ZYWlEOkF6mMX2a7IOVdVlYmzwOwEzlBi4VWnGneM6md9gvKgSF2okOq7vz2/+Y7V
0KuNjzR+sWaUW16P2JcOwGZvRnMDqHf9IRS0vClJedNaQIYPWlBMg8u6/k2hQ8CI
rBhg1UbcMa4r1nDyGw0NlMeUE8MJoGYDlXDkwZ76li8Cso1JJsffDFR5hWr729R+
EPXULlpHW+GlS03ZngCg/PPZ066oYVmohRyuMdBld96Hwm9C3fSUASkIuP6BYapr
f6IpwdB4NhuDIw4Nmm+JNQhua4GdZcHtup6vuVdqG5Oj3BeED0D2lSTaTKhR6ypb
7a8riObYfVYEQubo2/3awdoJ6uqbm0ZU+170eAUYhuawaG58w9LvTqruuwAB3W4B
wKihicS2AI/8GoPmB0ozDyN+BGh68P2EOMYMGaNUYfZiDKkdbWGXGnw3G8Fqkzpy
aAXFIvJGYlLXJKCyoVQDcSQkm4pI0Qq2L6rrle2CP0j4a65f4RMK71ANDBBbRZrg
2okRiHbO696PBnwfjIABGHnAcgp5rKJ4QDWLepTc2yjBcqrzgBv6h5NJLu2+hIsX
T6H4vEpbUHLYi7+q3aweNCMsXRaZzuVZzCCiNVijj3tuKvezZ/f9j+o3bqIBoa4h
Y2FMiIVFw4gz2xDZ5Uo4gJejLzdX/5NQaANTz9wDYC6TPVXp9r3bRN1aGdoVoMUZ
C72MxecqapplXUZuzAWBEwdlI2kN8pVtWKAm3PWUHiRsDaZgQnVzvpas+2zCg4FM
czdXNv7GHZmRXb5NhtKKJHnMCj2Idnb1HWfz7yIGMIOD+tg9EP8APSWTa7xnYPbV
DuSrqlBNBfQb5W42aFKKQBDJUC8JOxPnsVJYBWFEhEhVyFglQzDCULZQXTB55obH
wr+Q+CjPi2o235GHF83/sSp5Pl63K/ErvXQpzcHpu5eYRb/iNwaS2hJiD5s3fG6M
Oa5QfdnGJS0zODHJq8UAWI7RrelzD5MxXJHuWiZ8SibNfk1dIib7ia60rnbuDWRk
ozWojDDTBgzU7k2V8oAEIsk8asc7p+ymPlO+Btu4wqvydAYYCf47B6HAyq5tDDI3
1x7CFcovPWYTAZdJrylI4CtYrXfvRt6jUkirydzL5IYj77s/fV3CFdpNBGlu3h5A
Q/vTS6qDiq4C2ied6qQSLLySQayUbqoxgIcN3wOOk6/64dGpVLHlbl0qv/waPDG1
AvelkUO4ax5AFXlUfL53lbd/tEBfkhpQlKDMjr18bbgjVS7a2Msv3FHEzf2sPmfx
a1M5nlScproZxVJ5z91pC8hCbLWYM1kpX1r6fenAKK4Q3qsiEcyct/O9TENneMz9
IvM1BTZQZ19coMKMRGkOhjP/VjYprhIsj21zmjtEwKTAp4f3h4gJxedbiWxSOKas
VNtnfoLiBms5+lMeSRLfs57NhfUiZzvhB995zeDJ2crGW8u3WtGeAeNhAcO1nF23
sk5qK7U/M0/UYfnLkVLwRoszGWOIN+LJuRBT41nZiQqKsYMrN/M9J4y2rnctmKjx
dacLKUA3asrAfZBGSuummq4OuP2uDAyUGLc0LnkrgYstmtJ5eygfl/Sgln/Zwjr6
2gxGsKTfLrgkgJ6V2IUcGGM6u76pYixi/TMGElO4PE8H77w2Kf+Z/VpFoUd8/fOy
1Q/hdKxx/tA/znxbBBMCUxWb/iOKEEMeaiLCgxGFNsIbbVoWI6VbGNe/JYZ/slgL
mffaPiaH3Z19iMTxM6MgX7djk4ykluBm6DTJnvqCYpDHUF1Y7L+fUmUijX8ZCMud
hMtCfyiixoccAqyuotnvXNUIGga5uQgqp65yjBhgBveo/kqdIEiWPPMRmb75H/yl
OytsL+Se1TGYRQ48KG/gR9AGlIE3neiUUp7O3YJAEAadoB8sKIb1ZsSC8Ij1knmG
b7uWw+1oyjqxYUsmOyWVD6CH9FuvsPYxKTtN/DNZbozA4CiKEHrrScQuToi2Omu3
u+5aU/cRspBUtYibinY4lw4/w6ub0qchN9wfKvdXTaqS7/5wio0WKJT0ORoWEst4
h6zSHmh9RwnkCr4lVlPy6kpTJHZF3Qa7pwGorfJeNUGWTyF/Ug40rJfVkY+kyFNB
TD8jYh2OmYM/YVDTpRJQ+SFg312F/+5PQlyKm0OnIAV+UdGcFBfNvEvKKPjI357n
oLknv60A0kHqQmZx6dhWSEk5lH1U2AGWoeYGwqvqEbYs6rQ1O9ityZduUIfM2R8/
4Q4MN6uqg6wX5EWZ0INn0zybATj9MIBklv8OajwDcLU3/FHzglcaQTJyuZ2DyR7v
STdO8aVR92tCtmYWZV+lDjy7m3aFeSvivg7Kb/NXg1PBqu/9EELo3g97OjgC8/IX
o1nD95f+qLm6nrfZGWwpYMfAmAJ7/nkwst9V5HLZ1O6nombBMt5+9Fu72x1yWBGo
CZVQdwMzH6KqknXwEq3KLCbUKKisEt/xGVydjXizIERu+G+UNx8BtL/6gaqzgt3b
dSsGA/lw3xHSBeUmttyEx25WYW67Ae9jz6qikXxaSMM8lYc8nufHNydVI4a5Lpzk
QdZH9jxegzcUYtAz3J1OXh52e+hzE5Jz42hsMeC8cJf996CTFlbejE615f2nU6K5
qo3DoOU96AeN07n2Y8XRMIlkznIYe8cXW2FDM63C+Oyo6ahIq/m4cYapW+GOfjxg
LJI/zL8+D22F6b3EaD5J5yOzl9OuAT6WRDs0c1SNcXW95Q2FzJ54vnM089cnewNz
HWqTJ4QTc2M5qJzvyMURWLXzJkaxjl55zoLTdVPBz67EG+PdUScUAWsU/ql1z15/
fciQ9hnf4LRYUC0UYjDEXx5vPIvzC8jRIgcldpxZHibqCE333ESMsTLS//EmG2z1
B6l2gS/COcOhMHkwQJb7mmr+KytoES8mPLfs+1eAnkwOyqqDl3vizyuO9eMXHOKD
rZlicmwajPHjvqiHeZEerp650FRF5VhweHQvbLqgYk0W3fkggjIsS7kpRad61GoP
zxu8TnZMBvul1XrBJm8GUEV5aWqF9AI7x1Pjw1BQbIe7XYZ7kWFKvI3jypnmJf+T
bgRtM3Yv6gkRM9JQ4/Diah666rFbcCYamvItyPa3Ixsv/5gJcqm1NbDTLWsmHbw/
lNkKm5RChc/Fb8s5Hg7Wuyil4UTKzRCH1rqv4wqORJ2RYZ3FNJEz4qXc5toYWi2M
IsHi8vuyFdz6eXJtBdY/XRz1vw0zWUa5bx/cUycMIq5RBIltm0JfpCfd9HZMKjyL
E67AvwlRmb0PYDp7bLHbYJZtfdc0xl60YS9qL75ItSAfNBgxYr+TbgEIKeE3qh/1
MBjen4+MtKRdth8WR4xgflC3Rrbxn9ydbYHhLN+cmF1DJSE1Kc5weitzxokV9TJj
SI6Fy7F0bnNwEYxK+c8sBBUGyDFia1w9e2b0zDBXhxe0Q60cEt3905D4PgdRu56m
UXkXS3D+NgSZoJpwUVyhPFSO/UQ8CwiIbUO9uQsSFaSXQ4NJEPFJQO2mSrb83dqT
hJBj8KQyIb/duemObrMm25/987NQ+TiuwRfJcCAVY8okK4UeqrQK/PpPsKoNCBhs
Af2ujwuxqLAv5Rpw3zVLDxWHP+heb0VCc3qr5OwaqBtnxeYDnmM3Dw6gmR6EIGA+
O22EXAjLLFO67qEaDA/O4asqhhUo4BTbZ1W250w09+Okg8NFlOHqjPj/z2eoOVc4
x04DMOvvcXZu6y7Yj+D7006lHc4NN0fYc1BaqJIzxB1IuS3AFmAIAgdaSY81knym
29rh8Jiir6IEvQW0Ziq0pw04hAvTsnZ3HMe53W5v0XVUrfejWqer9Rqxc6qv2RF4
Mz7Ijfu8dYQ5opDuH49F0popZWgCu3rGo+X2PYrHuI3qnICmwXs5NGJw75phTj5w
weX2e+lxWddjLgZRv+Kq0y+IsuxiOkyeC8IPHCSLYbAWOgqrZsUZUFRxJ72tVsbN
g6oHfroYNYRV+oXBMab2yxdS3bPeCiUrsesCGBpq6lbOS+lXwxzoAAHxAvf+zC/o
wuBgomA6X1eeEygJ2gx6TxjlCoaBjoH8wlUosid4+tTGqPr8+GMFhB5o/xsiPyy3
81AjKba2s74ZQ2uKX7t5LOfMQdPohposNlatcZuf5sueO8dIDH0RploWYEFEADXg
CWwDqM1IiVq76XVC8gLSTf9qCZYj99EO7eQRczxGRE814SdD32Z7O9i2Vk9mh+tU
R0d6eQ0v7DjXGeyP99sMiBu6gPRN5vWMscei2DFWoWl9sLOFPhQRGmjkKkcI5WLN
Io6DHgCFnafhCar4k+rbSkHUnHKIbSEszJzIaxsU9VCK0DjFcgACz201kYwml+/W
glbJQwjRBITCox551c2zXJT9mdbDBKUQ2AbXXVOFst0v77vOcLFrbVbTj4u7fmmz
ZMioTkQSZ5Cr0PfSxPVhIXSzI3dsHF+xPWqCAUPVqSiH0AIYdPYjCw3uutPgP5Rw
yr8iHSsgYHrKBuY+UQEhi7jcr6f+aWsvkVTFEClXHrWqUMlMbSnGoZup2nXjJp92
38Q5QQLCyXt8pmCPljQQNkYk3qOPC+BRVWrkR4b66uAtrqS0Dws1zq3croupK3bk
lIRvEB8RmrwHtQj3iFlWfsLVJfwOyEbs2t09alK9iwFudw8EnlOdNEMFiuJ3BELQ
7rSOyqtvLGl6kuy5Atbnyw+9fHKzH+rp0Qir9FSdOwt0r1bU6VlUHrX/R+E23Icb
nHUYkEcBn35XjEkw8tjQULaeBkPLCJpzZVR/C/ErsmE1wL9+d1Ut1qplXpu/MaYR
tuT4/5v8jh2pKMYXe8FnQUPhIEdBwVY62LMpuzvXiAnFJ/jQh+pGXbLG+BTbZd2s
ZptmeE7ewkUOBkDPqEJ7XkpR8YZmtddh0+NgnWkaNjyCAOZYzOUR2lIRkfkjQ+u8
pn7BEToVz0eJsRtq1F1GPOj/eCXZq6BzC/FGralicRFxxOnE7pdwTsL79h7o5qyY
BcI7PMpMSV/lJlvmHR3XTlKczbN2iWr2HkTHxZEGVrE7uAWPZS35jotRWKzAxJrS
OYGoZJ2eYSVyWfV0WoqhFfmTGTZt7zCp5WHtV0F+woXAzqxie6lSvMXLs1MSgMOc
+VgAIncFe7uuzJwhYzZM5ZqI6aCG0vIsfvLbthJNudM7UxO3wnOdM2mNOdzYAyj9
a3/CoBkmN1tm31xI2dhu6l4C+UwyKhDGwdqjPnbkqnKc5BZJ7HaJ81LzNCfdlnI8
nw7NblLZ/NJ89aZR39DfqVaMSrr3atPjFVkUGr3JnlOtb/cAMIfGl+PTRgE7lOli
mOq5w2VBGyyFeYJ+mLMPMGDDfVldVB/NyaeK3WgjTLU1A4dWAym+OgbqBfgvrRvU
ADyw58laW1KPtbJRovPinsqTV/xI9sNJ1XXWVwauM04SCN/R6TGTXORIP5G9z8cb
bvRO17SKHxBuSD/mV+bp8pCG9doTtNwvKL0/wTF8VHLZ97W8oWCgQNel3183A06i
bQ4t9HiCQS3K+LE1H2O6lVc/MOPjdbbVyzexmDsxHBxLU52DQp1hJcnkDiITCdAR
7lIXMsBHyDDtnTJwhWUbdH+E4PbrUE5o52FE7uuobd6paT4prlWwtOroBQeq3b0d
NptdKwk6Bpr8ZOr/HRVzrQhy8ZvEZR7prgvaQFrrtADIYZzwzkUGFTar98M8NCJY
i0LGDc3J7orZTvUkUuYQix0E0HVliDOH5LIMoVgNb3p0du1LF2gx4MVBparXGKNq
BZSFRCHckD7A/nSTXYc7iJzT3wkevOXua5gTkGip0+hX7kcSq1YFQTBthMsqZXyN
letPnSaqtQj5VTV3cHnVFEK7J3lzAwyl5jI8HO/y3pgjVbaU3frCGFyTcJW8ge6w
TmtIAOj0mpbtURUE1hYx4ma/Bb5AnQ4eAnJ2mRZQZjtUJvY+UimY8luDmOFZxEXy
sW7ztXMz8WMeselBxKH/sAx8iece8MYqQFBIZ3hXxqYQCg3iVdd4mR5AlFd/iRbM
ZMfXLMojPLCBCRuhiuo31SW7ta6UZy8NEgShzgmhFtXAlTtLQC5Mw1B9dN4y8j4t
m+nqkHQSu7psPz+f8iRpKzcr7kB+5FyU6E1pWZUVuatNx6oHEQnAXICt6LhJylxX
lPm16PlLoUy5hcbWa1mTTLmQR3YucKvGH3pvhbXMHIrvXwGTlwt70bjW1PvnGclA
bzcpcxkYz8KvQNZ9yLljKq5teelTd3PBbDk34MhsinpyGa9hyv1n8MNn3A1U86qV
fXXxb4ogUzm0uQU97Bt9mIOm4l2lEx8zfVlvGU/clUKXoRcV8wwQvrQr9JKddfvP
Sr+yzdZqoMKqLtlgK/0WDCAQuCt7EAxM81Lfr6I2LWNF57wwQ6crXu5/ZIKAEfP5
mn/no5H7TE9b7VRgsJV/1Qx8iDt5YJU03c130I6+77AWajdogYh/xAEgUIm1HhVq
xc5TkxTTF8f0VcwRnrGbEDIYaiSm40UkERB+h74RZ5z+SA6ATDwBURm/QqLal0xI
L6I/XzT1kAJd94y0+nPvvKzDdt0yUUvzWddUtPC0QVe4r9hF/S5Vx48pzVJFnezF
b2e24Ph7CnqB06FQ/r2AL1tCk13sGQnSiWOjxE3SZSGFwZgrvvIKmnBvVEfE7ZFe
O1Z/8/QKJHB+m1Y9ofw22Q+E0NXv3R5sxos6VRKQgob+zDvsMpFNwfrCPG8PG3YL
hUhKY1u3iY0IAk8ggftxOTJHul4F3MxnQ5HrsKcRJn8=
`pragma protect end_protected
