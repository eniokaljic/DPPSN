// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bIgiQdm692fdYBbnwHnx9FKeYM4TiD7pfrT+zuAeJR0WJHeNzism5bt382hgjkBb
sVVPU3ej5udkUX9dRGKZJGFJOqlx8PD5gKyV4WnEixOUgYsVqjow97wOhjeDezxP
LqN5Xz6Ug/sLfpwiPl2uwTb7PeKXA1JGQsnzQwP42y8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18352)
ACWm96hHw3GDoC8fFRCk3gtJ1KoknEw3Xi3WnFRz1EKvJynmWE1bBAuKoiGMLYf5
gTpqj8cGQDB0zJ+hDbvmztmzQZl+w33i9LjDJUqurDIytRyz9Ngm8TUFJKairErq
hCEoovfWA930A8GyUPjMX3C8gllNm1qknMuLBBI7q6bapwbM11qj0rypq/Rag+gv
Nvw1jB0uE3tXePehV7/5G1CWr/I8pcHnCgsSrxqjuCOce1omLiBGqau1jVXKfovW
LOTIyF2GSFqx9pD01hUX/bTrMuATzJeBFYJ/6Ph06ZWZtXRlTyQacGt9XQDk6D/w
xj20/jtxotfgNBALleYhzwwkXJMz9dQhcGlRKWICx4NMfXLQtSirKRgZ88WJ5qs4
9PcUIfnWq50w7sR/hxniVJDNNVm+VSw6TSnl5/solO1A4ssv5Ozp6mlFr6b9v8e6
E0RQDKCmrq1bEmLSa3LW3wRUHNMqXPC90Faxih9Kf9PVaKU6KRicuaiTBpsKQfIY
NXi9Ama1NwV2E8yZEhs0++oTzr9uhvWViV+BBTOzN9D7eKFiFJcmRkyfVNxBMqaS
dwnEYR1HZapejQbYI6GMS+n83hqlt3d/XbqKvXwUubQ4KZMiWaemWYrAFx0lbwvp
yGFKIhpISN35TAaulBX470ZO5So+svTjakkrN7+V6SodyGG9iLUAaQbDj7vZsRki
I6vezoCbjtAOm7uWyEoVACEvgetkDpz0hxmJiC75PLh872xvP00AQ0dnOTHmeDSf
9sZxbpXV2F0RgdvWm3CeKBVg2r7TcqdoU10Hn9gtaOSZdqL3V6/bkAt+34ncKSPQ
AKhCQ/eveuttEMD9ujNoIxv3592G6NrlcLSIesWQWFsIMPhoEJ6gvriAEGITyjUx
WuYYjyucqljWSmqN5uO0NRn3IWEhnsyQKovmfG49MJ2+6qd6NRR06WFEYxIf//8L
4l83bqfb480ONINIEPYysE7qLrShNj5G58/csOeYlIdFZwkKVXQlwUKle1qrVs+q
/FKVJ3u9GD0GFvmoU9MySID225mZhUVvIRaoAFbC0QhkvKsRlD6aRNKVuFdbE/JF
BdH6SOp/yS2k7YW197mH+6tuc6Nc1YDIr7nmS4DAWSP6KN1MYMQGtqnnISDB0k+o
qF0sylah/Q+pwG/iXNcG0lG3OYGJUEeoaF0UOW03NaGwKIHyxYd3LGpyUc0TKuAo
ZFnFq4YBshKK2odiluZO2qDAcXu6NoO7sL5nbSWUfqyEwxZ0iqHzDBFKpaZfXMcS
0dL3d3667F3HhXHD5Qzu0CetOLRMpJxWgWgDwXHruJBgO/S68bcj79eqnU51XHv4
5it3iQbbs+wA97nVBFj2Y8aQfAfzQvSZf/Wv8dW5/CarAujTvjtIE9KWeaoTujDZ
8auEm2wQMKmxLgPzkmtRCy5nsYzC46nrF1HRZq9EZ7kceHNmBDK6klH4ZQVYpQt0
OzLeP4tRQq/DB5BTnq2HbZj4bl2LuWXVrQz0Q2+BEJQKk27L1Ys40kafdHwE75u5
eKcAc5+3T4fvCCOe+Uf9gSTDL26LGe3vo2Mi8SR7+F8UzCw2KabcrjmhsVg3Uo0K
gd/7umtoasjIwrfcUNciXhUNjKjRJ4Uls3SYmtuEYJtIgoK88Z+HJ5tztPhfhmj1
RQKgY7wEM4qDUXyIILbzHgnsMTRVBG6RnBbegHjD3z993fCcrL6VrD9sjImjCUaH
qhfBnaCNrgACH8CYtHg4Vw1/iiOJJB2mmU4Sg0DRb0ziK44U1Dep2zipvuSwzW/K
5dYVQAkq1qCGYDrgVw8QDompmFFxms2LGFJmzxbkPHSuYMJc/a8Nwo/rg1F0+cSb
PENCgruC27UxOXZzb1jECvwNF05GsSCiH1/OUIDQCL97yvNaRaBMTLPyhilJwDz6
JF9EYCQ0388HxI9pTrydyiNcKeWK6Xkd9LPSlCEkEBBXTjfAlBqoUqPh4n/dRK2w
cmnECZTD7MBpcw1TVg6tdlTIMBYqqIjSvy972KYGWdlMmmDK6fG7OD8E//NjDvQP
XPK6Qxh1jAdxG0BU8rCRS3OPRtDcSiEmFSfaYH5wsiLkMEcGogJoMdDO76DFWMNl
rZXeNCm6GNEZ6BJxyo7Mf4mlnVpyp4/Rqrt8cG98NQthr/rKOEEOlRKT+DHMEnEb
8rpWegIT61Su0QhWXB5WFiDLeL/zLxXwADhNEjcKD2kwQOnCV/R6/ltkz4O22WXG
oZNVoff36LOMTMCPLztuo+uQ/eyUrcpCRkWILTqMrlm03HR75bdiPw5Dy7KWKpZU
FY/hwY35Qn0vcr3W/73MHgPZsXKlnMUDMmfgRhTjiq0w/jvEQMdEJ9MYbZKu5sUQ
pa7AxMXWKE8LpFIt9aThhnqog1mEjQixBbI4aiiC6GpxsCAIYCZS3BP3tZQDkr0j
B7tUebR2hG8ZfBfFRTEeKzo2AoJgEliBC4Mo+DDlPGG2p+O28vZsTV32E03mfrTp
4vgB0V8tX32WDIa2pgW9698qzMozPYY1onoX3S+TdDWJ6wNlRmGGMjxGpiRrXhlr
OsvsaACj6MiYZDlX5nYzZfv8zGSNaKIMAjZhWz4SpAMjHtZrMMplqGc+rsg1cM5x
SY1s9bvcPnFP0PwViW4VHLQZxZLOQpEeLHCXFFRQcvMpTT2WohBuLnZ8AotpCQLb
qjjQ+aqp75du8qYvP73Cd1zLb+caMgKaWiskr/PcGKWImWv1iOTdPnRLcSz83MWS
L2QuzLynEkvph/MqdC3+8MgmgIopTqgLXuYEwuwYb+hWxqdEOtPPSvaEedbb8Ymh
nT90wcy7sPkH07wkyde43jO9vt7VoilHOlghvna3NnQQFn3xAAzoSJURrT8INtHW
K3VPORE3oRWvA+xXlHqEPxdbUl55Taj5mranlN00bWkiiYb5rlDGheeWtKisjfAp
ZD0Vlzj40QbS/0jJ/7Xlkw5uTwMJk6+MBMgO7gqRwU+dS6U43v8MoKFkJlbpyPFr
iIhlN4yD+rrwM/RnmSXjbIjLjorfsDBmL1gkDtGomT/bbL2cznKCkRfwJldu+gak
Z/4DwHYE9y9pxMhmfz3AjzjLGnJMYQMPhwrj1TOL1f3QVCvwSiX7cuUGm/eMyWcX
qslpl1efTHvgEwxP6pcF6l6C26BitqTDR6pM9r9iS2DLCkdwbJsS7yRh67TNrUFp
BpMQjxvVladbLH8eWWaWHB5aLpNrbNMNtKgK+mn71u6J9hUpiy66ErTVBzW9b1xc
MvbxlkFC4xo4+6SJ3GnEKE8j7huPd+aJN/BohBNf7y9BCuglV5UyCucPADc4C5DT
6+OarALMwd7d1Lg/4E8uwMH5qa+Hlg0RW4f6J4x9YGr2OV2NgXyL9dRhevq/0BbW
lu6NIKi3r8EAYjjwHd6r5xEAXhetZ1Njl7GJiIYXMAuSNDt+CVm9BMPpzXX8FGwO
3K1hzsJxCDlVSi2oxs6XDNMTP94JWT5DT1H2D5aHV6LmqKZsbXV1uuad6KBmWsdu
eaqVCO3YfBrG47E9nHTsKoUBvbrRwcHF+h/zjYJ98u4IxUZTE1AerVtZdgw6k+S/
IZUgkN7j5n0Rj9+DLDRrHstCUVdyj6I3GfmecKxVJigqvUIB5k+xn6Q0iWH33gwc
kqtuoLdG6lsjbb8oPzPpRFHXFrLam5/SoJEs+UXbQaPgZUr27Ct9jLcbunwN1Qom
yVl82JmBNFGOEN8+H3lQuDV9ZdXLnNC2+GS1nOm1rgv2UNeJ3vGkZLt3k9oo6A3l
WGM0e7dZBMv/XHqEetXi95+KAxmqwVouS8JfwuLAAcy9R65WO/RBCuzLWj4ZAFhR
ng6p/94I6ZsqhGAcTiNCkNNAjkUywpw98StY8Nk62+D8p7XlarzGNfTWeb3mXMTZ
Cux41cTphWChJWdzONsGgfACzab7V4Sg533DKL/LRW9ksiPFuJPoyJPcVQjlzNFQ
bMXS/Z9iZB/fWWRC5JODkYHRteEgsoa3U4I1/t1EM8aaEuWI8aLR6ULIohMH+rhU
samKefrktKNSE8qRRDGQeQERtZcHrsdpIIGKfPyh5FxVJe5OO25ualintcRC+zFW
Ss+8EMRdAFqGo54OwcijfaXMbbb4zSeZtL3cAMJObvalVyN7Rlx+xi5duRYrx1BI
25Ss+7y81n0XXvE3JPtPTvRNKGswY+DDRDgmGTNkXZT7wpzM+0/7TpemHv7XPRX6
dZ5Qf9RFNUT2iUI46b2QBImmdRij8wfKCJijZ+lUuS5zcuQRI+9RnLdJPEWIz/3E
KPZOzv3GRGy9WRn852xqJX5M4X1l9t0JJ7PWh5TsIanBKS0IRO6rc/TdkhD8sQ+A
nhFjL/cod6+D74CdA3xMPe7pznbPGtsD7rOjb1x44B0SktBV4p585EeHaduSEURb
Nb1n3hbrF3o3QMIdb8CnR6SaP3fVFv+Lh0gBFtBfoiVRm65HG+QIvwDGmKD3ZCWO
b+VVyw/TTJ0whcjSRxAAZxvw8Z+RnzJpMaQbKgU2wWV4Yy5H6mnF8xFhzJbwR5Ro
PLtlEUmczgyYAtEJiG7ig4NYnmLwkxCe0jQAR1BQf8DlZH/KRhmxWMJ7WvHgrTRO
sk2XjgrhFJr3Na+ywFBD6m3lfFzwOtjOEux9LyaGUma5yiHYm+FUgkkqmEHkeRmG
laMMiThMDmcJhLxHtMxy6358FZZaeKXFFN1Gc7TniJoC3rOOFuJs9oyJNOfChEsK
UWK9TCxjY576/dLG/tUqkBaFA9w+TEw5fL5AOf4aCQ0mOi+1P1xRCBfGU0jhURIF
7LiNw0uYgCdBw/IxHRmDZMD11YcwuTxhw6zYOvZB3dKowHV4SYfkY0Tl79jfTLxt
EVZ+mTxfFeGlHx9ulKjFtMra5cV3ihGdyasoBrDoKh1y0yzc2T2taHXYAcS2rlKV
PjdmTi4a88uTKAPTht8OLSVaJP+KbQDDAFaIGJA748KRqxNVzPG188S/0CqtZ2RA
ceLjgkAAhu8Zk4TJf5w/Z/g3Efjl8emKIKMZ/izDQFnhOTDv6sjIDR2h4Mvc0e5F
gO7F3tizjCeW25V6557YbdeqAVDcZt3OsUGTabEAj4hYsQcrwEm3BCiOQUOXOPBE
XcShFHEF+lse2kxhirDOfHuEli6ERX+A/LdM9UGjx4GeyufVJNS9+yjEeyU7v5Ul
sN/Dwmn0drRmO8/7bU3LhExuZXaNfIr4spVn3g6l7IlByWKMUna7c4XW6LzCUN4r
4R6kHpmKnDlMay3CF6RUFLjEf1MOblInlc+JtxAYi+MjMJoujbxCAP9sfW5h7+rl
ERhdpOxkr6manglq1Un2MRKwMOrrzE5n2++un5LfdAwDgmQgc0RYo8d+Jyc0yYkf
9NtY20tD/dUtlSFugKIbnyweJyt2l5nkpdclj+qjrtPItyfYt7YVtIOcdpruTvsR
MFyjwJ41y+TUcfwBx+AVrYk9Y4nxRIplkiKxYglieTRrA7C7Cp/zXzCt0ZUStxgH
oNXuwxOcfiSZPwowvdy84VRWFfSFYRC1w0oeYmT0922YyRoBxpWW3/+a2Z7ws0Y2
40sCq0O133o40DImMveWQcKxkUbpcwsgoK8XAcDnavdpXh5DQLTsjAYb2+ejVjdn
3CaTAL7/b7JghHTli9T06ot9VWnIL+1OkKm8hsjC88EGOyped4WFUEq14vvXtBhY
f1nMstWLQZG1t2P5KEoTVOSND5xua8bA4kRffhMRo5FQxWxmdwtEZNe8eK5PCn5q
wQ631raRiWeKmwv8LneijPoJXIF1jYshUnmugHOpfCosisgLdDdWQIy/UhEG8nAz
la4J1ga+RvUGxkY16KlsRfUOryHGMD3FMoAgOH/XbUNBDySdiV+5lMJDpfqAtgra
k5JEO2hDxyrcPGwB7FPRcq8ZmB/v2IBtIeqRNGsB1y0h/QdI5n6yas8BKN3K6YO0
KuTOsnyyp5VQoeRZ4gygVhF06zuNKGUyt26t02VB4W0o7JpxS5QqGk9rXFeQ2x+S
J8YnKBI9WQD5XeJ6G1iTI8WBOYH+RBbhObQu/LRUuWwIAOiq4FY9nO6syD5cCHfe
59icW58DxXecE/iPzwapZCxva+4EBOkdjmYZf4YXqRtPY9VrPmdfF9CUybUO1kZa
yMsL76jiBzS90FFjgd0WFs7KIrqOkS8OGcth7Vblm57jBE3JPf/ol6BfToprCMHF
WOQYpps7fX3rLh6jkRlo1qQNoL88DSEXZZ186VoCnl6StmIKUYq0i0gCPE8lnFeM
JzvW9rTVbvVdaw0qjQr69HBWYqfofKSHDcAuqDjOaaaC3nrfHrxHa8whKG9R1/CS
8JKJEObYZ84DnGOenoi16rIi5i5b6+Ak2d0TV7JZhiVWOQg4caOqsTR47TgJKu2i
nML2Izj584Rg8CRlIDlipqcxXAjSoFMWpkiI2B0ynZ945V0zVSrK2/BQ61EsGny6
tDcNCs6f76y/QF09JTYTeaqwveIlj4hDN38VQkd+OFgL6yg7gzGQhXh7f3x4EVz/
nmkzuboHqOxqGXLHOFEL30RdOjQY47p1BzFrDrCZJ+Tw2AfMIcOZa6Dx+E45Qs91
rgyEzOBhIuQd3PcuhbGqAA5WpYO8jV47Uum/ajnWFYPKK9TID9nZHYlMLl2TeLKe
q1TkBVcldSi8tnyblp8dwlSFvWI0c8ehlSHPekwN62tn3IfM/rTMsT1Z9cH2HIGi
7chVxWAH5XHI1ByMi/XpUXapOk5dSELAhrY0Tvz9cZsYO8Ycy3F1WzDThVWyo8nZ
heL6WZyKT/XAQtI/N2mInoW2rfYZ5o9xVdu2ydDqgzk0E0gDsm9zcxVNWK+KBowF
e8MzhC8oUW/rra+cziUzk+rZiZ3Ta3SnbsCuS2agf2eoA0jyeNQPTw8HwUNu1FpU
04JTOIUU4ZYylPBYjxkD+vyLZnTogbVVnjUFX+KL885jHw7XnnR4I4ZiTH+i9Q+u
xnuwntRTzcAGlEsD5xpO9AYQiTavFvGbK5PE39Bt6PONk/dy+m+wyMc6JJyKJnvG
g3hIFUXxmz88hiPhJL2i/m0Jt0JiZmj3m6bjQcbRZ/6qwIBZIh7qnzaM+A4hfZ7a
4vTlJ0d3bD4TzI1OsD9WN5TUNOyMBIL/2ouhERIIS+SFijWSXzRygveK/0duA+P5
8JbEakfNGLks45zO/mxc9mAEzGr58hpsfDQqAsxeNT1Q6Gryh5sSSK4vETZuD/SO
mFz4Mbd+nzVku2C2HpNsdzHFX0Jy9pooA2ATlhKLQiXw94bhdsOBlylEhmeHzPGo
CpDsde7VcJCP9zMq+pGLaqn2F+aZYsDguagiF1f1WSbMENOCRQwcujsZVm3lrWb2
6EfYdRC+S70hfP6Ylc7fTp+D7mf5I0CUkBinC49z2cgEO0vXKnPBjUKjpQPcMbp8
UO2WG7eJtCa0IWN04TtuJ+2hOjO5z9vzT/I//Nflnnq13FOxj6bHeehzEtl7Knge
d8qKpPAKaWaIJtzHhRqVklYaJbjLD1uq7IwXtfYzDry6H1LL3wBCL8Xnl47hRxOV
xfJdAEq62EoctYu23yrKWjHcQUNfxV8/og0hu6YhhF5SoqiZI4vQf/vCLd7Uemwc
zJeA6aDvXzB+SnU9/FI16XHojbvlOmy0KjaFvQJZB5YB60P8IRDy/3Ze0L68Evu3
Wt8adT2T/humWo+MufgjlboumfCWoGgW+dITjGfNRZTmQ9pk4qYErFJDgDQFwHwR
YEGdbDgngrygehcundILZDmzN71rOSCifXxpPuGXBmyBind/9ekb4RzGLO5MDBRs
4tiyRFCFUlHQscPq0JoayFRRG2KU9dOT8sp0MQWBLY+JcHhaXecXUcPrx0CTMU27
61P5kHEHY6TpE4pdL4hUuDJi1r+ihdHRJOW2atyct2oKcYS6Oz7Hv5pen7YuSqIQ
YFHmucnE5+p1AviqEiXHDFfO7SBLUC/mhK39UZuFY6FvU1ykXyPL99L3k9pypPpY
dNNrhTiDlhlpMGSjJftrR0nbq2qXuq4ciOCxQg8fsZPI72xcvCVpiiK5k7z5NrjH
Hu2V6EljR08i6liCIT5uZXyW/nWkJZpBRZ6LMfcxaY3MhYvXtNqDhk+kB7lZDdrB
lh96rvgAlmqie/kIljl0JZQ85NMTqXGA3/ISivkH7c94BXfMlqrT0cRGDvgXNqPT
za77NW4aIcsiJ3ikgIQW2Py+2iVhwlx6z5El3owtz6iR7cgI8fK0m2VLWWSWxBqY
g4DGyduq/RWc9evueGG537yYwbzw1iMCBUdFOox7uKBeBMZqQyDo6vHgKkHWdrbc
xgpfssySYeVWth8wEbdtm5/y71AGYhHNJJo+pAVbNHTcifNNZGCc35abJEdaveTn
vvLBksDNlVXwDNsClGfabFuOYXrHZGuh897kKDWBRhh1Bxn5XSNqj17GfSvak93z
DYuHeGI2S/6yMeY4QGEClOGiqn5D3W6CTL1DfwwyitXiJJ+NSjGcZ9olOJ2C48Wr
pIAadCj+daFcDgPKdY4/yNtWD6h3+Cu4o56illmAN5P+rZklulqU3ahsbiNWjHWV
JSPB0klJwwamGEahbtKBn3IAbWXsr1JBUKACl8czKqy4uRJIbzI+r9F3EoLMPNMK
PWTnCo3xHVRQ3EFHyxFl30llZgO8ldwAwtfBTivO0YitbThTCeMdGCywqrUsz4UL
1uNgJqhgtMg5XfjDxQ0enguS7MXRShTSVKoy4q+IPqleqlD+He+zHdvitgk/reBp
rB9hefjzA8VUP2Lh6lOFPvJtArFyJuxdv1OHF/ij2qAZM5prGA2NJ9tgIFpk884X
QWSruFpvAm4+QjJNwwvw3JX7/6uVXKGNHgqZ/WIsY4R0DSd8/bp7DWnjLYlURiPf
2rzJiIvilLR9AjHrsOmdsrARfZaiXhFPbJ5XM4hkC8hUHfXiBPotn9gpmgEDPxY4
Uf/8U4NxVOWOPV5CHZZtWRTgeDKqGXRDZke7EImi3gYhyLmkQRnWaStQO+NRuewP
oMqIRlZnKenunvAoo3Q7dw74TWxBSqIVNE/pH/MeA9JIGXNSpHhuK/iB+67G6goi
DGzZODCTGBrrgoFasHjqDSXpaxwNXxmb5KPtACuU3/Eg+fJS2Cycki4Dn58uvxaI
FeVAT1xguBu5N0WTle6JjBpgLwoJfnIUFIjm9DPC1JK8pukQuZANZryt7F/0BRa7
ubvTwSjduqXn0CphIW5CgQYEq+sqqub5wFVJBGYTfTHyOT7j0jYL0FlPTQCpffHw
7bo4MzAEwC01sxurYAJCpdQT2jcHLeCzTk1S746tkqFnTDgekTka0MySiUDkWjSS
UDSHlVesiud0kypvdI0q+NgZx7AIA/9D+h7heT9ryQ139vK2XZFuZV0IXgmOFKuY
wrGInGRc6ZNeSYq1NZcZwY/31DEmDMvhHG18TRtGOjk6+9l+cMXSESqnpFNJH/UH
zvW5R6h8wchGD8ZrfmpUh9QS1CnvXfur2kxtzInB4vvR/HWmGY55mNVEfhFTwc/V
Zu+4FHxSd37EwfUfSzQw58SvmD8Wsx6Rb2JxU1461UuZaZPiXUf7M/WD28Ip+LFh
X4vR5toxX/5uDnseugOg77dHDAOFNhR97tdALr7jcXt2n4YDnXK2RcL6vPmtEE7k
sdONKWNSnrMfmrKtEkvJwQT6YDZuK/Z6jaVMrtGjVQRUDkabzcUx/AYtz7gddkLw
fjFlGxgqP/S60sOIAtTU1d4ExptX3XNi8to+RWny0xcJ6+vNa544bJmuUmQHLQwo
EYsZbJJ5E9vJARP2ELMoHdz0XWmWopwzeCQhKrFS6ok3DHxVP60LCFFdL0tHqFWw
M9z88G6uV4XFNuphe6gJWrtjbIDJitSJ6YUUREd10EcbLiEcgJaBWTpiHbps9BMe
8b3qg9ZWNlLwxzJT+N3mJeW/LF1v97OuMoowrbSyA/MZMxtZpMbRjuuoOZyaLV/g
pRrtKSWPXL/MRLS694B5OYKUg7Tnb4bwFBM3UWvqUvTChuTWwQXbV0AECKvdGaud
uZi2bRwM/VMEDmoTNKbGkMWcS0f6vOcdc7yB81vrAiyFR7ebPi74AJtUa3UlRWQa
J6Xk6GnIu4Vu4gIK1DGa6CE/qRpweVb/IIaz5oyL97MaGfyEcDIXYNuj7tMZGDwQ
kex5QQUWc81YjAvvyGKt9NZIjz0/e10sEo6h+uEKIc46gPbM1Y3Ykj+lj6ZvPWTC
83oR+Dva/rP17+uWrVxixYCR3T9aV+ZK4rGNcJyXuApmnAw8bTlKVLPz3sMN8ifo
/nMKM66WYThaSg1w6qUTYtm9CSet4djg0lSQKlBuVpjtjdtJFScMRI0MkhXp+Ri2
XIOx68gUae3STC5VdOtmEHxAUpDZ2JyKb91jVv+k3NhxHOjSAJpKP/psNDFiFsEi
dAHxU/VVQDUZndnJSASZQ0uzWsf5KANqkkMqaaogBoPpJL3g2ZRTtROiWJEdQwL6
LYEhYMZqAZCP+U20ErNRzA0XaP3b8xi3768zO9l6oGzKdGd54RgGnfSmsN0/nPzf
mPgScNXlGCCt1aU6kkK66qAV9XAlUhIeJYpnZ5TBBbigeeshw75HC92EVv8VbSDB
7DhK1pwJr6+tGoG9ShuvlNX6QAPXscFzZ7erOrQ/e10ROSrs6jMKA844teQLazbg
7b6oUIIizvdmOQuQgnOH717t1DI09hMtm3Qq+7mem2WAfIdmnKJubsVLxaiCerIW
y3Yj9mZbBI7/ypW0vLnHRIZT4W11gkHw+BmfT+ifOZNfcH6VeZf/MXXY/N++hwWs
OuxWic6N+/xtN0vqdbfY9928xF0YEKMYnXEvLYQTEt50Bd+ai5isConJ1juUQ6kU
t4KfcHRASAr0PEJh5OGOLf8ZSTvuV2UokYmkSeVnnTInD01L/jIVGusjqjGJ8cQD
wHux5RLBTIbsqq3QGe9Q/ecpOOlrCmgiyV7MADxSLpNslZJymfIZEplzOiK/MHvV
JnNrqPUidUlywWwav0GiNmOJSWG+yfL3co1iUSEkTzKf9t5Dhxe2Am553XFgrFNp
23C7Jn8PnobdlEue3d2cy1xZVwJilsPXVZHLXGIo4MfZ7nFHxToWpiCJy308P5NR
Jy16IxY2Q9sMtIeckU3+/d2Ts1dKiQcGD2KiA3G+VVpLB6Mc/sGGHE2Tx5uSpwzP
HwXrUjxc2l7hBHEImBIZpNeEAmI9NjTcPJ0yZ7Fs2GywE3yfWxgVgn9f53I1fyWD
/2uV6JvvpahkFJ/NOW3W4XUqn2gUHGKT7AY06RkNqrHZA5yo38+Wm9AjGytdrsCx
Nz1UgCcsomtwA9fDGneYBEtWMmsiAZ4yRwXsMs17sdmnBKSjFndhw4HH/Zru8F+8
muAit0eIatMVzWPaXHcbCbukPHpyzo8z8HSBdnRnPQSmI5L3SryeYRtKC2PpOBAF
Dfze/LS7JMN43wyOKGBXGxiglOx71v5JLcJFVbehGuVRPKuSbJMSYuAayjuyz4yT
Uu5wZaE1zZRYBRNO+Wa8MJ8lzVh1hU2akBHCdmYghJZEFbdiJskvAPmNFQ4AYcQp
Xs9IZDbZk/ABI0ONZoYF6Yz4jPUDlfQnwOEFNzLgo8gcN6dVChXvN2oST3QiEdUz
4cW/GssSMyWdQN6/9dCUC4uA0P+1J3S9FSt//wmPWlObrB5keGkpk0T/IFd7QKfh
6iHFLw7JVPjro7EObStlDx9PtTP3ROU61ttXfIxwWTi67uFf89O7hK/4vXCd/RCv
BJGH5hWN2xubEOHsnc4AlQvxISgGlE8vhec9X27ETu9Ij62jRimrDgEyJjMGwdXZ
EX/SpNU/8aNcj7vSjoDy+8YZFKv8uTCV+jlVv5MUECW8i00GlexVpLS0EkA2Ydeo
RYOR9Mbo6gmgWZamfB7K/9oL64d72MkfXZ2iQU0hzZ9xRLlqOZfpKL1R1wPjF9ms
s6fq6DEdKu5FQb91PTzrqEdt7zgd+MfmlpFvz4o6A7JT9i1YFRehEY7Nr4TTp0cE
XIdottCET5iyJl2lkX+nDm1G/INqa38h/K/Rgj/So5ulRGlMPDaxQOLFzQDLJSI0
ZVBc41FBJ9U8Z4XFkouzLYjoWGXH1tmnkYqCUaLvsXSLQYuDTLHExaXgM53k/+3d
tfGW0MK34r15Mzod5uYaz5xHVBwzGqDQ9oVWWwQ/0nEXNTaf51PJw+og4qV7Vdcp
wAh3Imvv9tdWeRvpgOijKS1Th1hp0b/Jjl+wXtX8NOfJXy0CJoPl+b85ky2oOD8v
81FOPQ3WWNqYtt+vMxQ3cdOh8xhW+z6zx9wkq/HfjFNTHyko52RJF8kg6yng6f1K
8xB2sGfxTkus3LJUQ1SUzTN9/o/CP+raQuccjJGVV+IlU5GYCYMH1L+tuFm5ZpLN
ZIMEcg406ishIUw+dR+1X+z4not2PO/4cjmSeBeQ+zJ3AepZ6PoUU4tNPOZo4kX+
axVu2a6c5cabImu5i4hKXg4H4YpSQ6MJe3TqnlIDPAsth5ctRY2MLncV/Hw4vs0X
mm7DKwdSvPUATRyoVJbVpNSXcMnNLDnPahO1qR4AsIiJXk3nqDSWhTHsD2r6zaEE
TM8IrwWkXeLPNsG07Znq4jZWqbt2gd3FkwHP20fFwstVQCW7PuC4S3f84owr5Z9F
4j5yCp1kPdfnljaC2PdLwwrfX/qUxTTBinBfuO7UISBDszrwbue7cd0zSgSfoOSi
vtcJxjNHSzINK8JDarUfBl81kb+Ka2HDfHJMjqmX0YncavklJwDj8v5DMrWDLM39
ZrCzqyXVKgmiMAOj5XzjyYRueWtJQOBD0eo1zbbCcXg+Reneq8kvFcqtULL+clYS
MC0FlfLaZHLGvtF6UKaC2DNVJ1vZevs/Q4x5bx+TKUuI3wSSE0+VUGGEkIutobCW
cEmCK5B+oG6TFpufULMwGM035SlZpMy2sDi/p7c6f3CcXQFoV55MT/SMuvpQB+Aj
FpztZF2cJmYzOrZBMQl0qjktrXTsGJFhlFmqho1mDWaTqFgRpaN9PziK5eRIWufA
icymN9XAC1fRBDU0A8388LSDtZf2zdy3rXOYPyMb3Z1UuM+fFtr2fF4JA5VU0U3c
TDU8scw0/Tv3dz6P2bbu+Uw6pX/e1BEkrPGT9XlMlwNaTodM/GAe90dTGvyz5PDH
mj2U1jiadbihh2yxB1CW6HeojU1P2ZgNeqtVPV6G0EFqm1dKPamuZOlOR3hyCdnl
nZ/VbcnMsFYehV96zL5JkdX9ck5RJc3cTDvd45i7Pm3HL4WXLh440tOvQczP9bYq
FoyMSaGzCVqojV/Fa/4zMIs8b/JRohVL6ZBgoQcgQ0ks3g9rNjfssQqm9wK8NriN
FDERkdtGT4Ykk1gwnZujOj9ovvvdfGVR65OAwfgG5CTZ07lVsZjtT+/nz7lrbNyt
N9niLQlBcZnGA5zLxJhioHeoM0cHQnKuvN3mks79ZddychuLb6ZDe+hqxZV5q2KQ
rollaBBXeM2ZijHqsOU2gzjdpgo5/9uijA9wf9v8Qm6Qk/LvDmlvRPW6RnFzslYS
7dgujnTEHeSLngDfprWKZzM8+LXtOX2NSSorIi2XOxVWLG5WncabdK4ti5FNojBT
QOwQqdQo0gK9is69jBGX6jqXPKoFcvBY8A2oP2hfYEU+nHU3XmOfF422UWZVGR6l
PGdYxxRYhLCvr1t2d5PvxpcXw4pqyM0OZG0rA1wBDLapFvGn0Mw9PT1bdtSB3k+d
bm7FOwg6h/r8ZC2ZdNMFdmidCHnpcklbxaPom+wW1361KbSte8T1m+aMh8f7KJeT
4NKa6Q0YNp2UoUbHyiqg0Oo2GnBY1q11abfpq+cjQfVZ8rQfK2yAZd82kJyUwCjC
NEjNZq2uaPtkQbNMNPzHIU6z15uF3t7MhEaOEBdGDkE8sXUf65f5ncFSi/s0xZgH
gOlvWj1JwjjGGczZPN0o/w/+R4uXW8nTR6iutNVeNaS02a+n/aAi0efRFlsiILGJ
W0ek56Bx+cVBCTrcKSH9s/Dq0GlWdz33PtDsZz3m0mWl71BgJGBENelm//mZknJN
KoQ39bFnNk9ZXBHFQ6Mqqa8Rn9tD0oDRd+nwqFLIcZ5YEtkW1WIMf/9G69hSs/Y7
KbkOOFRHHYR40ZRIZ9ZoUtATsZsUb0ekkjvIGpeI+T2hpcx11WC4eRFHOBrctxdj
kHUYmM6878sP/uswnjrZAmgyY6hFz3GjiBGn9kozCiqozKGnplYfzPvXasGXTC8S
4kp1fmkKFIao1vj8X5Q9A3B57JpvsUmqhVkYwIzAGo1CNgdpmw9qeNSNBEx0LfbX
GU1Dym1KmTFtDmILZMkDshZgEx4giOKSP2FgrQc8bZDmsVqM4S/cO5gkXArWvEJn
5x/tKfyjYGcpCw4daIVa0h7HCGKBNcrXg5O+a0AkmPZME/crfuxf325Vra27nUZ4
i2hp7MStejAoyACob/B3HxBIjfXdfYeOt+3RnXwkaVTlIdP6s/RWC+1rQ/5BtE74
vASHUhc0tUeyhypu2yzy5Q85Mg5LIDBMbuvsGvI9ZxhFLpGIU8Lj1g8yUGxFrwnt
i4qHRew6uff1VH2yHW1JtB4AiDqLqpb8fPtyxT/T56XIL+JdzQp1zUuvt0CtCLXR
IWr/U1bRqiAy94GQGVNP/w8EUnLAG3lTje8ZN1G1l00nnWJstCQ5fr3lVtKUyZui
YbeVJn1OVNSm5txKOivkS+hzZDzv8Ojhd6YKWsbxyD0Xe0GcumD6ec2HidBGEts9
SbSczsNnfNdEglOMZ2l1vQPvsMb8zz5M6s1Co7ULDOhLWd3ZoiVlYPq0B9sjbWWj
mFyBQzAgzvo67ahuvucKGQHwu06YVZI0oGGmGfQ/hReBthPVpYhFOTwjp1b+Exkj
S2KZ1l+l0IXTgWcvxTSvnH2Z6wjD9HX1rjZffPfLsN1kPQhogl16Ynsdxxj41zup
4tF+cuSfSJB4ubvC6LGDm6+Pkk+K70SOPppP98fuGOyGKasbKPOCpbno4Opt+sCe
BVrnXQWLcD0Em7q+wKLUzX8qhO/gaX5Q+zoP4MwkSgvp05js1H5Sfm+iCLBYk7Wx
aGPbnOSaxeka8AS4KpCTws1B9ziXaIM00SiumsvxIfvfOAbjO6GcGfE92FXdsffN
Kk+TF7iPktQ18MJcd3OIRYMmTWwTueuYc+/6lZ26NBuqJDSDgLWwjFNQKSBU9uZy
/rLEmh+SBnXqf3z1SdlE+k/dgNUaPHkb4B70vR/8HHBotx/+MPyxmYJSI/WJboRB
pFif+uxAUNUzMM1eT9vvhQu6W37CEf7CY3V148pWJ4qIXIoyDuHHraPJeIUr9LBY
MgaKXmN8OGDAbPEChNzr80FfZxTTq5fq+QAqHNEBcxaNmakOHDWPinW6r6JetEYy
IBD2niFRgROaicg7WFk8clA0rGbaHeEF8iIIiGFGAJgbgl6kHc2Ts4DLNlS+mZp2
0ZKbnzCiKyrlcBecWPzXpy0PvMeX66eTE5MsH2MamKNnZPS9GzxbBDJhPt5qZiPi
+xRzVBrrihShiFKApmgPk34Uaw32AOLOMYjnd9mJsUQr5MLLTRsaaxwJ2r9Rwf5L
RXX7FNZyauslyQtWAsXmelNNB5W7NHcIkyVx5+Oix9ut19sotWr4ieecmitY8Daa
M61cNAKPJMVDFmyHAqDb3uA/D2lN28e3zGwr86aV3CD5aCLp6qzc0vUI14u5NWuZ
t/cnH2gQxrCBmwWTREXA1URDPV5nhS3Qp9CwlU7mIlKhxt9FuvBqEnhF4s+Ox2mi
yyUeJf34Yd3KN1DLwtnEu+lQCZtuMSs3rB8ZYKMF1v7F61lekyIB9N6rZUEyLEKe
F5slWd48A6ppQZl8ILoy56ViAAZT6mpkz9SjOny18N8BsMz4t/z7ka1LLiKeAlKX
7I4EKuxlHPJ4BNVLd/A8fIKTn136AqXB85Q9Pe6csIPNICc2MMwZgV+ChUg2E7Xj
e2qCpTC9Ep5jesNAPjCNXC/ozt+LuO/H/Uof2Vlvz3/hIVHZOgDb/kmFoEy+Ujzg
a+tUh+jFPMODddb+83AkwCBOh+A/1PDAnKbuGF3zeNVm3obgOheySiDOONV7wVao
ocr/hXvLy3T0AGFsb2TPV4nTHJWzYOaE7ywCMbDcWSSm957h2qoBd0turUoxuIKY
Tm0VjA+ebDDbekr5NaFa2q06l+fvV/yOVNfOTaF7oNddmnTSYplREDI9iMfIlHnQ
4DzZxohF0CJVo/71E8+yfAptNkimiERVTrlLJIngi9N6JG+q2lJVN26idwQpxZU+
NrMNOgTWEVtjn4OUdVb3adZNNALUPfLSsa836bvY9DgIYogLg0mo2cUGztcScbX6
i7rtDi0+HrM/hhPiq4bVQ6dDu4BnqsihvZoNkUdXSdZyWWBLX4myS3HNRPY+jSD1
UeehogmPRsjmK4bcoNXOQ1UwTt/gNOl8xs6JBXajkD6YUM8zQpm/gEgpQ5CXz1xQ
C5o1OaF4NGYMXjWdkNtRIZt3q+zwqnim5UjsFA+4AdvLyU3H3r3lIWtRY2t2uI7H
I1vxQ81JDkx5wXEE9ZEbRzzL8UAIP+SCnudWk2KO5/PA3KkSvuVgM+6E+2gYU4LU
S0iKfEK2SYKF/Li4AGb4ZxByjjFjb+bXtVH8F3DNx4VjznarOWJ1wxY+SqFn/aql
uhh3QA6Hw801J88Q2EEeAYJNySqf6lR6U90GAmn+PiIT2mRNkxHBYYbASCObUngQ
wwOLUzSz7uQuNYi5fRUu4xuT/noc+mipk6hRL1X9bUO26ksxfPnq4eoF3yINhyUe
XHJi59PRCqijti17P96G8M0FEffjc/ox54LfSUSbswqkZiS3dYt2J7TAzKYCeiRE
OmNEXkaalWuHOJzgaBi0nEcG5dMjKIMz26oCA+W/BfjtWX3dOiIR3jSDGq0rggim
DAsSlTprsauGJao2aHVyRmC9F2NRrlkZgx+13P4a1bJ1LXWwATQoOl2BlhZqwPjv
opwW5JkxZmnwy9RX1B2iFiZvgFfMsDjakVrJYXgal6iDD+qHZ9U+wu3twcyQtyZZ
KGndOyulzouPF0tlnafXIepZWCW7epG+f3VysgTUlPCbRCzR2kEetNKvxxOeJA9T
JN4biYbR59eZEGnRELCWMxKw2Exog5KsBGmUW+g0AHjEc+Qp2M0OqcRZIZgoeUtD
W7IvnWfUYzTkIGKmk6mxQ1nQ9y8+wmoGHrvxjzdixTqUa0LTOtqkdpEB+X8x2lhK
eHeIA+ixKdGSTzu78l3X7jByycFeLLxExqLwKMcsOvrO8FbzTa8UxXwoYUMJhaoI
rtQaiEyb7lJ5vSAJy2TaWBzFTefrDqIzf3AGSMUfUhFYzuLbHVJGu0YJp7+EkzMi
vKh01LivYN6Q8+aoM0wdpAWVh2kds1/HTVfBz8kVBioTSDp3/4AZJdBHTO0c26qb
6F+0QooO2svQTIhlwsUYIGqo3ew5aYCmWcBeZLv8e14sj09h1QWpK9UuS2FQ83bo
rdvDNFYvAVrHuPqf9AeISeONj6dmAJbxMxjd/0WyAcq/R/U2FRYB/BeNSdn35ICh
Pp6XgKdIICUcU0+ljO/hShzc+6ooOPJQQacDRmAcyN0x5oM9OihO/rNvyFFMz1We
ImJMsGhbN1cNPOESE8ema81rEGqPgcABVeQNLi6bxBDW92HCSNN2QDcfd7yBu4I7
0gcMPYM0hkuWcB+GH4DS545amQvgtMdow1Zo84dweVZnal696klfNnSKHr/2bqQM
tMLqu0yC8JgFxD8hYUKoqv8zaqZ1LlaHgelwNQeJIlTi4MkyrEGyeyI2GWcmlqGI
ZRzi4w4xQSFMCw+Kqioj0x4G1VtRId40lwzA4uk1UYcptffPGvFg86YNp/gYh+WO
OcE4UbmXFIxxSyXszPcDg22Rl6mGrvdCkhtSwEtae+RhYGxz7KRYSJqKlHGzJu0v
kqqynnXv8mPCcCS7DLVtbFhjAVVXQL9/uGOEdeclrnXMWj0MaP2mCsEF/GusXWsO
WUElmy5tQvhqvE56g0ltkuvFXPuR/1JC6iNInMKA6+Cgnes06c7URB1TKXa25t5I
TpV1Crj/o/90xRsjDbaZE0ctDHlyBvCWPDuvz+A1cNPTEu4B0JO6kG71w5QuNAhv
eZXZQEJCK37OnP/OHYro4Tx1PdIa5zciL11oJ/g7Pr1EczV853di7Znig2Omb++4
/xNGLg/rD/U7JGl8dXOl7hFVcy2w4T+DoQI2IfTAl/EK6EhSPPO2Sa3l5jfZfyVG
kkxG27GcarQN9XbPVagBCIB8MBZruGJxaQcpvQwbkQpVqBAvxFm5i9TBOGvPlcFD
lPqqLfLV9o8QttzN5wAfMMvL65FSZLRmDi4Dd1bE0NBUe16M0BnZ7cEHipACzpD7
EsEghBoYf7lWafnGFtRBAYBHoum5Skr7dE0NeiCpuL2ZOvsPSyNjfqJDxjv5+iiQ
u7b10UdPlmk0UD0D5tfmgz5EDbC7lcmhm7rc7yMp6PjGM85Vf6AdqBfAZY0NMdYg
0riZ9dg71UpfTs1BfpI95KqBTHgemp/BwraE3s1ybJZWCoMfuRadBQ72tOjEkeYs
2sam0+SgZpid8PGO6icpKa2Q6VCEqiyoxX8TT6g88RhtyEqr2J1FZIk5wwQO4SZm
jshensm6EldCjjauIYC79nLpOORS8HtJQ47F+cTBt4IbvQDaCUNALxAfXzI5xWT8
Lg6c5H68jA3z+EcZb4L1ZCgVDgT5/gGwW3FX2fnAm/X529eZFQdEPMYO7RdtnUgp
4gQuftnF4x1Q7m0IkXzpKzW0lIyrkDaDFu/C0IrpVCrS3udUa/KC1stJOoJ3QpqU
fJjao64dmnBa8bHZlQwUEN4jkiEJPdS/pAbpZzilgMvwZfzv4rnVxttAABnRub1Y
ou15BHe4ebFlSF0rty8QELAjydhGjravkuHtBw6mN1GRWXqrMDkNS/1WrOUbvcTK
owkhTm1v0P065Z00XIvbPXkKIA6K6uSi23lhKJwEET4lyWgryNwGnZbdihdrepLS
055XocT3Cs2nN97tYKi1PTZqRwWzrreDARema96DVQJ5kjlnAiuO3iBQQCPt9nZq
1lv366Ya6a3XMTiRKtlIvKtBSstEU7XPGh06yOBappjwzyDDNudiv351dHTmc++I
0Zm8np8mZTG8Lw6FVxTJHjtFEAl3/pbyqsUENnvAVisQ8wwbtMKV+XCi/y5GcFZJ
IHGbT7NVT0+KaXNdua/7w9JsctE6wCyjc5XyFjfHidI8s6IBD3775589di9LZ0Ec
eipBnPi5ASC1jwRVG4hO4l/DeHSDLy/nKqmKPqKu9O0SlBarIH8E9H829HUWNDEc
A8XriGquDO337Tgf+9T7vaXW4biSf5MQsU2jZ8Ntwae2w09iBkuvc7j5IqA9nU3Y
0qP82E/9srY7btK8O6ni1wF/9w6YhhJiVXOVQWQFCajNSqbp2FWOPwhSUfktubmK
1TlbpZUAMj62RGJYvC/AHQxkhfnx2OZ+8XhWp3+B1Cu4e6y9Kr6cIEcstKXbuEE5
coTJorJjFo5ix99eSuQmMDHrxkW40fF5hLdG6JP+DN0tTnWJB+kpdUpxUN0u0UGO
/O2YPTZextRkn9P/fjrNqPIJmwXxUDF2tVayduW1Anwsfc90KubWmz7YyntNmhR5
Hf5KX540LhLWCV0A5dPU8ymnTxD+KuHYCGGcnktLOLGPcRxj9+R0dHyaV7jFtTna
QwRsZoRbeCefUIZ2tmbMrjy+k5JZnjdGEKDRFRwQrDUCSeI6/Je5iXsO2U3eq4id
HbbcbFc82JMqtVVsS3hneXStlnVtM+giu1Vk6AI9fGEQOWnMx46T61/k9B2P61mA
GwyzZXR2cT4PMjEjmMquN3Mh5QguPC44lIq6SWdRHsSbVc30BdzOqGrQqFhQt07E
Wj/oOmmBBXLuK0g/xyeqpZmWod/yUFr55EwjLNlIQiqaFYGKb6Zi9AHqAck5vtv7
NDai13v8qpa+S+4kzZMEUdntDIzidsysDSRbvHKU3XLq/JsP1/ThnkUlVlnlw0KU
L8gJy64OoOB91CTbjywwcJ+XaCQgsKh6RDvn2KT8zRLtCuASlvesy0ERT9ZW0HwR
LykdKX8fmgx689UhBxcNCjzQ1L8Xz73UyuZKBjo6aw0dBEQZk9DHsbz0ho7CSrhf
OnLN0fiozVITRj6vHhCIc0JIK6t1UrwlgMBMVZRYeW9Cyr8UDFhl7+Ya2duVy5CJ
jWBT0OBVxE2wPQ9j2DuOUZZlDTOOg0BMrNK6gzuSiRqHtLuqIgvV/CE4f/RhnKKI
YZ5iBXz0Z+wr1gs6KGVr+6wgtlbS2Eozg0SZtqHfVnER2sSgeye7wniCyMVDW/RT
Ku8TjMxs1dF3WYot9lNehQqpvWzxTxv7WtfwYzUGRTdzh2SXGds23VZhzn6TMhCb
8V8QQStbUngfd9Pt7+5SFG3UEdmnHEvUSFWUJQ5B2M2WNo/prafhmvybbU93WfIh
GL2S02tvwRjQKZt9N0UJOi+dIbyPbb+1C5zqLYjZr9R3hTFdR5YcvJrxb0g/boR1
nSzhNNy+bN3838XyHbfZw3mkZ2pRteG8ngPjA+2wRRXbr+/WagX/9Xvy7a8PyUBG
iQpO7GKTgvdf4Tx+Jx+RN3YgqKbj9hhVwfA4Tqkn46xePgPagAgi9/pVA/kn0bEF
Oyih5DU4Rdh+/1Tit9uMJEc97R+3ggMms3JZNNQryZdOKoBU89dNmxWhTBSmO4/2
SYszMyGDmVMh31ZqmptxtH5PViwn1M9pqNH7MQzvkqz5u2mlJL6RrPIVfAYjQ+s+
nK3GxEv6duwT7Qa8PAIIUV6N0Y53KI0DDR3AWjVo6tGiJU+b7De4n04p+Rg+aICC
OK1J7T+3qnpn1fARj+xtIx7Soj2ORtYBDQg22KOg2d3f3NCOPPVpCk1gH8RuD9rE
wK5lSstUD5SgbPODjjGzte2GXS5JBCMUL4DvYOaDsKv3QFAvAaJ6V4TDPR6rbCbq
F1j58Zdi+Cs5B0PhDnCa/MbAzzBWLqJwV/FsvTQnfZaFD86dyVbdpSynMPvYbG/q
U6q1FwI2VN9ufbjS4VHCT6rsXTRNsIJzbbJ9V/rry3m8/8HlyD27J3orlZvZP9ub
GeNG9nmvhBDIqptBADuRrCC4c0mJXvoIHke6XyzbfwuL0eCh8xLnVn6eJyd0Dp1A
vSm7mjxz+mDmmONnsJ7ckoeWPQ+ggsDKgNXEKkjZF6vHHpdOS8AxS+YnA5Z2X8Xz
C26qHal0DvkHami5y6/swr/Rrb2LWl+pGYv7J9pTk4UHbyGJQYH2y/JIif0Q8a7u
tjLaKoBs0dG5uWR6BOS8U2qTQTNntqUc8UNtVMlqFQ9SwmngNt0mslnzZnMIwneV
ckFdeUyiiKuHUH4X+ZOA2xM+k07WGX64mtpe93+7NGO+1SE6i7AXWaxT3zXCqMLY
ZLr825hHuwBxHf+CKYeBWSmmYeeZff6KVSG3EGM5voph+JR8NpeKQaws9XulfbmV
RX/9KFPS5NzR3MtHhmPg0ivMdqgmi6tMzePguyzQvLbg6RYZCE8O7XGDhBVjPaww
aI1Qs7na+Kf7ULVGjwydt+WZq9vwsCpHNq3iLdk363faBX+y3lvOBmrUlk9M5HaN
wJ4x9BZmeBFaUUZFOKqpwmUokMBlWEhr06GfPi+jAgGY21K3mbK7MRajlZLfNCM4
4/2NL6il7qgypCx/50mNshr/GaMnh39Xu6T5OliFP5W0gpzRWZFiQ1EvMtJBfTzi
8PajvR57x1xDJB83QdBxd9UY7nzrrMpG5KX51esHTTKB1fuI1Ni/NmpuDAcPjgxQ
aQ3A1Sq40oJdrPx4PdB1xF/6CqWq0rUAh5g6ClTDfmX0xlqqWXoeckBNGlP+1GtQ
191I8+d+jzk7wx+pFkLLuiF/nAs5tedP5AIeBwZrjWR5DxWWLCkqCW6P0KOWlz+I
fHwy4IkQvEFiSUkZR6B3vSNgQ6y37T+XWZ/Q6ey0LQWp4m6tG2DQCrnissOjHHa3
Hi4R5OHV1xL0HkVGDd8q5VOL2ylyg/i/ZpouzaE4yt4V9D9feDWvFHTecIZNBt18
A2k7UBf1zKz6bzblAsibBva+4kQRJ4q/4unVoGvv5w5DI4w0UEx1ySTLu9AK0CL/
FlOVGZ1vcGFdqLN72kbYiqYuu1osGM5E3GG55Str1Fh3LlU4rmmJ1x300YiNsQHv
yG2RQbAGMkQEP+jqA3cIKgSShVBemEXgNQin32/tee2RCPKb8JxO4crf4B+j7tgs
aCyZaVROp0t+2ak9qYNf7lv2KqGwHYe3T/fXZO0YulmNry41ytzeKOxDlDffqTCz
lPRTEMIA3dV1lApPYljYa2O4MTkw5BWmTG0HXRzvqCrU5OUYKvlpxjR71W/LdJ1C
vIvq+oCm7nJimQ31bnS9++JkneASymmxu7NyS5hgWcSCtOIG/BhGFFdyRLvySebW
9hV/eLKWwTyZEivRHLeekctALNITNKyAbMEp8I5pccm+B/7rL6h3PrKyXqW1DiOB
eAt403oeo7KZ2oQJUXjQfGgfEKyym3ZWzURIRN0lHZSJHWYS2Hm+sS9dLVSWZ1GE
Iwlzh2LamM76ulCWd2Jhdb3ftIcgonAiGU+bntvSpfQFYmkasm8OPLtqQui1CrZS
MAdveSUfKd+DL7vaGZX2jP/h0zBCkP6gulkVY3sU2M85hYswI9bx8XMMnGdwiibg
nYzr9ExiUOwCdaptqTKwyV+XA4ySX6mMDoiQY+rFmhQm4F/z/6CveKJflAWGVSPS
hlYbf6bNnqbpwYl3CFP3j5hlqtpH9EOd2eCobWtgvotv44/zXGJVpFt8tBs+fpGD
Qto9kwpLr0rciUTD02Aey7655Zk4WQ8M6qj8rjlIpw/czecfR6IeJGnDgyVQJBWl
kw0IRnr74DfBdo/3LPgRkQP+kkIAANpKqZ7ePcppe1t0PUTD0iYjvWUEJusiF3lz
u3oWYumstHnqmcH6fpfBqMjiOrXWVYuKCFFwliXH/BPPdNieFGiGmkadd+cjSFkL
ByyWbLIitqy9cnj11IKZ8AXT6J/bBnvHUy76G2Bl6UkQCOS5Q11zw/vgC/DHfhRC
bTgcLZYh/VcfXFRmb9qNPOO8A4NI3EO0bqp/cF9aK0wn+7XunbmMS4wUfjxVgKD5
lCjZQBmSUmxw/zu/WX9p8A98ikoJh6jhT7BnBQ+jfr5BiTrSaip2LpFHkSLzOx46
dzeQ7FQ8FGGDvWvLBF2fCbkEXqjWk/j92oqxPJ9i8mRZc8/mz2Lk2esUp9I2SHfQ
8cDCq7yoNYpHsvUhshfTVRaYvbRBRnJwmJpWFRd4iW59fDhIaXOWdsPnQIiw05L5
LOj9rf3LGcbAszijr9caH3wWs6HbJayt/GU26s6trta5psoQOjFx2swOQlt9GdzN
627FOof9BypD5a+ix5doOgvd5WaSKUXDCxLuNuUVAS2xoqhVIL25lQwqunGPpTC1
1TIfBTgSUnmWZGwcT05tfeT/Mpg0GfZW4gVKTYj84Hh/atWfZ16jXFQvqErU70bI
sEZ206NOuVkxdvyfXJ4irihwyp5Xcjgz6gff1TROAX7MQwab34ws1nqZKJDEg4q6
69l2KFNIre8NbvwE6mfgCQEKweiU6tvNCNU4U2kDntDGtJwD6pGE8flbvmIcQTyG
D/dRgp121EwZAypQOQsWTDxrYmsQ5Up/h7QWfBhb9yp8Stcae/wdO6UHmqWe3Ok9
5FJAUuKbhyyAsr9w+0TfaK25jqO8L7YkspqkQLGCNf4neJdwQdi+bo74vjJMWTqW
G0V+vLsOMgfn9cHpF8OYJl0s1dJyxg9ayLkQU6hK9qD9yvLg3O9x0KZVIG0gbNdz
hjt/Fqwf5zCoZ3HFZwTGVhuaueLJSCos0tdJVWHa7+COAaJ9Bp0wa1csrsj8+A7p
AAs9id5WOjmrGRyhNmJmBekvWTd5DvZQHV7xxVuuj+CXqKzfQ2kreCrWh0zsW0I6
wSI9hjRxdkxzWd4A1iCCpxx/sjYj5aSMv7LLnDYK/rr/35mGK9+4bABi/zQkqI6D
cRzhZrhZRLdTbeI7R9+3k+AMWEqvbpRMNc0bLBRSBW3HHsCDBjMchNpDPU0yNK0j
QfX03JncdBSH0UhKDE/H1fVCGNtpovw7I3qnW+U5XgceCZAlWeXQbs0XvkwgMNOa
2Mach5SD6kVuY6vtWxLYtP/SL03iIuH74Kq7ENOfM09hDlz/oRYK8j33g4cSh846
9zR0N0WcjY2+68/JUG3sX+Bzz5gvBoNPxXbDg3HCMy+rzDAhC/KcfXveIQ999rVL
DVmsh1SNxWIVngcvYI5/dzkNukjmNB41r56ctxCvB9yZGLsXuivuJO7RXFjYswMv
LDeDBmmjFPmxHfYbx7uWWQ==
`pragma protect end_protected
