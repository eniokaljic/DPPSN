// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eoTkNbn2RgNzJyTKYQJYDoV7ykjUk6tmrj+vDYl2ly01bt78OkXokm97tSFEU9AQ
p1l4OcxXIoPgbzP61yrfw7Vck8/ZWBGaF2HVFd9rFmgNfGJw3Z4kpXnnxd5FWM2f
KdFtHssey5iNk86S26xuF2pO+E5ocn662qX+looMqkw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29728)
mPxHD8g32yRWNyjTQFA+mAsqL3eQV77PXAmno5r2b7IYNHWz2nPxXKIkZSTzxMn+
3OiWCXFjVAGHUEAW7vxvrg9hlryvHYkrX8/Fy57A13riQ6PvkRhmDmicdM86mcd9
TasLJJPWIQsx5VgpA8lq75o//rB84loCKuwjB0xqR+aNze4acVNFDoNoOl3+pUAe
9PKriVhAWJ8X5Et134OElPjJgQJZGHiueGPIwplZPtjvMDRp+YWS7mvsvZtgcldj
eJiujFxxT/HR9rWUdmggi5T6nb7PzeWReoBOucUN+Che6EvUmY3rdFatEVP33Hui
x4hnPtoEmhGqXyH2O5XKuwXcxIf5uxnaSHLh6elKFiytqxu1pfOZKP030n/ZpUl7
THmtG1J01+Ya/muiTE1bCAH4/VGLDPkfZbUfsV8shJlOTizXl0+CnuYxVUrAjQQ5
1jHmQxaxJ3+F3s/QXq24uCh7RX9xvIUxWD2p82x9a37abO3oqUZMHRfisbFVWhjm
bRQ9RJM8QGe9zbgpcAuLnQu07+6uD2vpuEZn9gRd+2jFfYuCK/O4LnW0W4g+GC9O
BgBJ5nBMerSdcaiwk8+q/Off33MfJnvWhZn07XTYbAk9YBNHGLsNofBs2JL751kM
9omn/T05KjNQlm8Gqj5uD/dMNIVi1gkKw9Zp8cwpitqBfL1TNqykV6QX9gnwyezO
f0x01JSEds1x8oXnOH0YHa7G4wrCdcVYJPDQou3bqOxzlSnr0xdlEt0AmWLgCPyV
oDEfudGUEm/xi27OH4BjQiIjLXR2wcz+ko5TFc9yUCAGffL72d9czHlxkSEX37jz
CJurgYG0xPgN/GgFoZ4yx34QwYWnF7+SB0d9rarjlhaQfaX1ukEgZqYP8CfYbkH4
rGA9AQymVmv3RAOxNmvjeAw1PZ6UH9D2KatBxu6T429JqnNeXGkonvesgWLx19Oe
uuhgb9vkJGs+uVJkHFZPB4DYbtXv4fW93qlY1un9Su2MgIr7z21y0UU+gsIZidWi
WIe2n3WtY/hr5V4hceFJr8Ypf/WhVwztLVmEcthk1wMRsEzNwVkkF5wD8vXgz5wk
0E6zY3qevbV7UxyUAyjed7HM/D0uwU49hOuc4YJnT3ntZYWKmGW22DLcJ1J5J0Kq
3f5wWbSn74QYqduKGxksFVzf9ceu0HTOhAlARVkqOXPkFKcUw8Vw0bVHe6G6eW0Y
b6HlRojVQuPZ3psIxECaKSHMZFLCbeCjtDt0L6459WKsXgx7KpAjLnjqW1q9mD5O
8I79IVxDWgVN4LKvonSOnvgiZdI6OEWK19j663grzXxLydAmUAn4fiRUQKyk7YTH
T3wwQo3fyVOcyDTv3U2eAzRubrKCzGNxupjIe4lfpQ11IbHYnsg+2Sw6QcUeN8M9
vDXdAGvrD4SbvOjuqd6gtB9lfcyv6CT3YNElzPM91QqllFv79dLp08UcDp5w3ZUY
iuenGJ5+LZQoghVVMP4iC+mw8uv2NTqu7C51sEBGosUxfqb/Xi6ZclZBNlIHheCN
AipUs7Lae6KxmdPr7pp34ByfOovTynDhv6w8f1qZ0/8SBDawn7E+qO+oBl0CwHRj
V2Es0L8GZTdlidm8FfxK+5ta6t+WgFfEu7t43SyCKiyP4yI4v8NKYZzVC+FSZD8m
AZKa6YJ5g1PpiI3eb2774EY1nm5G6AuTN6RDSm8tpP0Rjz8Jw5h5/+kVHvCZmCeX
6BDekZYmVANT+x2NA9hHwq6H+rr9HEeWkU9IfnLS25DbpFYBGJl8aqAuHtcG16yB
Rkpe6LjWTNmxS5Q3f0BTTa3KS0BrNdM204mZSxNsIYCHzz4+uW2LqiGzwYz6qNxR
It0kIXdReuhNtRQsf0hUbzV6d9chfQ3QrEn8gQPFTHPksy15YRUnA6TeBm6UoRdI
53iaFK1IvlS9mO7AaNhlGppdzjcorihDNyKAis+U0Sl5nzoxCnT4GTndBBCI/kPl
DbLt+Im+NY5VrBsLAJURRDgi42PWi7MIv4OH+raaLRJFqp9Xwpdc1Bqymv2HcBiZ
eePMhPDxcbaOyYBLHsjOf/9wuW7ypawPZ4+uJkBug4qMFyrpyBe8rm6pHf1xPiOH
xMrjHRbG0W0a1TdxfnOFH9hTnDsLSiLDMhF3uPvwPPfInz6g/W6pltz4DmaX3DCZ
+irnoRH1pJAiflfV6UD2inufhNkcAefLNbVSdygXTqGY/yftH4oIA3WOmGpv5Z7B
7QzvQ9cTJ38JfRcr6YYEzsQkCWVojsfbvRMbIKd715cBypgbq7rm0QJ08caobR+O
ZbrRqiYwgiJKCEFX/4PYwkNMB2CVmqccFoaNJ1bvCXB2TUOBvqHLyQjtnLyVwsap
GVNDUJdVLXpCBqeRCwjpWsvC/xXSHpZ66SPZlClbamW3+WPMbuHtpP/P3yxMTXk5
54omoRqNEqnIe5JC1q09UVcLB6eHn4bbd9xYbyvkY8tMwoCnwScPecQLMuuzQAjm
n18JrXdnbp7AlGX6qQ3D1fF/ELZQ+HxYIlm7Ha+qqWGNS5O1P2kdqF+xniI/LqQY
V8HRRxOqpMnacMOo5cs+W190DvIkULANOsHURnw2v80K8/CUKvjlCNd7/cvAVJUl
l17xrMqOPE8kSkfshw/aaBjDBt0PZlKdZ7q1muIVEKWfYJCWa9AhbqFYaK8y4djt
2jOTVyeI9B6+P3iTogQbjbAOUOaIGMs3tiP3d3NRccb9H/szXPqtSqKkG+qw5peX
C30p56YgomuiyM42FEunpL0rTyBjcXmGLRSihKBb6fxzVkEDO6CI+ZDe7DmWFerc
dU2n4R3lIUDrsbXCZIloC6bAhQVtDMxPgLAw+VUIjPkBrU4pr9T7TwbXoxL/TWR3
IK556G5RCDA1d9l9DNoXZ3Ot/Y+0hO/o/pMR0Z6xqudnSEdxKCjnIZTDNy2qq4KA
IIsUh/tZ6io15W+42i/8WBRt5MKNnEUtuzegK7GUaUlcLnzbRdXjgU+mzzIVWO+o
OYD0sIZtMkKH6VmHSQZBDo3MQn1RmkJIBq8p28OBAD3y2vb/qsFV+Tyn9JKIvUBk
AiEj43WelFSTxsH1yHPzFfH2PkU41gGWp/YSaDfloCyWWZtjr6jTUKzvHvX9Cycx
+nsghsDhJwvFZ9KQnvW1QIhWgbOUhNwxz1Kw6HJSz3ntbmG5P3YTWi/ivUS+ZpnG
KOeBlOfgOVKAn0cDXAiMJVmPQMoGXk6oHx/6CQNGaCLJAbH/CKRHarx0byIerJw9
XEfWfqPOpr0RuLkJ63xh8KXqPCHlXb1G7u0IEUJhm1QPDlQn0XYRbfeDNEAvFt9i
Zw3veelX6LPfI/YhuT1oMfTzdnMR7VFUVh6Jed68ehvO803wqhA4/lUfg+FIWAcp
tzB6Qfs0AkJSE46tcuC6erZBI27QpnzHCm/p8O2ATRoE5Irucnr61GmFQ5L8SFhQ
WSmZCIFEdG6DlFN4HBrpVGYly1RbKA6uKsueyP3TxzK/ElU+rKwzcZYyfjaGM455
gPVsd4IvChUw6DDYjze10ELI0AM4FtPZkkr5VklJNDeRGEvoseF5XTc+aBnlS5+W
z82joeNyHJ9YPrd88d8J4nrlF4J61RNMTT5NtYXXv9AwgsAZmFIPG+devSNKDJrf
fYdtlItVcKVxd6n/Q+027AgZ+OQhV8AXbycZ/gh9cXL6ZWGuUXIk52zgB9UowI1w
YfTFOBXt8ttnqT97cFuy06TNH+Mi3yUo0Nycr/XROBCGr0j9xw5k4casTypXM0CK
9bdV+YNplA1tzQKeARfK1CzTF63VJuYK2MW9LeIhdkQRemZ+rI1oZ/LLWks6TqyV
dP/RriwscW8GtjrLlZwHaWxu3QR6eLMAjGhJkdZc0Y1y+Qz3Uogi1nDlQxspJZRj
QTHCbobLAJj7oIAGITtKb9551uIlzMXRBw2ulSkQdbHDiqPeKNRyI/BPpilghRN4
IkrDewdjgzROqoEhqZmNVxHCOV1/buTgRfuMNXehZueC0zTch3ML1zlVXrn3yddF
BoHSXGvc5rpwTw4rLfOWAGCb8dbAtjcTY0/a2u4kvm5nE5qKtMMzWmxf6c+gnkND
DSqIrjWrgWmolyFnjMAc2l5uQvrdbXEjMDsr1uJi7EGA0/+B//rrpGIBWwSXrkB6
CuYEszaHND+VN7YaDYcXXplK5/Eug3xbz+hboUdJu82PxxJdm7eOODGH4OyhTCGZ
VzQUGbxyvhDGgIfxwzcTdN1kTNxkjMoZN+lkJqkiz8RIDo7GN5pAL17d2bnsDrMr
NdOMMsDmDiSW7RSPedm1uP/zlVI9swS29e220LQvnZrCpGTuUg6Z0de3if0SAOuv
hQQ+zwdUjur66wQPDJTfP2tlSeFiOIc4f+zIaMdM9xl9VLLxjNeHKLuQqof3Tv78
xfvtnQ5DAH0inms/Lra0Pbf96sPuOxmENtTX1scXU1YWle2zw8jnU976zo7Uo/Lo
kSs7Nuwx5pbOIhyCsWprVpDdpmRyjGhNW5OQtKTrNyyscDhqHbvYrpPKpQclZnN6
iZjuMnlxnBf/YfaMMquVekdMwJxIrZd0NVTcP70rhE7Ogk1e+gRMjQkxfTp3phGb
KZifN0+WoAQVGJEHu2v+IOGIydNEbj2uO5F9Nkz5Dj1wY9nj2AsawhFAxRRPluqV
+mpKpYgmhOGY3rjLe1JvvStUSdGQszXS/zRSuWeKxOZx0+kUCRj2cuELiGBwjq42
WG0SLVWjuhNTGoDGeBVyFg++F+U1FdNyqXbtBmNLuxZDO47fYR3iMxVMEtV/tzgF
kCofhRy+bBx5bpaHdY5UVBikR6NfUrPHCSHGHkj1lr6vbRpdghALFywPfxZbIiEW
rtbboPyznPZxnazCVMfg+flaWcaLfhAuIHDr/d5i+T8VTRgupccqYqH9uvVKlJI6
bwmbH4ihTPBBBjiu9prrtPdSo3MLIuTnj8gpsPreNvcTBNk3Bis6aNxncwdWvfMd
XB5z2ap3BfjOZ1W1u8SkTfCORYvdZ2r9LZgW+n8HQMGJBIdNaoGSnupLUT/r79mg
opbc63cApw6GVDtkgYko8S4Lq8x71hAH6Y6JgfztAh6xFCu5bt2zyN5yGAIELjMq
qwdRLEcdwaaGGf7oNvT2/UcP/q/WSMRZx1iudlxsa3kfX3tGaFO/PGZNZM6JgSRn
NdIPzsb2IBbURtTKmb5c1imHMhMD6Cc0ingCWpEYGG4ZQ4ifdjVzj0XOa02bY5Yr
k5p+32mgKcEWaEipdzD5gC/JeV+Rhi3E2o7KJR6eGJr7RaEqx2PvY9C1Osp8aG4J
4kqBV8dq7oFn5lV+RMIVlZFDE3hBston4bi5sJH8JOyqwHlP3Nnv6pBUqH10CJ61
9pXoXdNh997hrOA3hs2szKq/t/h904JUOEik4TYb9nRXQF1wsswU+/sJees77pU0
I42TDJOAM4dXs66T9r/d0TLwYyN4nSgZkNab2iAdh7/HK3ZqsNHWiAQ1Exvz3i+Z
ME5zs5a1y7IJ9dfPCE2/flRDWxL57qz8HIuJGkXx9tfFIvX4k55XsBN795bciziX
rANhp6unB4DHhVRLIJDeO8rDiGubLN1V/IGO6Gw679iw4RdCGDU7CLtFfY/Gn7t7
xU1WHScXbFziE4+m33eADXdvwtV+KZHIMU1QTf02IKiBmgaWLwNKUqTmWRoi9X+e
DiC/3EIVl32wj0gjXCwLJ26rF1+8lpc2LCXeNe+//GG8ETnCfP1sdaOwLEIeNHUj
IorB5hmVbUj+ax4gksnPyv9Hu4ZS4R9AtqxOzhSFoVIdci22F+ISG/sowGdn5Nym
rJGf1+jlA86mM/dHXwzXkuZQ2UgVAJn5r8FDQy2iilqWe2p3qdBcVJsrbozj0GRm
PpXN8JVgdrEDpl7imXr1OBd/Infn5V88eArET7sH0AHAjvBG2VD8YdrXr47n4/Jg
1ypyJciqgZ1pxAnl3pGEweUolJj8xGHbYLfAfPrWJUopvWRCDWCA8AsAtpNFWcDV
iDRyrtNU3ZBFBPET274ilk4ynbe97XSVjfCYZqEr7E4cH5Lygud+tevCh3hGEUEh
+F35QtOCGprMLnvHRL16qqH7JbjU0SzH3PTKGXeE2QsaAHEMAPfWIu3SeJBHTtx1
6OGj353f37Ho4ZUvZhjjQYv5PON46690ZqVZg9EMg+n7DRtRhJakKd7TiMPUPNXE
xgy6HZ0hgJ1anDtNXkdDoV8C+BDIifi7GPiSmhZ0KmeI2KUm+5TMkYb65Q7/CmoZ
EfNpWYT9P+8H2rOqsv/HIFtZAT4/1IcXIParj9M1A12TXUmxri8j8vzpGc9PnUEC
APs3io/rGuXkY4/1nqF0ieOKNNvidRp85aP+/NDY09wMiYr2EkSqEVqrUomTs/8Q
5YZmrGW8DpwxODh1Dh/XaVZwD1qRzkI1TFxwzkVG+oFxvhLnurbKZ04KSk13zu+L
3hm5SKWDu35Z2ftkwafDlgswYBm94ubtWAdH3HXdcm+6etHRO+4kpFLM1DEdUxj+
UYfD0GJOU4KKMEkOwbPj7QnAoG2Q//UfkYSXut56PJgkgIcBhNwP9DbrYpRGBKJH
JORK7fPNUSn8T7heqf5OQ/DM29685hrfiLaqT2VAfF0d/JzUek/iH57mX3bApuhu
69Jc9v1X1QKt/x7YQjmMU0h5ui9NngV7Hh5wCQXGQ1XjxeCQh79ujg74NdJZpz13
UCYnlcsLqGg7VhCArprO3i4EEsxhDJ6k4UrEJzwhW2k6UDOibgWxIl4pnyu1soNS
SEBlIrRMBZG8Uy44dNVgABYrcJN+iSm3T+Bjvx3GDCfy1Djf51mWpzThpOHsWg42
UqJ6AY6Cfr61VApukjIvQ4onp21do377rSCCtPjiMXtjtADWFz1/GSdae+eJiEgh
2Ne3DjtC7VOF1kyYlnJKDE5rRcgaXRYDFC/w8j00FVRgLB+IPn4JcAfpWGQKno1A
k3IyAzhFKHhZCyEj3Bmjrl2fdiV0uLwjDTh4EKe9D2l+LVdi0Wa9/G8bLP8Ui0me
qwZVIt+OailzlBHtLqZgAzemvrINKiyRiPbpFADLOgZBQnugV+iwqgqnQ4kQ5JhO
a5OEjVq0wzWPhBbkrIoXt61XEQgSta2wJWA7lQCdXJ7UMGykrXEfwG5Ejt6FCVJo
xHBeXg5cby26EIhpwIcCG/c2itizYGtSg+fVdxZQdFQDjcUpbGxuKJIyBkpjNIUd
GOvAEWHxhxUXY5fa+dCG7vyhDMLi+IWdQnErDHd7j2SSmmFjzIvS3nvhpihl4jyR
aB+ld0khUgEv6dQX3aKXlVm01my7btbECLJGrxN4nRXchRFt8VjvmXgHClbwucF5
ZnyE933FtfjBG9KmtfMQl9w5oomFRFzFe2AdrRLfB+t+Z9Ddk+tCUIHaRD3E2r3y
Be9xPh/GpcbaLSKYAznUctzo1Toygl24uHT3gUj8DvKhMaUH5vDzKynWsrPPY12a
75POExzEUFvhbyOo5gJkmuT4avj2iypq/bHqKAE5Vf7K4Bq4PuY6EJzOOOA1ilw+
aMv0IVCWOz5dZ34/+nyJ9XD5t+UDUG2jLoD38dYiFIzLM3ReuhaszKvFIRk/EoVm
jYUWr3AQw6o9iKebDKzOrNWmJ7ydEbjnnGkft4unLxodJFO3fc0BL/tc++5rw6L2
oGjJjAbn4MIf8LTgJbfea9eDcHLCoYfObLY7Ys9li+gsp67oVutR/rC3i9Jbfh6f
rQ/9BsFHyqDJpo7QjKlPUw6QewsZiATPdffhrQFEwBT4B+7+7K0z3bhIhhQye/3y
JQnEImDGSqnhpsV6QDTHvAQwk3e0tUfgG8uOO0XgT+VKPQ84b7xoTvQJIbAJjPtJ
hWFoy70NMA6TZyvKnJJOh9qlsZ6d/8WkCiEsCAGbg6tatil16ieYcQchpGAYMRA4
N8KHVLbngTYccFzPh0gWKwS5iyWNt4e+WDl7ML6ItkfefPtT7YRV0yKDQjpnPKkh
oK8S67JjUayxiVPjLyr078hyicPCrDXzT1Lsw1UoAAU5q0mahjncqYty3lo5QkVn
iboQtdtlXAJmDgfYOi2yB01mrBioz/ZmFQ1G9Gkt4o1AkzpdCQbInl32a7lLL62e
NwzupoZFs8ZihTUK7+x/Vv/JJJt19EleEfQCNV5TkJQRaALD3Fxb+GqzS4qZJcL2
O9ut4VL/XKKJ999+EOtq7K5W2A2d1N3inJU5oNBZ+nv4mW3+AN/dgSWLVTGMHFIn
PnSuNYKTNJSgiCBL/dUHFaCzsyX76+20Y1BvXgLfzYb/OCbHyNrWh7ZjrlOJ0nIP
TnoWGB8fz1Ob0tUds8w8i4f/kDkNbOlAq4kF6xcO2Kfj2T6IIRi5wbWVYuLgfeh+
03LTX9Y2COGGobg0ms3sFtFTwClb02re1bmUdpe8UhVwCWTmHAy9ej/WeLzF0uvb
VL0Aahu7KlyYf5w1Zx1VvbmQjxs0n2eHEhMhvWrZ7dRw7tBiScN83+eMUxdGUuc8
HflJVbkV8TIUT1PLrN1sdZWXfMNf8w18hti7W14KsUsE2n3gYnoIx4Hk9aibASnM
yM/vOuDvoiMovoclNj1NrftHgEGo613R9XhbPap5uUw+DjTCyO2Vd2uDE69NbLxR
Q2QbAm4bAg8JrZn4yA5IFcI8PPYsgMgh9Hn/TcSzHBZFL05WzXMcHKPpE3oD6wKC
vPk//GfMeb2YVH4oyufbJLThs0t4BMsm9q9VUxBd+4OBqBIRF92YCb7hm404PROT
Z9R9sDHfOcF3j3/sGGlNORqhNVtKoDFwM/BAsN3/cWbjrjCgKodEAcKjMEpSsO08
ujLxAE+upjrjfXB29PgN1GYHfURL4awLDEgptWmaVAGgU8pdMvwnkYWwJi1sK4x/
/nRzeMm4AYuHaAhqoeIqpm8esqh344Xk9GXg0XaZefK99dqPM54nrY9CcbWW3HPa
6G3SaA+JTYpmW0o7Dc+3fKXLSEeWiuDycdwrI7sSxjLD/JOcxz0yRB6Ts6l9zqoY
Sw8ao7ieXGp/g/IVI9N1tFpACsQ7VNUcg1ksALm9Cg4fLTEdaBfLS2lIWQwVAlWN
R68LWcxAOhzS071WyZPDtmjWGkS9H7t4prSIcBtliuwMM1MG3Ao+ODBNqdVp8V3C
Fxgv7x/Gv7npihjf0f70zr5ZGlZjkf+/QcneVIU/A4EK6G78YM+hTjm+vHCqwt9z
MXciQxJ4l8IbWjYV9TM7xlVgmD7zaCuq5Imgac2Jn42kChK6Dv49wwmk2bMrJoPO
Qeuk7dXHjCRqwMtsXd1Iuv98c3MqsbZxcdoGc4rCmKxx9Rt6CbJLmZO5ciFliBb1
fxegHK3Ib0yBlb4/3mPEt5NQfLVjv1/8wNcfNrqyEedwZIvhMzjfYU0BwpV0rkS4
ueqpqlIb7cvxl7Vx4DOex1P6IABfGZJFQnpm/Vg7Q86eUAfd/35GBcF5XnxAsEqM
H0dp8lcYUn+ltzlgqnLLatFkKQDl0reUYgZvMJrAeRfxIHjtbpUEJ6OlPUleIpkt
E4es4MRwo6m459rh6fQO8URcEHvuJhFyh4II/G3eV+nHfhvaOfW/Nj0Xggq8zHv5
frhhZcTUKglxqskA/kYQKvUybMyQ+rB2K23vKHjZlRWuX1gfGYKPGbx4hIUfnq8F
JRrkWd0oE3dOd2UU+tZGsd4Ssu1YpkUrpwyVC8QHmzyFFLMHTlWH68eOXuwSTfHu
Rioj7FR8mi6aC0JK4z7jqFE3QD2mKyCsl10W397XF9fMxht5gs4AZ9Y3JAEl+10/
h1s6qNDEfsZQXZsx9qwHPsSGRkcZruYMMKgPEgImcSHMJ4LZtObhNFYRUD/3EchI
z2QCpVTdR6Q4aypDT8NqzsvuYcFZcQcK4zqjqeZUxTDyfGudCtwBwj6rRRS8eCEX
E5mAFIFTLIFjF16+pxjwBaJrn7z/LYKqBs/yd2Ot8xvIODaOuFFHgadB69N0RGMT
AhXvETJb8GneaomFnEUVOlwwWWmPBDrHxZGIX9oaVaLU+avznIxRwkCltQH9Anpp
OFnWYOza0SX1DVhrneybFiGXijFusyW6nrFHlwTFuN5PUfFRvw7OKnlcfECSI2CX
QVred9ZN3wzvLWzdNZb3H4XQxEXaR35KEcrrHu86wpS+rqp2GLH3p68voWScwRDz
88vulWfUy/UgY+UfzaPgKr34MvA7fCC0mzxdjDOBGLssIibv4NBPjcZbk/dJfR4z
DQaAh8yB2UFi/arn6A14A/0VdINGCJ6SBAmeZZoLqEEablvCvo/ZjFDKEtB/OU8A
+eDoTp/TQVE9BZX/IyTH3FlGQmWZq6JLEIpqh84N7ESaw8v7u3lzjCqHt9vwLa/l
yZUksAKubyKtt44uMNz17eq1SLIn/lYQsewQ+gpQFSZa/z5XypcO1mGdxQ+b3Bp6
x/K91UcbRFxsaAeon3NtkByyrZXzDdUdPa+roUFDOzwQjthlvcg+FtKQMutBzl9D
fo1J69/LxKRdVsnGKJ9kCsi0w4MsCNuSBxZZyg7ZahluHf2V9cQ2lpIxDmUBP2iW
UEXU8ywTI/jwydya0DzCJ/uP3TzYixCxEdWE7TJutLjkO5Q5eZwNIzGccWkOwtAQ
j2a7OkJRD1sBO9APmsBEcAdldRBG8xqY/XObqkdT9Ajf9t2/I3iVsQn3cZevhdA3
gkrLnMg3vK8kwYUqI5gjft9RtHqqy7EJxPcxypONeiKybNgM3XkJRaR2q/gCvuTN
8y5/93QWEKFCvqqenwqV496BgVjvOVC0XzSZztJjJzujMk58rxUcurjjjgWqQF62
d9OgNisQdq2EhkrHb9gelLRmrdPJEzRmYT1jEKlF2Jw+l1GTsVbwRj30gGWCqXbc
ZGghKS/PHpKvp9niI6X5D7kQr6+eVbOsxws+YMPy7IyXBmyrog15L0z2GgkR7sWG
Gzazv7TssPvEoqbp56iDYHsQjHuEFZDBvLZIimIe0kGh24tb2JaN1Agz0Ome8I0V
+kXewyU+k+rTt+ANeQs6aGAUh332UvbIMAshO4QJ5my20AaklOdZJ8j696+PhU9i
eMizfi9LtrG3gzVpGhArdTWt5pe0d6brZyI56uycIbkjXEDxSoTKa7ONzmdFUyuy
K//rUV2mHFTKHbGmI6WBDyhoKwyEcPCFgsKKSvGaq9LmPw6TgBGmJyd8zi7U9ssx
x4K0ajdEc8nIZ9LF5zs4OTH13mu1Foi1zcJZk6wF8/A5C5iVjn3qlrIRsuH40LFR
Q+hcyoh5Bqg9za+K0TlVoKWtRqCB8EMHwKh8Tvzl1Pj3kOQ4rPIile6c9GweRwLb
mU1ZXP6nJGMWZeKpY7JrKFHmWiy2HjsP7/Ms/3yVf8pXYDeQGj1cK2l6e/FkDehA
g1tcxnlcI4aQQhCPUeBIR5csOrIFPnJl7oiYGo6NQX02UAxFwCmYvLpTofl1ZoKs
E7xocXDT+OC+hzf7rglngyRjPWPeHzGMB2NX5tgiiD9/w4uaDdDCKi/9QpVeIcFv
nKCZf5TywDiiM5BN+oJvasP6ANb+muRGYHB71mXIOlxMrAm1+kXPGoEXruMmrzZL
UQ2Y6I/LAQCYdwRwSY2KEZBlZFF8WKur1XY9opVa0k4FCrGFe9S47KJvvSuV7LFP
x9EyUmO7qNCTYca57zh7y9s2opd3FdnHm06xUK0x7pXnRnV1gxUyZhsDLNUbNJ0D
oCnMnbuBNgEM2Q9CPg310uf56jNasSOEEo6fxB9X/YMbI2bfnLeV00Cr9VoIjZlV
J/G2jOsOUfry5CkZguVPFoHrnNY20yN4RMxyltP9Hwz/GTZQK8fe+NQrFaUgtH5W
Z6e0TQ3r6oJLoLmi1ze+aBmPY/LMykl+zbOGactAh1uAdTzNjW1N7hHEoWSLr+b3
H3wdq1ZQA5fA63A1nZk88vorJpQj/Ql8jAop1ulIqsWnv2M15RQHd4THiwWYaY4s
8B2ZoHKDU/bouBZ0VFsAUAKb9gSmkB6wVLdriudcBVQRVaHBA4wMYVrqBf/a4Vs+
sU7WeZ58aIMB8xnRtUUW0XaeaieALs6xyToF6MWIV1LT7UcOoCQEjh4F7aeL6K4D
XrStGGqv7B78aoJc3RcrIn/kCCQFc4V5fMVidxyM71PU198N1gdpAUVDR55IczDN
0vlABNXxn+GRGV2gOwhhmpo+p/qzVC2rkvyWamqzPVCkUv+XJZ5OK7UPhspHnH7U
/XHoN5rvlsmIE+mt+v54aAVKY9oPK5RLB71JgxsBEost9cHOW0YjaoiPFjazB/9v
puizWGwGSul9CK0Y5tygbbZ4/jNTIsmwr5scydqhK4oVmBoYvaOR16No43tzQZ8Y
89IltM/JEIGk67R7nNJtGQpQ8osYZ2slATkojY5DtXJlS0RmP5EXsTBxcWEfG/Xg
zkmGymfc82Bt905JtkViYDwawQG7VvZBSrmEH40dLt26OewpLj91uowoNPcGsZFf
zsbkVgns5G6hz3W6EQv+hggp9p0kSzd4d+uWhQnTVXbfvMqZxWtD3Dx5aGiiZwLG
ZT30K/+8lfGY9YZF1vFWCJlLFENGtiWQFeWyiI7xVnDLaX6n7CTRedWHtsl/l9tk
RlYYTQLXOEIrJFL8N/SJrChptjAjUlvKOAYqGD9jI5TGeROqOlb6TsvaOBDZ8PUG
JSlZvyaWdHviFX2H+jfOzZ71okxmNDWNSSezyKFgCwFxi9aTCpx3FRWkN4XctjLl
HZ170txYdmI0qu1yUPxflVal3cCyRomGuYspcRKtAUIk6kbBOjCi3KmLMTbO1YaA
HAmBEZwgK9YAYlcp1Adoq+IpwInARVdGnfAf1QlmC4dZdW0VjzcrSlH/LYD77Whn
3EHTz8uPEYK5DWtsWdz+xjUm0aul0hpJfrwmQQe/UcaHulpENiN2DnS3imZGCt4O
GaqniB291oCn5HguhyhBj2VXJq0xrLSWGOl+lTqqFoxoJeVp3VoVW8k2dZADJOFp
HFx/ISEdzQ/wglJI7v1UaNeIl2GSzVet3/UmyCoGY5OJk0ikz7hl0isZX7FOR5sl
bQWDMflffqkgPuGAZAjAylnFvLACZnqTkG20btfokx8hFiGehawZX92/igUjkP4K
MiDD3bJwmRSyhrgxmioBFtwQgM+Y1+GrNHwy1Z/1atDx1TMWia5volxLsDuXIhb1
fV2+xVwM9Icc8tk+N4bPXkKaQSAiC3OLZ7g3OHWUx6PsO8ld4iG8IbGoY+W6cWB4
Ivo+DiVS/XISfGwX6Lmxh2E+e3Wz9ggxESU74OBSBbe3kprF7F1pREnjHtaTpHUk
exiOBsY9iqXEnZfBs4yYf/YvGevX2jeoqn6sKwrue7AittQyzQFHONFzYBKvcC9G
J9usYEEx3Kv4UckKRoNztDQ21ZjfhyaTfa7MhsMOnAXCDGbl3+srlTbaX1JvPoXs
A+r/mg2+y1puOzuLqpSzhjlYwYPM9M+U5ifBkWGDH7x/4JcezjgqlnW/6aBWJLFS
bFEO/2G2dO+A791noo2gkS2z59yP74ggmpSP/u1TsrKudsRJXxK2oiZRig/v3hVL
vy9Gm4+VtxMlhAP0iC6OUuz6YvY2enPEzQYAiGV4m1NW1mwT0DJY3QCMEk4bOpLY
0JA063GLHO9yn96RphKckT495Q/tHb0KViaS1MnuBJDHtZy5Ykqcgro6RJvq0nYx
0ygAmjGJjqKbzEj/FaOHGn0yZeS6Zzo5/ftPC3p61j7TzKhV1hiuvQL6rkYEeiN4
DI4Vw+/pQx3ilcShuvScYWZkEAEfcMB/rI6NRK7yxtC416PkypzXtrF8OAEn0WHY
vd66Ci4dpcRptQz/DDwTElVE56Z+DvIQ/3uQdH+Lv4/ILqQ5nQCiU/b5ewDv2Qo9
ATwtcCkAS9Hf8FQQ2tspCeTiReQyIQkFPVz3gZ23L+80DJL9XJ3kAoqgkIhciwzp
9MHDXlg0icT8oqG8RgSHULr7utUla/6ZR0D73b+EgB08Yw5H8kIOb2lHl7O5jk6N
GXMH7Fmae5+k8Z9XND7uv/vZULM+iKNxbDGoZdxHxZqNfmkSSDiF+BDIKYJ9vKbx
25nVazv7RhocRQHYYeD6ypT80ZivyCFn/idEsk0x9vCwPBxtGVLdxbSTtWDzATaV
Qhlz9F6klf3qlodS2u9diNehSvKUqGTfgTQhez40iUorAdEOMaEvWhJz7L6tlPvm
YCXg2QhTKEpJiM5tvp/Qr/Y9jueOVOXnFNOFx1GI0Bb0rfGbqRtO/SkNtYhCu4ct
X6tHiPIt+3cxt72U2hEvYa9LUIIad1S2BCKRy1vWnhtiRAj91YAltGhtRe55BuAT
LK63BaWUqe5hlrriRq+/dswCpYno2vWZhl5cnj0WyzlX73nG2z/eBdylIZCtRgvh
2i3Q6vQ/hskgmhJZu3ypgpNnEFFdUG9tkGCBUaOfJQHC8iMKDVVrArtOrS61GMiq
+Fbh5JmatnenWFPaxng7CNUxmUkUgZsKu+DG87mdXLJd3P/2MFEkaIJCSpN1LeSv
jO2f97+bKD5BpfsUYsXxSvb5llcnUJDmWWk2IRIJ/XQLxZd4cF01Q7tqjAlMpGid
Tf9ftJ3rQ2X34j73We28egt8Z3AqWr0kEfHC7d28XkHXG6zVlGfSH/Th80ehcjEV
e6+5xcw1QMKHDBYi2wMsxZxGqJb1Sp06XZfs/OOG3ZIZKoiTGDvOHzCoCSFw8tyM
9cyqMuAkR4Z6IxP0z8Lh1Ss32A32i0IHJ1c74kxwNTbajcJJ+himbgQ+rys+pHOu
QkBsj/l2M8NvfShmRvhWx9OD0vL6ZMFQQVKle7U08lncYpc+/mcraMWRkGhezon2
OGbLSjg5uAgmPhnPkqLq8bJGb71iK/c9/lRlzPTS77lZ1h7pW01Qj0yuhHRDXydJ
gZuFyRLvPfuotlOMW5H3yRfVoGNQQGDXHQRFdCWDxyr8QazogyONl4gPaGNY0pAF
T/9VhjXirLW/wQCGZdrpPePt2pAAZ/mBEf9T2ZEjBYCBC5uicZlHfLyrtsqzPHKT
q58HEu745yq38P+sblimVTNthxpZiHFdPjHC5387O7Tdu2D8JzMeIm96+MLs+E95
5LQpxDvAFNffeNa8ZdBkHNkK9sznvb3OERiS6wgb2p5bxv+KFF1/MXWGyFRVsHSf
wiUSguQnTkYr1makD8mxWM49dnwCI7wRDEEbgC81q9sSBHA3vdo++2mhtbNOgGjB
11SQsR6iyM4VkZEZFIxgnsFHQXFPECEjMxnOqDHgp2nYul3Alychpjn6oHoC+zdU
UUMotKJOXvavjWiIPrBjmp3GjiBQG4fuMe1dOOrfiow+9Gb7PHfToOY6sDs0OxLX
RAv9H9fFRiwHAt9M0+v/HCIWYwAiq/f4vlr7NmxGGzY1XEQ8bSYmIBLOLkRrsNb4
dMoONED2Q+RzhoORxcba46YLmb33GxAx0gUlQAJujqww62ooXyCir26heT3TTPDY
chWEx3i1seEPRw7p60vVSRY0YRHlnutS3AIqoAWo6KJ+pdKoQbgaPRN6cQlfcAxh
/zmyAz5+/zDo0BMSasXmKObMZX7E2SoO2YrRlhMhJqOfOjwuIEMRFcmYWbhNlywm
yjCTFQVd2nVfbZx7F+TXXU110RxEg5StzC+aK0nzyoV137oCR6tQCComUFUAlnNl
9+gcEB4kitUvlIwcSpvgv0RpBzvbAqtuONROKc0KVBcdAoLYbm32/jes+m0kRl/n
8DHU50sxwV3Yn9KGHumbWhkAyJ/A/iwcm0jqSVEtIkq/e5ynOhLtQo4r6B7gkQRp
xsZm4nZ35lLmHz6EIeP2PRddvCszz1JaDFAfI+c5+ycmqhC/baUrGqWoNs2yDzzu
fzow7pDujDh1CVS/IgyjNbPkIcDxER/znS9vxXX7W1+nkGDj/VvmH1Foib7oAl29
/VU6pO799cYFYlMe75fcRjHCdpesHKa+hyHW4mz8LJ59YqMnigTApaAJq/jyF95F
yOQsq87Fdk53ha4yKZduaDvDuTkg+8nY4Kf+SkCaubdcGf1LiLlfutMSELuaYmg2
wCL1df+TQ+2u0uHOSOCO/1h+35XaNTg3S5BdNGNAKoc3+x4tUmBTBMDgivgh/RY+
aWQk8qX2qWwECk+5ISSbLtAkDhRWJ7I9aeO+/p0RefMmx3VggGR+kX2nxeylFWEt
/GNOTDZMuMV9Q68+q041mZnB3huPCu2XZDO3QvZ0kxGCsvxUX9w8NTfxI6tcGSbM
a6ATPagH3x0L0Mqu9pLS880quDiXSR8wgPTdlXZmXviJGFRyT0DaZqDEDTTTZQqJ
CzCvZ5nLCvOjBxlDr/EwpGkbCyO/OBBUCITBc4XBu0ayCmn7260JMUMDv1p1hQYM
z63ZS95z/O1qwkiKN2gjumfRRVA2hXOX9Wy4y6cN+okmWGz2W0SmxEhw0FrEfm8y
+TFTlNzhDE2N8srNd6rTMuYPsX65TUk1yeqsX71YU0iRGqhVpQJgbLMbP6QjpQxW
uGfQqxpSO6CMV0V0FCf0zaP+ns11OIZbgFyCRthuBI9rRqBjrxnUi1VjibU9clw/
Q4hPRhgToEheB2hoUfIs+1kS4BxOcPWqZgkdb3tHkD0ebGM+bQCMw9CS/xlF6TSk
BCaLdpe/GI9Be2QgDsxELEb5V0d8kqKVU3C+BUgnDelWPyd7u36rhEW0j2DS1SYK
qUAEojNPNESydreIjeFbemw+WCfx0bWIKWtO7XA0OTL2WjOZQtJjPB2CprTlah6g
loj5sMEh+OwZMv+Cf8UkN0I/MKMYSq6RcqZV+wxk7PFhwvxWRLEv3O9LR0bj/gYo
wm+uhOErrXJztvt0BnxXynNU0KP8bCUcmtdyXjFoeyiM6yRoAcRJr7wGzXOrMz0Z
vCBwGeLyrEgNn3VmUDE4WAoMo5LLfyissEDmo+l2uRLp6AJu17swJffk7ycFhQcJ
05wzC7lX5IZzrnl4y8Kp8/7P32nmw+hQ6Uz7I79PX6MxBT4xxaKBGHdodU5wMAfd
+grRVCf3mr6AgOHz9I5OJ8DP05gy/P+7pRquEXZbKtalutPtEUfNLN2Ia++Nccu6
Bh9xrftA9navrxDkMnoVs47rR+GMXMFGpUT0a4Uz+3h7G/NoP8+zfoPkBDaaKaaK
+2Geik+2Sg2rQJc9/0/+FWDFO8zZl7VjW/REc25k+1GxmRbfi8jKg4564mI4wXd5
oUgNg6ppenFNYc0eO05wMD+/d9/O5PWvqkvcHkUC6TiGOQY5L06lOM6S5/lnQ9J5
kNCsshZ1JJsiUyP7BmtaoYl8adwo44ZP+iZEX6VE12jh+wcT56f3P13wafrg/u1i
ZpB4c4Aeq89RboLz1Pn4nZ0VbUzypQ0uaAqriuxwNH+yzGOtIwBV0Iv3YOLwbsF9
OoSUxsqhNXIL0YYTBBCETl0uBmrHe6Ajfmr+wvt8v0tec8TYM6JbQaE1qFH2bXy+
3UvvVj1UBTw5qhlzO1OGJG5AFnp0J2ZtAx1GqjmmiVFvbejsepcPl0NqRtArlswR
Sh+IEyrzqKsxuxI3UjBNgGOsqdMC1oeM7trkNKq7kCAvVOjeBr6lrPA6ZnXGFKkk
A5JDvGpGo34R7nwc/i8akPL75Pp0q3NH+MfWocs2ZfMaSel1pHh3mv9qJ6o47QZB
OqFHLkHSmu1B8rE8MFIb+eqhZPUOT4EbF35HLGFh6iVeltrFsv/pZe+olt6ShxRi
sq4AcREmgz3IxLjyNso/19iPmnJ7gLQvcOZgvUjhCw7IMsoZY3c/dLzIACiH1yJ7
4LvP2FdCC9939gsBap8ZdDWHFRAoigf6UvMp8sHo2CEp8VGDWK0oXeTKSn0DBptL
Cb3q23kzwG7JWEsya2PDB2QPnszk7OrImGxSOEnIMlEOq7LOzJxyI8vSvj57oqrj
A0JhTMo+GZ/1DK1NO0pOD0PBwmi+E0IYkpgl0MbKwVLKna12GsLzbv+/cKtKpfts
olSLiRePKPPugSlRnYsz7x1ACOz8kGS2Fz32T1VhL7pWWqPaB79a2KbWwvwduX9r
KpypBWe3G2sdlxozCPT/HbtE8+Ggx0XAEU/192pdMh2Sjvwa3/BfQxJehXP/k1e/
QtX1ExT7z+q0a0bYBEXIeiEn2zaVmQINBfcz+2Lpjo7NZadMjG2johvftDFwms1T
dqc1Lx5YAMc5015qUkFWibe4Zs7gX+jgg80yy7rEiZAiLasSf3dYLQUwsgIBpm+q
KAaR99W4AyXztrKVIUM0IrYp4m3iXTHpnoO8a//jp2skaztibKjQvVsi3GzCaxOT
/aWtVDwYX/NdUtlMG5ekJTkcqma6k/nTqAGd9JyrivPSyVhQYxXgI8Qz0drXIpUH
zXsxuWrEpVCD8RO9mrW3goZp0ffQAQ1uNv48MryXr7AQl0Maa7KsrrI8QlqJysrb
qg0dJc5oxmdBisPYqJLKUz45kvzHEc1cGvFr0ssMGmKuQjDu0x5kgASr/2qx3k/L
jG4sqaRoVt75NRxe4NEkvJQKtHdnF6m5PaWGgHm9ONjVWaIUTcBsVFyHSCwFNZ54
WSssZbF3zHeMJldZstAjTPP0my/mh19UNJOXq2PN408+ZR22HXHeO4/+NAkDPcs0
MZMI4/O/A/KQbRVFHGR5iwaYKx8uYnLK3Dq3SkhmW5upMR7Xiq7Kqm+16YjX0rXF
7E4MS5ZqtKBDGGHLKCELIbvn5XwQCO4KRDUfPu1+q8oeaLpwowG5ZjuE2gPoi1WD
vtiVXPMJj5LyCEiEO6nnjkLSfu1M1ifqnKFFeAtQztQg/Yl1lVrX7Y9ukXm7UUu5
MHZA52r8g11yA44r5jnBcS6ADH2KAxzsDGMQiKeueKGVw5xJyDincYlHGxe7k3Ml
IG1hp9WL0G7S6sWkxF7L8c8OxRqzpNNpCK67jBhTuKxju4bCWlGYhV4lDt8k4ekj
LdSOMPHM4DcnNP0OOtjhGOLKP4P+57Fxs6W+i6sTkTNKjo2iQuf7WHe6AwMVhUbK
G5nKaSIon4lDECu0pu6gBItTMKEjhwmPV+XU55wihprN0Iys026vqPDRhiPcbp0s
rGur01pWv26tEWGvMI1sdNBTqb6ZbloGG073MAYhn77Ip78a/x7f/7BPFSkEvGTC
Z+suA58zxDXvFXFtn5pbNwqmSE6KEE1uhhfqHJRoS4AwkFHRy8OXFIL04q2V3B3C
NvL7Q0LIc09bHFwjphukRDtWRMFz5K+6pVGBQjm+D25SYitC26WZAZkLAW6pN/OJ
fez5QjydkjnrydlZg//O9a+4Uwe/MiRy8LTB+Sltahb4ChFHjxh9JScQO6YvGf1D
uFwhNDyJaM68MW2iQtyDzDvpbBp1WnWhVL+5PmNQpwziA94Ng3kIXAYbqL4KpLDh
lZxIh5NP6So+5Izh/gJY7XXZoibznLftUW4rgwXEJ5YvONk2ZvkCMwMq5Uq3l5xd
mcbS6CWomgMBATCs33xNCMPdAnQVCsDt9nAlDFAF/Upms5+4LNdKdgRvHiGDr/nm
6Z9uRcdoFrAoEJ81Rrj29+QZhR3MAP9DTvpiHfSRbWK/q8cGO1apaVdSBu2FZ+0J
R5rhDZapwlCtjPCQffmKhgOJPSCECtzYSi9X775ZbwYjOj0M2rZ1mV4CjvTC0Hgy
AGnXha5ZK0kfbse+/jSxXwHQkA6eQCktvO3GXSI+pZvs+AgE2hrCYUWrchDrEy8L
+8zPPuSBQB1ee7VBPVNT4Aqm5SLCjuNgVw1HIfG24wwB9udE+6XOWcGDRqUHokAJ
PrbaDgiaDraJkbbzXTqJidoBfujtmj5yuq+G0W5u8AdxGhv2exZyfnrlKrJmCndC
XcLhuTfaRor/vWDP4gD/Z1L0dHvA+dwsaijR662WIOc1ZXiKVeaiuqSodNBEsfsP
yl3gX4t25eIPSd1l3BU8HctU+IqQ0Da9q3pd2E/JYyxk8GcZBnzWmfA40nef5okI
v0tXgfFr1nxnExlRPyeuus6NEl+j8uwvq3/AvxJCcvI1C6+5PAt304M9ThsLHXeU
Dmw4MByrlYI/PVBF7oBvXRFc0IDsrGiKnhfOmGSnYVTlX8sex1xYtlZejP0FAEVu
ns2gmMj6QaKicMiJpg/nyCB2FHLGC3ltqORJ9b/TmUQEUEy9nhHBjjBXz6e/EdwX
M1DUZy7DH5T63TRuaSvmYmrha5ycOl0vT4uIfT3rbjbcN2eFbcFnTstR3rqajtA2
Rc1pCxl7YKdlmIehhOwKpmnXXwHsWOB6gVlgwjzI3cWg4aKgJvPekvQd2WtXWNoH
2pMHkooAlIAaoS+Hm4GEtjKRK0vgXWjIMhHuZ0Adv4ycILG6n4KEbpRx5uW43B0H
9Q9G1NX46llUG4p9oyhQD7fEWtr6+ALBvZhUjW54GppExEyYL/L1ALePCeTNNuMT
n/2760SVINfhdH7IdVQ/9V64XwFXITJXEwzjufZhdOLpL62UqWYTGqRZfXKGn8+1
8ZPsnxNDVhShQuhPFRgY7jvrS2yLTBEbb0oAQkzAdYftfAirSfa+qXHJg+o0n/dR
cyrEYke6eG8NcvGOQn5ZdAUlr6yNkZe1yqoXKPJ8G7leoTMHg2NtHAZF2W9N3Dww
FMmhRAoFNKThkI4ezuwW5z/adClfoUzTtkZ8DQHz01WGkJinpEEzdV+aNwOJAPWo
pIOqQc2A2uhgkbrb38y9czSMo2aDR2yYSFgDPgwQVmt1wk7NjhsGRy9tZvQ7aziE
OT54JjnVGwa/lyOwbPmZPxd0p9L69pNIr0EYCSKfHKF4igiv+ZvekjnNt1HuAVKE
8DMGWQUVJups5/cse3h1V+VybqdsncogsAuS9jeVE3WF7T2ZzbH8XVIYqbVUFCi4
apuPxjsGOVJjQ67OqwCAJwUsFVzvzLPyW897k/RaJP55T8PUS9vlWcpI6N2/zfud
siyhH8fRB0Q4z+E+ZLOFC4l2cC6CqZ0Eb3o9x9hYasYyI4ksmS74x6fV6IPDlRgB
COuLUMdmJCotnD4qc+LbhO/OjmJJDtmYVT5e9OFsJrax6+eDL8OneGMbkGu3c49q
2isE5L7QwVfx0itiSBBbUFSPU1ItY7C0hLWpdmSC8qGPYdZ9hyo9GGh4DBvaZlvF
AFITYuaEoWAH6td2/oLLWZl7uX35DgkRwU2YnVFKRQzztuqnW+eTmt0qajE6Qcjj
v20pv/CvOTwy7//LWEuKBNIivrtfuFgEfqH0wC4/e1X1vA+D2bx00AABj3p3jipq
CiGaulNiXCPllwY5eowVGWJEk1AuwJllKZQ/hnqZ+q6cILU1ZMJeQQ3b21hw//kf
O8A2Xq50mWJqTwJjO3+Ag6s31JcVfWP+V7pqAI00m71+yneTVdWBQo5dC37+BkWf
IacWEslqpjoN4a2NUCqWTEjYz2iif7wR1ij6uw16V12huI9YRRVgtqdzPITpLp0F
agSIxHEeJ1r5bSCY6/0uZoR6wc/+70yiWlk4P3OuSu1uk5nFB2ksdn4LNqq/O5U2
N2EJ3D38ym6HL5whr+11F7Pvo2JhksUXDPjAs9K0ME9Z7TgrwMH/b/gk+CdY6BjW
BHfETVxhm6KiI6bvI28NrF4XcP/fW9tUss40TuuiSIPVRx4ruL0JaatN+S6pwqYA
Oa+JLcmozahMOddabfKrnixQ8D6n0Igg7mI2y9wnVoVfs/jeEFbZCFfDg5A0T+Fk
B8f2wct6VB+xhOI0A4bTYMYiQJ4gs7TaeCW8ILltxBoaS/4UK287YRjOT2d2uI+X
+XThlRTmKOq2c9NLgycW5O/Wo1QQA9x6MoEiXKrZv2tOkULym2BnVHySMsXigJUk
ctueYolkd7SsqP9svef+3cZeAgQWfg4CIfstB+g9Ny64lFfPmE285Yi0eHklvXIU
HSgMlchOCRakiwYD1rzDmfanTqEtJM71fD2jSgMz3fFA1Zrbukk/4p6i/OYHk0Ow
JtKjoDbD462RxuF6UyV7VMCj9BeSyCeh0KwUc6y9G9RQPvrjuRLqZ4hBEiYQfWaa
1jyqXx9j5zPJH88TEdPUuteiFAxPy14HxblQMmjEzWpd2AIN0DHPWDKHvknx06jg
juzgEep6iutQTYyNONYyU8W8Pl0uhRMqeXEdwpjhPFGzoS+0lpS5JQ0xCitOG+S1
hqX7Ttm1VDK7t1qBPKC9hdSj8IDs6+QMoeSn2r8AQrOtMmXj+xVWqT10xtlAXwge
L1N0lB/JtD8uJHyLtCOXV4ZfN5Wc3o/vuSZl2QVHQRkLrkPclBmkvxmIG31g94k5
+W/LWGvFnIvrnOp6Qhk9jL11Wgdpdz0Q8i7AnGcRpikL8QsXMB3559Cj/3AWYMXv
YnvrKVRPh5yj5Rgd0TPk8rTJ8z0NhIn9I7yQJX0K7gORJpXZcN5KRWYclU2qGju0
z1rnFL4ok+tbymNf2NFmgl6p7771IFx1CEHsxJNDRf9tQVANC1X+cwmRkIuqSgwc
SsbHnrn1vjKshpNXNepeBJONP6fA1LbykofzlK7ikMUxXGdSb0TO4LWIhYdZ95CL
/knqKPTa1pjkGstkikpuHLrXrPv2SSde9jNcSuxf6J7/IBga/I9JZOp4yapt9cGM
ezvRWwjaczgp9mla8O1F8Qklnhd3W+lxgXTreU17gXAEXgZiZLL5hzzOygIM0aBN
aMkiXGuZuGzmJhw922YClkFPDW8vKu9Mh0yGxQwRBmRa9ysc7AXEQUxSIsIJ75Rs
XjLSei20LwXswTv9qB/w3I1qSHLQfpC0YZayyAqs0+0L0B+hO9M+CRp4fTqgpprn
JSUt0yun/S26ckySbV3Uxp34Bnyv0K1jYzeuc8lcPKsWFwieYb4yGiM0pXtO0Ofg
4+6bSwcX8vtus7h+lWbYF+JpgpdCuGC69IVz9GAyktyQguK1SjrqeqvsYPgEBacQ
RN7dbL2o41HwhXx9cIlYutRDEdcCWKP0+OfzuglequRxLkP2rwUeU6ZChXAwo0cU
XDWDpWMhM35EwMQlUhS0D2TZitElK5zH343kWsPUuswrlXp2TYvWAWtqRY4bl/Qi
Hax1hoZ61uHdnIKIOhGradnKs+WqhQbXDklRyz9pR7axjiUoU3RLuBhUIBMblFL5
CsQu4OYOix1EIzW0SlAUq8Nmfff6Ix9FiYLvbCvBHG4OEDXcAPnURxQ/ypi2w2Ir
Ow2xx16EtUFdsPUDRVMnw3LK4lgeBjMqC+nRJnxND9vg48ocMVz/PfajK/intLJm
Dx7FvAIijevGR3X+ipo4NwtF0P76D24E3JQeOvbjVJcj2K9kWowUX0mkcoTxYsZj
PErErMGXYDvitgB3GXOfRpvFjtoWSCbiKOjMU+9DvIdpYu2CSNCraRTDwCiqVrVR
hQxqmdZzFNNiEuYOyvJo0GT6PaUVdS4d5456BZ6LFrWKF+MXQ1K5pInaila8uLuP
eySHNhnQ6JJm0/XD8nEIHYVjd3wwucU8yjnCzjvgswkf1HAPMe1eNzg1TJ1FOAx0
bzjC4+SIFaGuZqAjr2WH1kvexlzRcKLEcBYZQK4PPSuqvA3PbCT+GxSOI98Slq5g
C4lzBcwG3YN11uEIqbbFarAZE5mTOoX5ikh4auWYZ2+x8FpodMT24PNewUTI8juW
sG5w/s61TalruEYqWYqnA/6k55OsYozDG4rRB7+bXFLJS6KW9kq4HC+mvSQJ+Bd+
TTc0U5TVj1WmG03BeZoYVmB/Q8NxdG23H0111gM6i+wNlBPllUyfCKk7KonlGXnr
tvMPwQKwuRI2tHfgfNSxYVsn5LGH/w1gHhkDQ9RPTnTeuMp+AeC3vevHBnPGyZNf
81Zzg1cSfT/kAFwKM3jplWc6Wjk2nzg6v+l0KATtBBFWddPEWEaN4S3UPPd+Aigg
WXmO3osNhI6AYavmTCe+5zsU9Y+SvREuzPcG2Buusv490LmJeCPjv8gooZeN02VA
8mH8w29UvFk3XsQazaKNXwpVLUgXrb4bBWyrDPsnZGN2tVL/pfba6lYNsoH8drtC
YBO+wK0bJRGhGofsGu3rtf/UEi27QqDAVT5rbpESNgZb4VjmtEGacxEP3TmvA6X5
FSgmITR+l1ncoYPeKb/KBqUkSBjXlD1mAio/w/mLB4WSDRhnSBwhiGSMDq6bY3Sb
SH2JeKyOSa/zWrxcRWihtSwIG+G+XaYwZFBEpZ8/gsIKxTY9wtyPRq00VBjYfHg6
gybHmuoyD6LaEU4l8VSmuBk/db/WKUF3tT311h3qYtG67dOcoVEddh1ouI1IKyQ+
bvuAd4SS4Yw0iLJNuMgah7HZzMlwBPEyhzwulYFPDFslSJpp4XIg++cHJk3Xh/J9
uj9sNcZuZpcDlf+p6LySyW1eZHyEeGQE40nx7s+42H8owhWdRdkd5mteClirxytE
RrENUFaUv3OFNwQbF/t9GYLMy/LtiVUQ/iN+Thas+uYvg6Eoe0IlOHKICo6r8uqO
qmzX0Ww22weg9OM2RCT3tixX5nZCXhF9xIaSA4AyNbCfJ7e08C4HLvM0ytCkWyrX
ppXmd6KCGilvf1d1CVcDUkBL9hfC8yudvS2a7ao6uXetLFhDiLqk3AaHqYavlADK
ikWX5pX62xRhLE/Xq2UTlB7Bssa3gmIsQzJqn/X99AVPZfkOW4JkiGQ7x4EVhhkF
vmr+24HI++yaWmoi1Ve8Wy9CRkVRw6iyKG5k8bRmXO1wTGY2z42F+GR5kHIP9yJ9
Bf9Q+bmV2kz+1AvI/okVE9T8XE5JHNJeYaZ8M+i19yTKgsJxFaIoOab7CIF9i0w5
wxcWW7O+VJUlbtvgEELhUAtrbJ+PBNiK6ZuP/E1IubZbea78Kug+78PRgeSKbBSN
BTsfTK5JBdC+99RTrQB8W4w6IU4VGrSsOWvR+hC8+eK3uaLpzm4rYrgYc+ITGyDC
OE+tMY9bN9RZwSNZKnL6bpjrjmBlUDXRfiCKS4k0+X8Pp+l2ZQxKt/oingAfYZ2O
zERHKrPFQajo5TxyExd2He7VT2G+CsDkZcfOwsCPsUDHLpwisXNA8nOqzoKrPkwz
x+DXrv4Tvskvfp9fA8O+f03QeBoXxFCnL9Cuiatvyxg4HyB23SCJAaHOr65RNMNm
Yd9ZkwYFHsEUjT9GydUp9dc27X7AJddBqArtUhOkYPrAzLiaDKcH1Z+vN0dlu88s
7gkmHYWBc7V7pxmLoAQemNo+gHH3F6G8jvuP6qzbiQxJDErYpezLZE7QTfCnk1p2
23bt16mtnriS8u+d/KhYD5+HriGFCWmYNgp6m4YuZOX2/RwVZRfngVCC+vg/qIKX
PBuQpXRJQEc+P21XYog5HJRlcOv5UR0hmTDjQO9J7zLO0mCscBpYW+MtRSVsb+2o
5lug7YfCf++KtJz7Iy0Gqh8Rc5v5cyLz/LfJkRGGn81OwDn569NZXmHmJ8l77FFK
F0qrILOg6Ei5BIh6zzrsggW8gztDAK5FkYlIEO988Yr15ssLDw3HgkZljlk2BHww
bADfrlESqqwcnFhEqhO9o4eXYQIlYSlJ9gtnytChah1xQwRwqYHE+u4OSBZlSGPD
At7qS9ssmZ7ZCsnXMvZwci1aE8kv4XAxRPFHG8JjzHX63ufrs4Pk+b6TIz/FQtao
QZW7nFy++tkrLYL8v/VLmEt5RySR4xU+TXlaTbatPZSduQ1WW1RN+nOrdPzCSd7l
vmQeO89Swi9BOZa+YxE+fBSwgryee7guAXzxPbDl05J0iJ5ETLpnYj2t2csAt0zS
uAOUqRLzKdU8G3MJxvzrwheT/qvLmfnrNMugxcFcDnYPZQzhPVbAcXe2wteKjzXN
kpXZoEn5ON3MbBI8P4PjWgA7bL2Bm9L3omHd7h5LlrMkYBQuABJToT2XiRn/D6Wd
nl/BwQR5+0Q4n9gJ16hqMyT57JhYOBMDD2DvycUzZC1bQCKMb96lFpNm7E2SyJDA
q2r3uXyepBhYrftgija25s1aaPLskmditzZ3jo3Ln1LHoLZrD0pEP8IBy+Rl9LVp
YJJOl/Mo5BtrGj21du5VhfAON7wNZa+IiQUGk+Ok0kh2IZdFDB3wGkCpYh9PL4HR
d0Bt40JkjT0QRqHTCQbRyAadjDyCoo1arWueUdjPM4veID83hfGOZUwo6rxjgOCE
muSgV6sEWfPl6fqVOPcX56kFj6CWiwsiCtEhAqoLHgmdYWstwqJKDMG1uFmOVRG1
5z2ofjFVe8Aisju2qg7g2fD/AreNKr3DEq+JyDd4F2YkzkrUeKb1TYpDBHWnzxfN
FL8ZLjIcMl2vjTE80RLm2PKTyXuJsnAzNaYCk+X+YbJ4lIPbjfPAl8Dn0xjQ2qpE
QRJCbX+oMnKbg0jGKsPspH4B5uaR2fqUcjvsXx42KzZZ+cCFeyQDLMBqwKIb3fWM
hqkrqsVypiNZ/DtSASZ4v3RlqC60pv75CO12I7csotkUbpC8ViJII6kNXI/++Bjs
L36Y7WKgvPZCFARmOhe9anz86imfzBn5nWCMLxjoua/MtLW0eqhL31KEELnlo+BD
Q+F3ui8HFHr7E8mHts1qpcBWz0vCxvv/QaYlYJYuNsnRw3wT9uq1Bmz/86NrPugJ
XElXqSJhVDD0OYx8zvj1wEq5h9aVMs+aK96zbM5O2uaMSMi9ZJnzqyGMxFkO3yjI
OdajrjiFtDxEmbOfC875saue9lCqyUUJMwNLyr21ZiMdoB0cecdl0W+gvbT2soW0
2+8Awkbs20SRyuiSqny/lEJdae8joe8UqXWfGwbD7SZV2s3YZV7n5R3PrI4kU5/F
0VVZTssNeN7ksHIfOon3FXsodwN9fUNs3hL1FPwmILMQ7EFFdr4WxnLJ/iK4hcJX
VGXzB0Jvzy7FTEYSQWrNhIt5ZK5FseeWYIaBFsMNZxHGIDNdKPRe283IdkOXC2PT
LufkDwNmSuHiC86bvdbNw+HHD2RDdxtik/gZI4SZrvYU3JrhMvvQftK8JZfQUKcT
J8Fz/GgSfpU5FTZFiJBlpOakrY8JILbYLDvcuPeMOaf7qAEnk99AluDRyHeMBsnO
Wqw1RLtF9C7xJaAidCjs5drfQzy15OQ2Cce54eSv5t1X5BZKyWtN5C7CmtYAVVw9
hjrKS5mQdNdcV5xq96XiBLmFjtLQWGMyKYBsPzwicnIAc+GnZJO2rMV6c8bIbMiO
ipHOgijyTwEXQmYto4PebdC8f9kPJnMhe21P41IfKE5nB9jWYMi/F9v/XvoeRVJZ
+z25afIZr+WwqWk2kvcL19xdR6osgpwSnDsLqtoUM9uDOxLvXOWV3aroJdHnYg15
EFmjikXG9RKrWaoSEO25EiyHOMrYuc16i/bDkLC7YOUYkWj6XWtgWvxVu3v3PIlS
wETfwank1b2y0Fu9odSsMMC9FVO9tDylqddeSc+cs6wPDbZDZXeP63434uwT/u0V
Ii2aFCZFJOkP9PMx1xkx06SzHmXurlSyGo+Ugmx7jbyvOXeAkUYW3kL8BV0QyIHw
isM9KOxtsS9XLIpi4xRTPGHhOROuAgZZyaeIpLssc21iZuV3dnOjt9oKeIFeanHe
kK8110VJwdMh0XOacggjAOoX6VwSufXB5CTSY8Lt9pNvsAEW1kEOaMZbXdgYFliN
KA1R3l1visg+66J3k78//XaYjffhhEWnhulYrwf3eUhd8FTjHx5pPgjgNfF6dCR5
df9rUeBa7k54GbMF12XkwpQU6swb8c5O5ALrDlYoDrkbgCBVkcVcI1M3KjKqWtkX
oDJRrrB21H5gAjyxnP1tYNxSTXLj21dPC0JjJCbmBaN6jMWFGl/rGFquNfPeWWJ1
tNP+W4S6wMapH2PL1kL1GTH36o1sKwC+MCyJ32TWxibxBKyg8Fubk76Ixvr07RhM
5jqcpALouX9NpCQ+jRzDLyGfN2W6LowIzr17UcuSSCiDGlBkbNsUh84gtvz3+v+d
t+nKXc33/dtmJJercNY74Ds4wPUC8spGCG4xg/F7azdIgHPwJR464beTsqxfN9sH
0eyb+P24ShPoQnM179LmYpWscYQBDgpbJaCr9JwN33uFuCav+sCAm1bjwEVAxi//
v5Twfbyj79VfBuSLvvFH+bFTVs8SMcXMEIMnGPWNey4qWK78qcOaYpNWuosg45VC
WklI0vqDIO2vHGRp1AfI63zTxgAqL7npDUf0zhaLslPoSCx8yirOetvsPdjIJ+ob
qwf42xDI65zzY4bO56K42PCQwyLFtz0jr8B9C/AqKd75VcXmWq90LUji0usUtnCL
2Q4aEGPc6qDFYanvRHTwBhCcAY1qCP/NMfOIDrtA3iboYdhCqIkJTlafbAMOHqlp
QFRiGjgvQXc12tJOg6kcTNoxCyIbg/O9jyXgiF23emWmM6KGV4eQcpcRFB/XUxGJ
ntWgP1OEFkGBviVxFZ9Weu7r0hsv2Dqk1C0ozpPIDDTFh0JoBR1MmsY4aiNTX3KC
1+yeETKvYMrr2Yi9cmCayTinlQK4/WVGPRYMKu7FvRRvvLoplX7PP0LT0YFmsqKh
36qcD1TYsltSWS7eaFGbw2STJtNJUBH8XVUsLFVdVQTXxHt+kdlRLjCuZt6y36/V
b4BTvKT+JqZ3jJ5Yb42qbOP8V06H6PTQmRUxn4PRYBjdILiSl34gUiykGS8mT8YR
u3AXSrCWMVDUCL9JxvtboLU7OEzInZnTCOCu+6dVVS95x4Q+F8tFMGUH/cbbV1zM
J3pA0gpMV6w+RRu40TcImOOaas0IsX9al3cZEFOzumdouU1c1wLwTotA1lSHFUWG
2SNcPeTWrSe8zNGmLZAeXSZHMSbZ57pAA7gZLzIv/jsXkTTSt6ATKtAZNDO0Kc5H
gz18LYZtg/06m7kxHID6Gz1XQgod9knqFf/C1ArnbDnbkdiLMYbYjHB1OgDBxkWx
a6DqzLKo16zBmJClzuC1s71y/ioZqeQN121PBQUXzPS688lfYrb9j/v+Pc+bJX55
dxuL+8m4m1rsOiTPhVmQOmQ5o9SJ4qR1gCLOkbM7O3wrgsw+7E8MNPMjI+TyiRsl
QNwgWJrEwMt7+1JPxl5+TWDekK8Jy9fs3nFtqXkhGNmn+FQkBPMHNg4NnZIdOoFl
S4Mzi007seIcemNVlHd1Bz/ZxDy2KgYReaMoTgyYGJ02VPmEXmxGweluBpQkS5Iq
PHnsK6emHYdtbQxwiS5sHbAdk/xdDnX00oWSzBI5QgaCCkltxaWmr2ta5pWwSiDH
f/9Q6Qwax2w7FA6Mpx6O0b+VeyscmQJtm1b9+kA8CMUoa5CxNyV63eUmycrqKKM9
UQfnIPSGcbRgafjNk8zf7WeerXIqIjprtfdv/wuM4hrCZ3ERSmfJHo+HLWkmvoOP
H+rVxIXbcIhxj+t42wkG5oQQc5mFjN7JgkqO4auOuzJ3xKVup37DfI4zxogLniSj
avxI/T5csP1wOgfN4Fd02oGaiwfMaUYNz0ZBhrHcxg8irO3ADeR5GQpZcwernuDu
ccK2w8J0lsNPIXoQwDz5AaC3423tXIJeaETtjjCqORoC55en+50ch+wsf9CP+42/
z3I1veDhKG9xSWVkAA7bBVKDEPGd0itbIjmnDMjc3aceJllQKppqajfXfC7qybek
rOVM1Pj+AQyI4jFIVSnUMjpTNswq4JrevrDi4GSY/VukOZ1tPahuewEHvo/HxbmP
3O6q5oKoJAxr5P6pIdIS+bWQWy1Za2rPwZI1z5ctH2SyG9Mf8ZiRZmbgy7ePjfuX
naBovrCk9vUgmxy27myXA+Q3Fe8WiBqgh61Y5o5RaNu9Z+XB90sMzjBqGebWutLO
wVfK8yHZjOiVlgOoiyvOsyQuFa2NvWEpildVeAd3GcanJdBiy49/PP6v7QCXMnQ1
+6nVIaaMq7ObYD2QzJMWpTKc80dY0mWERTLb7wiPYDsOp1VWkUKaFcTJtM1+VKun
rrIcQ1A3CnF5MmdNY9CPi94ZrXZRGQgGTq6xApURbgYoHmmuPKejdBgnFeq5XmM1
Ev0AXLcy7v5gCNb4jLn5r0PoIMxLbnLJdV7r3Aek2woUH/WHHWf4VFWJfYV/sE+G
aFAct4V2OHxGMvRy8q93sjlTUK5Hx6h/zuN4kZci/9TFqKr+G4diVuPBqGl+Zgy/
rmtvOGWr2AJT1Lc0DWG0iD1Q2m9JvFd4XOWlVZr8NyaDC3CI5V7MCSDpFmgYCMo8
kmPun+9b4M9yHDs0/fmGJXtnrDiRc6QbzWWawm9zBYXIOKTeoDn4W7zmghl7D+6U
c4lPCE0PNWHaDHDxRK86sf+GGNMGSyuKrBVo2x3/kRtt5tB/degGh0oyQeFn6v/q
mVPAuadNluPI3nA7DYLkGxrJ48XidIwmBLaOvstFWzSC6LhWjZ8qicgkWjybPT03
gmEnHWifCpVCb1YWn/aE+IqNTeKap3AFShvr77YWMlN2SbJEjl7qCRonPFLE4eJq
vBSK0AMCEEgPWxRV0VkIylx9AFplyGxCYWsJD8XbuhTPeY/tLAZfnOMfuM+/vpGS
v6PcPGxXp4Kr7z7TZFYy+0D+Na6q41V9GetkTvcp5dMQN63d4nLD/QY06MPU4nrx
3X0tiQSmk3SIDEm7S3WhfBHo5SXxjKHy5LMD54weXb/4lCkEFf+Z6RvbfyLzTRoJ
982SKfajYnXweWc+yeC3BExythOMKoBFTFG8A7YWGU/26CV5hq4iAjF4h8ESIFFm
W8mEAF1o677IebUj04BEFEvykHtePrNoJvizo5lvuPjssqpwhZRRAKHxcgJaYDnz
Z+LjsLgAMSfexSO+6euOaTzpnqxoCl2ZpYATpIVDLERIQTqtfNB2W0RmKsbWE1vy
YIa3IWqXyDoRsolj9j37yB7vZ19REHlfeQcL+aw6CFTF5gGSDAhvWEKE3QEw34Dw
lGUzXUtnKRoRP2S581mF99I48NMMozg9JET2CMQf4Xq7uOUi2FQ/cjs94nKmkOye
iZG0aRSxm7leCSEsION0QVn8DrYgMUjU6sz4q7vzFVTSMp3et5LGhNIzhG5EohaK
2WT3MJGyAyWoUskkk0fsGuI18Aqj1MzNvbnuXBVcgX77fyS/8uxJr6yourLbU2O4
bGMz0on0GVbIZZGa/pIEhnQZ6DPfV9fqk0oDgkYR1k15Rby2VyC4KQMyymsJ//S+
DZC6lwZNpQcTkRT9msO+f6XcAz5cEs7nOXq1joQ8bTGJ7FhBQLX61WfY7xSYv3+t
cVsrs0mw5NLKguxew/+SU+TjqAtR5B2jNIHWWiEdmDeOzgCKypQyw+ryVzXrx+J6
htY1HEdfPy5pzOpNeYRaZCfu+PTi97PV8ll97b2lzBe1+c31n//T9lk017ttztsc
bruQYQnBhbRDtLnNtK2xSlUwVvHNtqikzR0teWamhQjH+8xtywrRpwCTLnoREEhP
MjGSLwiOfFfInFMbDccqcjJ1ySaLHCb5MqNIsJy7kiphu93qmAiSb6t1KwwIJctD
I6aiVSBwJ7nzzAA8wAwXUKd0IpWq23T+Yu9McsHlmWttCZeBJK4xBCDWTNchwYLA
aGfVDcF65s0rVjMp2gqaTPta1zOV0HhryYDTYSrpY5/gJz//5QZF+LE/IvXcmXCI
fnSivUmU1R9jLIjdspYURrlzEIA/whhClcZi4xoUmiZcPcm3Hv0NxvUJRdoO1AWL
vGMZvG0t0r6blFulIOZuFQ6EUxT/H/BN112pFG9J1lEX88xmiPpelpx/I6j8e8h7
uLUgHC9LkpJBgCZI4X2du6rnY0Pp2hs/TAzwGhgocRD4Q8V2wsn5S4/4YrzJEiyM
TFHGs7HthggsWW0tbGhASgpr1d6PN84BFw0uUB/dP3IiDoMD2qEwPhey9dixMzn1
aPxCQ3XvjOZhFYYVa1bys54OnO3hi42f7quPiSZ3UgEbK+LW42Ns6zS3NAbbr9ZE
qHfeJEtjAg/ES+GRe7kqkcMuA1GPMcoEmC9YHxxG5iCMOF8xy1HQLN3OzZ6GaIIh
S4uTVoHM2y6UaVFD6DPss9iCDtoe6p/o0lcG5BLuhpqXK/dsZBvnGAeMRtOPFgrJ
mYubEWKgnpg8ed2eCfJ2HcMzIDudpci20BcnK47q7ovSSPRX0XQaT3utzwv8Qpb0
D/+JkfN/1o4WEKCY24cx1LzXrwoZ0tq0CglZtdqLLVZH+/20La33CJ2RVtq9n4RP
s4krMzdnXR2CiZDSvuFsNurWQm/fkLHVkL6xURHma+FRMqSvNF8FBhfzH972kMlM
+daB0236zJCqdGx3iF4/hVl42FE5yCAnPgot5YDjEHr/OilKEWr0bUwiGAfnXZP9
aXt0yBRfcsTSQxrS5w8d7HmrWOkvskeLGEg1FzC/44d5aRw+LOOlra5ugB9YygEB
Pnn3RFeFA7wK+pNKIJKNWzf7tcBvB+hQ90BIGbt4LW+J5OlU+NLPREG61WGLAlfS
3pxz6nnuPdl/81pnRlJ1eXCX92fDOPY8/NhiqbsHtYdwvs/0g9jqWyQIX2ncUCQd
yNOz2oljnXreupFou0nyG2IvmyMcpQfbgGgQnlQOjoeXChsTzdU3Qimo7H1bDmK1
tFaTCAJbo/ZgIaovGRCHWAnaj+VWwkASCp8BdYqMfONGgCNwmtJizUBEf2LmN5sL
OFZhuVDbhFB+RiZSzs1bUs4Pn/7RrSAsvZ+v7kHFz+MvSVLwz5LzsAb9gjYRtXtV
NHhIGNaQFTL/xMiwa+vjaRyLbkyduE7tptVPX+c6Xbqyz1zd3dQqZhn73vsn+sck
XT5OoNzhfYbJQ3cX4YarttqNGvI9bJuUnyl1wS5h1glA38LBT7dS+D+lvlmnKj5d
UfBWjJqBig+Ci2gvEY+i0C6rkqLg2bCi8e9tYGd6jWbROX59wTDdHbsNr9J45vcE
ajc/hk7pYiMLA/2A9qndJBfjKN8uqfwa/lwNUp5wnKgrKor+XKbpuC3A2j0WM1kM
v+6bAEJ6U9R94rpWK3zmDcATO+ZOcJJyWnVy03hJQuNCsr2K3ByUcKBFtxjwCC7c
nlmg3C1fKiF7jSf8QSpFVEwsrPXlY0HfdfrRTGLyHVskHp32Cld4xoAGaKw4kzIc
Q57+rm+4pjoOnQ/phO224wQ5iqzrKK1hNBS4xx4ck2AnLHyE229iCkWewv+/oC6o
/SSx0x4l8mveCYMQuVlydIxuGzOmuTx/D6TUROf36dnGL0D/pdXA1S4DmuTcI3Wh
4JxXOkmBOUdMoCYSBl7yvftxiCk0shjREBAm777ojQyEzxAhP17PX/Gaag9p9ubU
jKwk+Gk+ypHf4dISsFpLVQ8fk65TYy8OUqFLDeICtu4eqqlNQjwdg4W67A8Q/GkP
tMPRWyJOto3d6BLY/qiq/tlM5O6nNgZsFJJAx6twNz2GYZJgjJle2eOCNjoE+6MY
WDcBOv3iFgasppCay93Ony25tUmPW5SSthfxe+E6YNolmrbrVP02OtFTSav4MpxX
wPfo4LEPftVrp/ij9lNGfO6JAOmdWfo2M61kenApPyDJF8wvLf/wRl8rlW+jK/9m
mkFI0RLEyVHV87DnaP/juoNM+gZz/USpQmmZFlhIVk5tLxDGQ9Oev81vypf7FHKP
mhpOUt2zXFnlba8vi9MjvC9AfOOpR03uxGxQc6M6YdVj5EWjirW749MTTRhLwbsx
R0JueLlRSRQYW178I2C5E7w56gln7HyRn14Aba5L+ibPcac7olU0TIRuMMQlhyn1
1J0rCC7zTEfCsSQdZB2KKWkYtLTAriqBazhmQ7UvzX/P9OXHuc3WFGvoF0eORB85
YBeCP2RvnpYH3Taj/nQfgkYiQT+mC6k94n7AGlZDLogPTtVdDtF5MmS08c2+ylOy
FmV3Vebz46qIn5qN4avjc0XMj0WTkXNSLxp1gD9PgXIvdF5eiY95nUrDa25osDyB
X8llLpqw7z3JA6SFzgrYBFBOBZewF3RUbA3W+bzKYIg4ihxGkoAve3Rvir0wQ9MA
iqHIqK4d0gmrd7T5chwMhBvxAOdTtVOc+qYJVnVl3gml/iHBkbB1TqA3fB07uFu+
iD/erPqzO8Ya0JwOpFatI9mpG44MLBK1RGCGJjfRYAnI9fHYVVvwAWIf3TqPy0fp
1L2mE4+ulLFiA4At1HHF4vF6zjidXRrOLoEtVNZVldOtqBBMR8oGc+UHyX6+46Sg
t93Ia5G3jin4dTOw8miyQ3po+MgwVNTm5ul5mb/43mA0ChV8X49LBwNfj4Me7PYO
f+RAS1KvUEZb1lO5oCjI9NKuylErjpjX2NmEIu9UwZf7lbLuTCGmW15ZzJxYG30z
Y1FoL+LnHnYoSqXS7/A65OOb2Nc6N92M+qGetF9GB4vguOasBFIjf9jBR9RUTha+
elV03D1HXi4+bO6vo8oXB1VZwgWu/eW5XeapkLL/viy3bLb88hl7bsJLAllLpLNx
vWNbmvTeXwVcUDx+q8F6SBxkPqDHyzEL/BZtuKBiLERFJJ8MF7jvRdRLuIVKhOpc
VgF2IrwMZKGL3CX72aJmUKDXDpE8k6VtgcD0ZtnPcqxTSVRCwggw3ndDg/VGq5MS
bdmmVRB5h8BzPURO6372O37W3tgy+W7dW1/H9lsDaDcJKhOLzeAp7kjrIdyx79zh
TzNwVl+LLNZ7CMY9gFL9yYPmSAuxUr24DYaZh8LzAgibD6IrGaCUqQA87Htf0bDs
GRd2nOqMltBhHbTSHU9fXg8r3nDVXKHxP8hH/NM51S8Vo/2psyzoy62veWcOJb1y
1pOkuVFKweTvymutIDaO5KFzoOVK6O5+P7DKdzb5EIxTmqIXAhRlzFMiEnZ9jzwU
3/vsoNob0mGivdvCmxxXGRb2Eu4oBn2kJ4GZM+7hv9STb8BpjvYhHHYeZ1/vQEzX
l/TgJjlFmdr6LVU0KmBAYauNP2Tk6SpQKCYDMj0nytYez3rHOmt1Jq+81BR0y64F
MNvrebF5uF957VfYUa/v7BVje1zCPcJmjNEZLWeyRUmxk+51GIY2oEIsoXxaxOA8
l2xZ9LvTChw1HotKEyDFpGzMl1kwZDNJzW4w89DXc8CEjdeEkMZ98+F+2lpjtrwZ
XhWHKhn+A7UodxzvbHSbnCpO4YjJ0hIssYexd8TU4qxJBQ3VsSIYuzbXbGvLWpTg
jrWOOBpe0LcVyWD9HWTatJAxdgZUGrgjhvDWzv1DmevzyfUdDaxoysxWDpJHGctX
LN0MuPQn9O1CRCFdzFeKzhTL1RKNuWlATWpM7ImVtK+RuPxwkHbXYK6vfaLtr81j
T+B/d2D7KsMwwns8nWPbZNWzoPwDw6UqbFbb8BJ3jFchuBxgtKCMUuCKj/4waH0/
j3seLWTmNYh4UD/clyfvzqHi0SSHac7a1Ys9wpUWfyMQWPcUHTk1l9W+6dwevut5
rwuE1xm19VfdznMK5nzvQMsCMK4BQh7EfCy08RP0PHhuDAJI8zKE86Bi65DQR20k
PbRgJS+zi+5AwLDlbXuUtFtZCtqb0cbvv1TseOJEWkrahzuehUTpqaaCobv1Cso0
ZQf9ZPrEgj7s9ACDBxE9iyDsH61zBFM9Re3/J6flAurZBVxSM8OZWXjhW5RM750i
i+WpZX4UILw3xKG+QGB2MLbQ8gQZPdeqxsLfDMoWkAJ/kqm/ap+41ND27cw3PC46
zbrXpDeoV542RUzaNY3hAKpVecZaSzgpPzTrgPS2TdygcQrn1URFYzXI1gIdFI+i
3orDRz4HCMyg0CCcnAES5HzlC8sjHq830TTjIugnf3bcPjdgsf1+onLnpqxOKZbW
V3aMYR0CGyjwr1qyh3EFtTPCx0q0JJK5kLCxgabOsDqjEW6SizYvLoa8RrAA1WqU
2SHKLM68cPgXIse4SwWAUXWLGh4z9CTz9d1ecxDRlfRU3yYxHCZ1oKHMdfkG0ABc
jIte1Rz+Ftk4tUpR4LKBfl1ursn0XFbaDk69sRz8DqJIdVzPPlZvD2WjqZAYcdGK
c8NDsrV9eAuIf7h0nJRpEk58SMXNg545B9loQO8isNF3HrMCiQwDV6ZapNWHBLc+
asIGLhAvILyNTI994TGBSO0mG+8/ikRUDRZUoH2E7W88rICutFC2rzR3IB1Tx2lm
5oRmC1N9EBTpdm9o0PIufiArEnqGDLrrQIoGc3LAxf03ExcnS4VcYhN1+ZyF9zZo
homuKX7zHs+p3YALbEeNs222LHrgbZmp8MRofZtNv8MQGbf6bcaAHEhcPsxfdBmn
AYil/PaPPy9xbCmbbSk5i3oocTsfxQGBL4Ri1u4nO5+lrgeuY9kaP3+eaznrHFys
1Bse5LGLioUH+9R25dlZknOYorfPPsIjweOdCYf7Y3+yNsd766YlFAx89qU3He6q
PiyIqGnTtdP3R7/Fd5P+5r5n79p1NNQOzeggqr6OwTf00xoIgj9A9z90HhjXj0Wh
14MIYnLqYn6itSsdbgdHsAvbSJPPc6KluuHw2ZQLI+c0HM4wK9sYlvA25fU9soYQ
c24Ii3xg1ijOtxTvvYLd/wT0jr0TxoRyDnI0OIv4Ae4Wj/u239vxuyMyfSRuOtcd
mk+Bg4E+z17JD7k9n3mVp/SswIpSVI4oLDVnVncVvDwDUyU/NHsIXwKrypolCP2D
/FfMAIs3rysn6WjIaERmpSwg8UJZH/5Krs3nFI0Fi9uLuZRiak1fhvQqhr413O14
8H1N/VQ/O5zkpcx1tUfaMWM2d9lXzgoqdD+Tt5lRuceENrVBb6/Pm5zmdfmbIAiA
JL9kh4F+BAsPGzKyWLk/VCkWhidaIKFXj646yNPp3gncqoNeW7LE6pf51ZI5Y/da
yWqMeNF866F0qte9X9y+o/gVXs1FON4Wqi54pB/lNqIAxUUJF+thb7UGLTbn7S0W
stmAq03/VHFmj9scBmuO8feV9BB2ITt9F2lrOik/0Tf7G8t5TbcTRBQrxDlw99+P
eJQxqpq/UfXf4NX78p+cDrNnpSI/T45En119YAeekVzTC9I1qsnxjFj2eOfShUIQ
fw4jI3pO37JXTwNSGakCSo3aAPOWpy2GjGLq29Alp9Pk3pbWoDPF/Vp16O7f6PiL
6EW2gUaGBEdfn/dGap3xJRCr6uLPwo4/I8FHPPl1e/AQNwPoJ1jHZugEv5lPpWuY
Whib9SKCedLEUVpWiNflq1HN0ZDefbPVPYTu2y1RLRJ8h+tx8Dx03CLNJmYcImQz
3Wg29qERdOF2s9iEFEPVNyaCJ/QJfKzISUjeBPrSze5G0rZRdHNjhyCuFukkGRnA
SWzA4qHu1llNMJtxOYDIVu5F5pt9xlE93z0yB2UxZNO2RcGL+f22F2GEjaBjxAkk
tEP0KpTwLzQrzHMBAT2/4J+A7xyNujoJtHJ6EweOIgM+x2Xy46OXsbF1eiZrMi15
9CpN6/uFUxUFem6WKnbPhonUk12mvDfnaxiXjLeKMYgt7GdN5QtI1nTwZJkfQXR8
1YhPutT7kUxDs/sp34WGNrLpYyPPJHZEQUXj/T89HAP1+6vlbO7+c276f7bzxFlu
B9ciFsjsw2P+UoTeIGtTanIzq4I0IwSc/I2JBa0WlM8d7zkXeWuK4TrnmdcVUKe0
SJOZjerbbJtjLNIV7LXxsnDBXjzMHpFXB5Ed1ibMgmeIPVlenc8mvCN2rYL4twrB
B7hOYefqgPSjd4ZhGMZeh7b1LEt7obsMWgbS5+R2LqkOe3ll1meD/i9kXJDbZjHr
O0DNOI9oU7BVfng4ypfOsVm9IlWe3EySS43CtPeJzmW2KgEYcIZlylym7ySw2bHh
ToUDBVd4vFen+FvTX3o2DeiNWHbUw02kjGlWATpsBRhoZh5SJY6z1gD81UeELIM3
7R8O6t48eskL7xET5b+0JpzgPnrzpousE4JIq5Y/cPx5KM72pGv91vHOxZYStKAE
/eU9COOy9iYXPcQhzXU27Ju6T5/x1Bm/ESoHNKfpHU9bL5D0jq2Lc8YzwQ2Z9XVy
2pGxnTXldqLD6Fopsv9lghIZodMT7h8AdjC9Qhz5gglOV2seDl8QMJkVT0no0VJh
K1wqpkIQrvyu3uhAYQOU6izD79Was4EXq8o+gfXieU6g0a3nLGoolN1UkQii+QpL
S5e84MFzx+rXeGYKrRkM7QIGNSwZltUyqgRFFyJhbFW/pXYDFxyjgzN3pk8tUDa4
4M4vc3R3ESQyOo2K9lKv49sTr8/aU2mfKzAdNgV34J7PGyEUVIZeUMKJqziyJenR
dqMSDULxvsuDXFbN6e2aEXYn8DNn5WF62j7KXK75DNNHO5XooQqxerW5FC31Tqsw
Gc7AUaqfjBIp5CjiPeENmKM1HDo8+AW42416gvhzAZrESRctXMd/aPz07Q2a6i0g
jBaLjJ0ko0+X53qnndRk2GtUWGJDwtvxUgVgrCQmOrSi4qG+ad9jSpsTkMSy+Ph3
xqXrspMRnPvaLUupWjxAelBuTriHallRQr587xfef8DLyFEC681EX5XDXY5bX0ut
BxHgRN9eUKZmIz5Vor2z5uFsBwL2ZTz43UeC2HqNqf2NxxZM8oK1I7y6bni+1Q4h
5ofUVas/mfqjnaxn/eTl97i1CzksS9g6Sgc1biBl0X2ibeZ8MjnDMeuEeOscsuqL
+B1lNegMKtVjAyL2Q6EkQTtWdcH2rJ1deNCo+kLP27+SZAxYLoxhYojQb9NKkI/F
13oGjVAdwxebnoZxZfyM3hVsGE/S3L5P3GxlK+Key4d0EtG5/7IOBAeLY5T/3pJ5
//Tbd07vzTdwazusTIAbjbnyeiSsR7QmU04cqk0Saq6k1OIZAa86FY9xlULuTrts
w6jSoqhWWoj02pa+JJiQgncLyZJmJVI5smJIufLdDAaxfysf1Gz4lJw8WACW2tzJ
Pfo6cLdDxyhiSuuqgdbAaHRJucWia4/xo4wslt4iAzUX9Rx1n+pSLpRaOnb3fpyV
2rTWFzpc4u50G2DBsAKRNX6cwAS//y7AVEImWS1UypZ5wb0Gve1sqXpH/1T8k26G
+MeB0I9SPh4k4/QD8/B6So12fxVRNHK3cmRZWl5Puy1tZvyKTKUoRWu/ybmpmIJa
0H2UffP7y3/bzqy/dFm/DJgaOZXFrvzkXAfJmJ3Dmzn4rfrdgCUcjFam1jBeTlN3
qTWA9pM0Yu+ulbfTeJF/t+3XGVqeZnFSSWjhQsSGxyc73lTyttXsIRJZojh3CN60
owWvN0qSy/nmii8/W4i0X1bv6mGDZDSCw0b+rHYcIccpe5/6aBd9/He+O6Grh80Z
HGzvpJGg0X/Yd5rDm9hae+DDYHqibQggy10EJvL84e9anEKMRx4Uv1l3jvUYzVwN
HNCpthyrzs5d5FRTd4yTBeDl1ZrfFkKVl/Hx5wDNnMfH9/tM1RcYEwuQweZ4ziXT
xHRyOm1UvR/e9mKJt6ZB0M8DLlUoJr9oJIPWpaYjhZVtekWBGeswFiowtgoPRZpG
n06TpDKn/2qgrGkKs02lwB+FauRuoVKnQG+4amDvcbWgaLD5iuhRN1pg22d36ofU
jaAfmJEmNt4zkKNRHFeX8sMzkR0Hz1DerpsUlmMOLqNts5X13/JiNjgivioNLvTF
1F4TpOj1DDB9piCXzeNmy8/+0MKdicCoofUZWNrKENvnIrejn8uz9SvZOygXjHY/
M971cmiEx6dAvy2ibGaJmjNPfJLiBsO2Wry4BaawOyHmbnP0B0RqB8Ozq9IwmmtJ
nBhhmshs+nM8ZsZS9DUjZg==
`pragma protect end_protected
