// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bizkVxZJvYVJflxRHxk8ailoJqaqc9oopGHmc9642pk9na3BbqM3Qrn0qTXccYJu
3UgkhcC3DBozXKgzCEUJT0Uh9iOFpG9LWLLYE5cLhK9PDF94BLzT3IY/cLCIhfko
opzFpFc1pPMQzYc2ZxeVZELWCDPnzfodIySag/leM1k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9840)
4oH1U9Dtr8wzlfXU1ILcHeJ+AQjRY9JFCUBhNT6SCcWwwvGiC9PYFO4O2YFFd7rk
VgjIG9SEHYR7WE4nouOoRCt+4rsWrsWlsmdtg8hWr67634Wlly4aszw9URdZCSWx
/CpVz85eQrZLWsqosHL11Uz4Zk8eZVeWyOnHvDVvc9kFr/fmsJfqcgL3TqfmDWU4
qjlCChbHeTcKfFQRbfcq5Ezfjj8lKHIMdSACCP6/9GtMEpuWdLCALwNUV1nQspuL
ervud0IGRaYB4qeWgPJtsmWWay0v9FC4v6Zcqaom9Wdv/B2S50+hSRtuKCnI8Cjz
qMTOy8KA7d2l5Ot9V1c08O8pxrTVl6xVITyzAkAMtPlZ1qJFxeGw27vnBqpu+z0/
EQhqvb1yAawinz2OEGBn4xwjZGYnsaUDztb9hyyK/w9eF5x6HyDv4y0Q3gNvSlUj
7xiBAgMQeEarpUyKZFxbVXt1eabJJ3TD68U7XYP4KJ2DdMdaYBopS0jCZLumKlHm
JZh3CrS/3qPQ64JCSx1YE39eff87BFVIv8oxcquw7ytTuYAR0UfbuY74gcejNtS2
w0d+O7FGEs8/EDK8DODTNQc1Ya+voenVwvXuGwbh8U005DHsJ266e5LKsyhTck0S
zfGmpRz+oJ17cow+8+SYxeDsM8JqriPnCfbeaHQs+3ZsLpzLQUTBJyKtDDgxERBT
8ycvUz4LBTHg2TLKCPaTlcOJNaA1/dPv5urpCbF+4ieqNfqB2C9o1ah8uzgFNvL+
7+KKRTzocaF6EUnK/Bh4Y0zVP/DlIEtMZLPsofv97UVfSPtJHNGF0/L5NRpBYyiJ
0RrW8zoQVBUinKw41gJRCDh7ab13LQc4+/tFjYBiEvufmM3ptUL44iNJSEDmQ+6W
oshPoTM2VCxZ59x3JOsRVyjz/r2S0BTSBNREuS3JaSM+gIS6qW3hJ7IsHuRsvamr
MI3N+RG73jprmwWvJEEGAasl4DwuaZQ57KCIbi2OqPAN32M2JGjO+JuNnGF/w/Zp
uJ+FIQ6nfvMzaEJrB1ToRqRPdSJogCuhvDkDlO+mk81OD0mb/yxD1WP+gdu+30D9
s+uQv4KxkYaEOHvvgM5fIHCbja6IFzucQe3lc7hrKtSXiB6uexpA/SNYrAU9KK49
WE8MK+pZJNZaZHSmp2LXkQV3PjEcHBcg2br+ggOk2HF4DgpAKcl9mZo/tMz4Lfdo
h9yNtj2PWanTF+YiETawaZ7pYiBjHQguMVxKE9w7oBiFy481d6oNXJu4m3+bM7fi
hNaRCcUr21dq5Cj3HJO35f6RronaCaGd4+ZOSQ93CoXRAOrE9vkWhq3rvEPM4RzA
TlXfY49xpWGed2kJ7+MIjUENB1Rw2Dou6LVFHbiUJmC9m8Q14/a47qBTp9mAB8w5
2NdgubpaitFDSMxIk+Oz7kJYO6ihS0QyDIWKJcQeXpZ+huxBljTZrmu4ppoQIEfE
zBpKMPbNj9THFQfk7M8CXrLcP0jQBgFGXxHx77h73xRPb4MoesMyDqFh3kSM83D+
VDZBEQ2pGx/YNmyM9JK8qfUZXjJXW6yJCuOAjfCeEl1K3eaOUp9VlxYK1sGo7Tox
2ClSklMwKb+L4+mZMgRNCh05Mibvo868GmrlYEEjlyYKD7dE2iSMz6UYk6NLZZeb
u7TOhy1BWkklETToo0wT78y4UNA1+vYDOwL+xi9XZH0gFsLIYXejGPs+RQ/Zm71Y
Mn09+imAPpOU/FQ/Yol9bLcIdGqMpOLKIK7h+PvoS6xly1N3/V/EvyELvz6MDb31
C3ypMrJvRNHnetP+ri/uVxZV8DfpUmMHAZjXQ3dXrA2lpbH5i4WCi+FOlD0F9vtH
GXveWR/aFBl/aJK1/iZYS4J/fIHAYPIRsITDCmJYx25wwEElSqKfURgmtjj5Y3oJ
o+GFCMguhTzA07UPO0713dNLrYawMC7wCbxd/3mS460p5Lzo8e4PNjzj0dm/0sRi
hwrego2tSQ2VRgkKpE8pW8UcvyQJ3a+5hivkLv56AryEoGeMEa96+M4ACx2gwnZZ
TPo6n0cnzmhlPQHXoK7XMvDf4+cOefo4CKvmWuYj/hWEJIGA0nzz8WgW0KN8W9ex
BmnD+S3vDGs2jTcLDx+WJQZAy6uTfVkNABL7NPpCV7GErqzd4Au4J94vstOMCiUr
N+/C4nI0T1XHxPGvCE2TgEYwYDrqjERSkkBMSyCvLl+vR7dwrQd4j+Hw7Ax8thLk
F0GHLH6wPaUKRr1PM6CIBvFC6iAwpmZ8qdNGbzfa5LjFxaVo1EYHey6LfpNjFX+Y
ucrrXt3lPj0CH53FhaS8FZQ9Y1NkBz+7Nc8TPfDJH6pQJyJwDAZ3ZrtHPImOycJE
WFDN9fD9AxQbXE99kXk9X5wVPqGKUTkMTXcUgJVrj/XSjRhXor4j1kcg2T8apAiu
l8FxSI/Lx9B7dGOySdlGjSJVVRl1in+aDI0pV33gBnCp5w/nbxXn94wFSR43e0vZ
iDR+ZnjysACdnCFKizIByAJkefcK+DWHSHzTi+vBcjBN/xZtr9zCOJmnA17CbT/w
WYxKOKUb6tPsV7Ay/wB0VCxxxFrJX2SyRHxzFVyqXPhRvX2oyEdiHwieaQYbbOUG
zOR7MySP+Ay7gX0PnPGir6wf5zlKNpTh1iGwWXRNF/yaMCIe8MJWTjuRDf2H8/fd
QRosVNQTp0MN/7McrAz+UiRgT9xhNZpruTItevtifwm6MJLWgWuCF8OY/MKE7Kc7
MNTWNyvCZHYdMM5uO59Uv5ox9U0V4sGBC36867R+kaudbIgo0bRbHix95fRDaml3
fdIroWK9IUYvFEADcCOK5LcDPwa3CE327zDiW91jd4LMCITKCb42xneCWHJ3k42E
bLgzhlwVXn/xzDFj71mDQOVSP3WC+a++tPP33wDVsh8I9fowqGu+if+JcpF/52uW
MUcnPHAYSrmGHKCEG2VYcQeVXdx7nIola7bW6pk4SZGi67v+AjqiP/nZHyLqmmc7
muz+EjhHNPo8S7k6eb8TCn7+zWzzsxPdim6b7pV0NEuaPKsyGkw1oGPuFxyapW6U
O+KpWvTz2zVQ0xkyqKzwnKySkg4gaR4cOd9a2gvXpNxQDsM5IRBQuFedcd3tBG4T
Q6gdUvMDpsaL0ckeihn/xaNLsJXSyX5MKbdW8zK4tdq4Hx78275zhI5etzpT1bvf
3x7Z6MCVCDSxT2nBElhIhgWZceeu6S+/q0SHhx7b22hqcDRW2tJKegBZWx6kjIMr
oAXnGcQRI9FVBLJL9EsXKYsAY8ukm+YYNvNdevwuYaYSCxg7exC7iqh1NtwsTYFu
2BAKwEHlTlnZQ9H4WcuSxl0FyuTnqmBl5vE4RFH/XtHh1aZsTzd1mzwqDQfgBDQP
LurKQU4SRoabmN7rBaAr+NTpmll3nZTCNHylDXVLJVElNo6CM5miFOZhYxcO2sNF
EozvhO7W8fowxqLG60oxlQKKoPFm4K3wPG7/TegdDtC2BouHFklnnDyYv6mpGNgM
ir0uU2hXFmJw2VRafKC89Vm6li71iaS1l1BZ2VGjYN+tVMUiirCFKlPYIjzTMe75
lby3D5k4gv3HEN0bHRcKgrlnUnxTrce4nHzo7V5wAamEP+1CnqQ52mtD48/IbuGL
szv8QiFObN+w+XNPEfetAm9IswE/ZcBVsjWTpXbtKJAMqgSLgNtENbYstodiT5c2
LQoepQP3s8vSRuf4PxIQrBjhL0yhqOPItoTEVMhzt08cgBGKBHrRUez+tSS2pqbv
Tep46YmAfGz+wfzdp7D6Pa89guyV7kPFmVoYZsA82jWz9s7n0p5EbtkkL53rHe1s
1ag9YVCmeXHljUl+Zk6PtFmEthly+u1LsT+KCZsrA2RiFBy09CdJci49gssbdxTo
g4xFoQYekYVRMc+VLuWnwmxi9TfzcPgUJYwEqnyVXQLQ7XtR9+33kIxKbBnRoh9s
fq53MR3S/VZ1mGD6x6af8iwoLALivqU8R2DEnfbXfxNbVJ/NsnU4b5c4ZzJYAKSk
j2mYksfZRd6/vTKiqPfOBYQkpztOSE1X+BWTQNn/8EDK8JF7MaOYoof8Zl7cWOVm
rNNA1PRirLRbEajgeiDuyEpoRRrk7sJuoUn2Jrzq7VsbKrxtUKfrNti/1wrCcIBF
hVnsyXzXs6n/W5IVo+7mQqnlT/Cfjoc5/1lKOmD1oZaBy7AWAr+2vFVAnJkoSI7u
23TQPHY8pBa/bpABJZ4sdq0Cm9Q0/oTz6JBssfT5FtglgSida87oLJ8sHTXw21qy
mTz4Tflj1zFe9O7waqDpeQ2gDngpzRAHpDIThhSzUPJ8A7Gm5iKbyRw8QAeS4eNT
TTm4kcY9L19YYUV1WZ4KYy+1K/14dyw+tXXpEoTIkOkLN3MLXCBJJETtw+bFDgnT
4/RaibrB5NQ6gFZs3Ku/sAYOoT0g+l8kXCHZEReMc2iAnMDPmD/cHEo/ygyvosN3
xJyKC50JwX6yBqctk5xC7Ks3yc7ukejTAHsjWlCE5wDzqYQtauA9Sdi/7fPXcyY0
i4tzykC5VrpUgv4byKqJ6Ed1TuTU262K7XRkEB25XWjS5cyPP/Xvp+Me6Zz26lF3
CCbrITmUUW7NjEucHQI9pJ/lRp3+qWzOONYoMtJZ/4eVE+OePtr0KOSuBy5QrP7f
fBY+OS2cnh+iyS9k4cvNRcH344QbbWuO0WviVnfiz8CTGggKaO4KFEf6W7HHKZTf
r7kHtejxL/m/QHTLhmEj+rgacavrlICiAcX6E8NN3HEOPWQJtNrXaZocWqFmnXZn
WSQ4H+un4VMc7+tjeaStYoUIOec61QdLFkrsP6qwLrhZSX1QnAMm20n5YF6csmBM
2bBsKrvGUgGgmHFF+412f8pk+xbNOXlyBeEl5BNqUXwgzNseiWgDFr0u3QcCbTlq
xbsBni1V5FqY5n/XOr6f8MYjDCfJnNb6/bqWvE93CQmOPO4a89tl8LHyReQprAjz
T9TFnq6vQZIBcs4hFP58j1s6U+pkkqWj4thvaEOFgz894+unws9C82uPqR9dNner
TCRyfuSkf2DL+0YD0k7p7EatKCuxeTWZyMmUMYFMhNNMWyvRCyQCUc1hvtJ1xJim
orOYAIlN6EPYvBFsk9ukpP3r7q09MXssnbRb0yK5vJyYnGP7RlLlZWoeEp6YsWjt
xqFQdydvZ9lAWAkTj9BquCqAj619nmmPoc+N09gJx64RpoRG2zmbBPfHVtJ11gET
W5ruBmU15OOnqQhhZoJY/ezegDj9VcZA39vYthp3sAeEATmhkMe8F8ObTaUoOEp1
p61YOU2BIlkQmwPBqv7XU6fjBMAeK5S3kWNvj05JAztD7DmC6qrMaokKb+GuaPgJ
6Du8cpmN5mjAjN0C4+bW+pnaUC06TaQ1sc47fg9TltpWQj9pXUe290iJbggKFDlk
fwP1Y1X99Gsqk1xerZ/i2KB4KpTlZLz408d6crPK/1rtptTmGnVuGcOgLQUyAa9o
Ht0FhhHC5q9zV3qF/+AffTxXmsNflZrQn5DGCAuyCV+uKMFGzPLU5dlLYOclT6O1
6XAF67FHWdfLRWOWvFfDZyiGZtca+Lx/SMDsYUavC6EHtojfRnQkiNHsz53i3vyl
gNjNs8Y0FrDMvFzrlPKnSOUOHEWNZ3v65dM9xydp7R1Jzrs3JRLEL5vc8TzlzE8W
DWqy9p4DE+RYKIqzwlba6sBDx01Ek69llZikFElk1De5sxNxECWbkrtFkHYJOWNp
qIxQUkkzrOM5jKoM3gByEejYv20C26iaUoI4an77NSFoJpB3qedhGLWKU4vRwwLa
Hmr7Y/WIIFIwDNWZAt1TRI6EnWpT9Ex1KreS9f95oIzTfd+2i8HSN4OY9bCgk3rR
MUdbpuj7SK2ZVAdTMi7XbVCYiWnsqBmtQ11yZl22VMl8fJOMasEhNVKblpqpVPD0
s70qaHegVDkBUxNpnI/1ITuCVGbHD+K/EKy28Bb6UulQoBa4xiHojp396pTxUjpz
/TKqAkPQt8e+WqlRReyr+qYeJfnjBZfb9zTaFrjB4NJBLmDJ+1+saYjW9tPOtewl
OJhCxPZLQ9TuqkgUaiZkVwl3gkb+TMFU3nvPv/g7Yah/jFHLMyRU1RTohEzd47hj
Q2wJC4MhRi1np+7IQmrh0DNABZHMRWgKWfa7JlD+TElCTijaWpevA0uM6D6sCOFA
CPyxG09lCOz5Jpv1+I3s2SytiRX484bEFLsluc0PAnY75qrr1zmdbBd25GtmwIx+
al2KaNsYng2zDqcVNq1vTLE8KP+imKzpTzRgkZdz7BqaPScpVapj5jSFhY5EcENV
yqRV9WS8w/IXrswTSBy9yMB26uUy+S4yJzBklw2QuS6Io7Ofq/ULLWc+a6lX8fra
C4sSBg7lcjv7v+Zk1Qq9Jsdb4Or9mOwbVjiQMWyc0VPMLSh4Etzcn3j0gweDwWBt
6j9pnoY8mTUl28iXU+nX4R5U+JQ6kQbSG6OB2X1EqJ6Cb2AskEu6jDMuK5Z4SMVd
ModGMFlg/4AuwXKT40DzpLZyuzO5RypSzaCWshdy+UFFt1/21uAn0qGtUABDvZeT
b5KQ6wJBkTeMw/aG9k5ZOVgbOyIO5fSbQKkBb3u1Pb762sE7MOaMKBGTlLmn+2Y0
iPDdRaj0NrqsQgFYEsUc3tGtvsHTxW88itNmTnMfUFA9FrI10bMItJEOaQfkV/Um
DCkJQO+aVHumA8AquHul8Xbk/5HdzMFIoAQAD9js8fyPx9Bjw8Bsp92Y3rMOIS5J
rYM6AR2vznRShdwra9eDyAD37T3HQVcJDJvf2wWm8O3Iwhd0Qg/qhuVgHTHxRWoR
OXcAE4b1pxD9lCB0i9uN8ojzwybQm3lSDoFhcn7yNR+CRQ9h3CdOffTzBfbaOw/b
xzvDqcgYw9KIdu0iTnNPmw9xkvD1p6muyMGT9YVPIeKgn9ZqdVm20Ihp/nTB8Cai
ziU2jqi0amMh5LAln5/5eSaU3lOBOyE+nzha0es5LlxT9QkLDdEsnD96IKTVadJD
aPwGvMYQto6hoHgcDIKs7xm/FKFmAy6Cey6Rn2p2rHx25UQzf/vqrRp4PxYaFv6s
yQuZkC8vjBGeG0z4q1vwnML4krcXWLJyrsNU5lhQJLxs4uz18nxlnYuGWLIcmYfp
OC+Huw03+fjBBUKDFVH5R5DV6O86jcN875YdkRi9re5cyYbZ8/fI7lGVsytdaUJV
RW5S6eli7YWE0qE2dOOBaSLyTCvi+bhxaAOjRY1/KTdMW26AnvDsgmI/tZzLI7fc
v7us8tw54cpFDTkokgXFiqbBCJ19buY4r6K0Olq7oFozsK4UUNLZvFjo6TIQptrC
Qwa5enytIdLy3FDqstu9pIzWYdGT9WPu5cHr9G6gWDzKla9QeEJD8v8hbzjAzGL+
1KJKMcpQU2wwBaKyLqzHdcIp+9cZnl06utzcoorL1ui9TxFuwgqq9JmL7HiiKkNS
6H1tHmkzAT2p6wb/P4pxeoHh1/pulu7NWyNd45l+gE4TBCG1qNox1QRp6m23c1bT
slpDseK9+Dl0pg2Ot0Xnzv/4ltkT0tkpvCwGJ2druz2Pb+f0/SfMuCV5CRWiLqPr
4wK4As8Q+FwEJhdzLL6ken/ZdgGlUis/DVafMUog8ORdyLGiJjChHBYdJSIIAQDJ
Hf9XEseNSY0JKXeqNFk3Cefd316xWAh++n0XxSAH6pF+1/pE70O06Zw2maLwi7/N
tAaQ2sQGSaVF2fteIQhlWNgrtxZLe82EAYW2JQcq/FVpb71ZBzCEvpRjP+UNHkD6
oDeddGNfJo4aKnCEkAm1BNRMuPvW0u7OI/ngd2z3hW9ZiSp29+4PtjQGgMJxwCBn
zJ0B7WMOac1Z4xFqdUXbZs3dC2snA+ZHtLq8D5hyUc8UbR6vmV/at7Wq/grLV3/K
VvAN0W5dCRC9ERM3P400fW1TJ2MchgAjOjzOJC8OsblyP2x7MRt5yBr1iMuAt92o
EcPKTiHh1qRN/sCBtakiLB6LtB4YGtDbfreQM1w1my6DQ9Z+e/1pFpMCmC9Ziwoq
7Tvoc6yXeaBHOdUmrzLHKnTOicyp5dBgX/kRZJsT75EumwP88WjRVgw3I2Sf4Sy2
yLNaamtota3foxs6HMu48euHODyxAh2sKFc63xmpKA44zkZ7Ky3biBWmPn989Iqh
gzSUQ/dbAsAx4qZgJc9YJJdZB+u9A6d8P1PARxAfBfbhqoT9DIeuEFG4huG86Pqp
KRgWOC7G3vkyP1VYWihAP7QzPqmM0UWj1FWUbiD4vMi4YUrkl1gsp0Chcl8eJJDi
D4ZVKkmmo9fj6MeQAHMr3Ji5HwSt8ecM0ds9CrXA+36miCitynX1vPt+hcwatoTn
bC+BadscHArXiblHEdj1x6vHPwLbK2W0FaXUmH6BKv9mVq2D3G9a7FtD47BJg15L
biDtSd71dRs1u3PqzmGqDAOcasF9xe7ijEGcMKIvlb6nF88sL39p6zJ4c4GMAJO6
EZfqhvrD4QOIlAnXjD6hEuoq69c2PMSzfTyGr6GUZ7aphRDzkE0pwyrL4Darfmtl
pKKtS4nKSDhYUhC3hz+CP6wfgonqqtKS1BCvzqBUyjOw+k7so+J98SxqxcTOuFUq
kD5MQYHM74A5LSKGozrnNKqzM+Y/CfY0a701mmf1NeImLsTQvpoaq10agwyU2ktS
WyzApllrrRWfU/1ejRPxIWcp2Bsm7DjGNAA79loY9rqGStT2PYpmRpr0Q34Dbr7L
pGwwtgC20amWzgQOj9b1u8OPhx0nrzRLdwO3W7xeP1WaWv4zmR4+PxY/n7QZt76p
sgeo/Ew3NacTOqKB2irfr46dYu2e50J3QiVHNHkVulKJ2Fn2bEum0tWzNKs6d3e/
MHwKrWvSf1bKB+Ekt+kO/AK2EvHQtv3ewBw8T9EJOh2/PAAUWOzTf3WJFrdT7qXx
+OAavg0uVyyNpAOjbeEEYK/IWjMs0kRgFEYOIRRgZN23sy3RHFsmtAXkx+A25tWL
kH/trPc+c0Pu4xEzuupHslFdIPPWr9BMUCnPbI8u4YTN4PhyKxrrROmUWiOrtKJv
C3crCnx/nnBCjNisEhHoHBS1gYObay9pyGMwT0OoFO2I5yHoWdBBAc29WUArwNj2
cX5Xu4FFdJAk7miRmTwFjdNVIr51q/xSPrTKbvKnTTlRZCsPZqk5Ih78jpk+8/BU
tG10lCJ5hbq5VCywDPvA+zRFuz8BSxO1SO+4q9jf9V/iEYMIjNRNhp6HcpJ4oEir
WVBbUA2APj9iMsAJRtryo1eoOe2duuSeUHPuWp/bUj5QLHAtquCCal8edfMqmWCH
DsHhHhSifDvNE+niZ3Ba0N/d01qCjRJ5ruBR4jr2XR3B80VWUgdQ/Sg7Z6XmJuy6
11sjR1fF6HKG0Q14IRVBJfYU5FQvDFUp7CuIndBY7vmzj8UGmwl3+agHsYk9bkze
iqXKJC0K5fLemytvXMbhL2UCAz4CgLLsOhwOf4et6XGP8gmkFX8bgFBBxvrF2UmL
pVrNraQVO3dMxdR7EckncDUmtTm17LDfUCZeuRUeZtd7stuTE2J/mpxZ6eo6TceV
HOs++VEz+yDchpqQKB67JIDvxzYU7NCjABMf14ATV0jCYVLKB0LhG1rGBySlL3bp
Odj933xBBv/bvEtS6pYdY6lJqxOuvr1f2MmxnpwOtrjegBxFZpB7e2HdpgWTG5pA
UeAX3fvygLOImLKJ0Dg1tEWjWkjY7wGLMUVSEuwLZT7YYKaASB1fc9X0moUYXywr
rGBw5+nyFUGIJZGpvYsKSM2agiBZVOzn8650PTQW+u+5cT8jRUtIqzAEmdnEhsZS
ErLxHpHq/lUuTg+EkoqxAl+6hJG9ttjK2ganQ05wEQVAphClW7p0EjrgGPQ1XadI
3vJtydFx57f0dD+mGKxRvCnRt6PSRmBZpjEqT4uqRZb48AHFqNd27PCmV1BVD1uS
lXtAem608xleG02FLYabJyboq+/A55emLz0z8N7r5dT/URb7ohD/TDZx6/zQDarA
fsGkHV0AXfLjqfNoMtCVzpm9ny4cVhoPPlKRKcqCL988ZWgwvYP22rypX0UzWfEv
3J1FoAQSX7c/PPI9EnEU49uY3QLoxAlpMl1EGIwtur6YiiEDdIa9KRFMaP9f8KP7
xnKsEdiKAwpjOfzstM+TMFBOfpXsvNDnaYnnrO0okWp/TnrVhf1t+jbP47jiTE7V
4m455JfjBYF6kFh4w3wcMRQbzMBI69p7O+kM0hrw0g3nHWDSXZC4BJOWk88LzRJq
DL+Nb2DE0O1oNRSIw2HIq1p9BkONHv73v9mssZhCInPUxhC8ibZi7hB24BdglFQA
lQ/BeSJl5Oxb8Sk+aaF1C0RK4mUB4obsdpVs3nfo2eIPkP2IYMdI+Tkzbv8OF/Ua
VEFlRGMrf5MjsFM0I+t1xAu2BZUjg89tpGxENkbJuFI/FZwI2PuZ05uM1KqS2EE4
IgCj4L/yhhlxlFqNOdOcBUSlqtZUK3P81+mBNcoArfXwV5FDiWsPDTkJiHlOxR+X
lonUcdWdguXn3EfsyFMmrQx6C7v0Sl55v7/l7JgUYqaKrYTx9h3EZGHiRo3Q4mgh
DtEQIvkc1iWlu2ZLeFjaCj2hLzhzdS6drcEOBwJ8q6ZO4/+fB2RAUHxtls2f7ahP
yE9Kp4GcDJmakgnnmQRQlM3rkmEVdZv30wFnbAWUAU/r179+97dtzDpcWNitBTos
DzkM7ruGWitmbkSf/ZDNzlfugrMGmLOOWjwjbmUDdJNp692aMY5wfDIZl6Nh7aLI
PMpUSA44yBBfVAeIl8bXSABw1KRacR74Dg9qWfzrGs3P3OuSU4kbvGDD6AMUiqhD
dXXfejQLBAeLduw+brt+0h6BXTbty2g30MOyZWKnTH/niTaCW6kplvGDbNLxrpyn
Z3+/1HezKCcLOkkHZhXVez2Sr6XjpwDmL+/Am/Gd2k6zHMAPFqtdHcr2FgtbAEUN
wXPkrPeOvbi0dn751Im2JZTDMQ2DhYbp8HOkeR2I/x4RLUd7Qwrx+0U81gP20V0L
dq68zqvrUN8kccUnnicmAYLDQszrcJkstcMRcrqrYI9/nMrYXozBzxoODOr0oKRD
4FeTFdggzAVIVyeIUTr8wLmfx6vdeKE5I+UFwuv8KXXHjLSGYC1OxObqCu0GeIJL
tB3xHxN6elXxqLTiAmxvhPXGWfo9nBgkwW5I6zMHIcNLFQxa02NXHbt6HmKgUN71
xhisk4j5mXSrzwxZcKA4zS2G6hqJVXtMZU7ORgQYinoNZBotTlb2ibaEfgNRLhP/
XgT09jdW+wjCWyAGsOFUAj7PftgeDHm8GA6Oiq7pz9c24lnIe5S++Hdto++Hg8Ss
7ic+L4i74fw/6PXkd/vYBjbTbC2Q+KeDivFlJ5Immf5/P3VNGo+gPnDVg1qldZcn
Dbc0fFQve1MPFcdrtWazD0ChiYeBUMVynhH97TBNeTS4SW++H8QnXK3L1YcMVlml
/Ei3ywo07AIiaPQOHD7OZ1FVEmTBYcT3YlLtJxbCkiPNgNGg5l2WV+7RwSzFdVtA
8Bpmj+hbJFNUp2o1gdzYwq+JnyC8+EnTwpz8A76D1s2vph0ve41d2g7X/XXOQzOF
AaSPayggeEqAfGlHPY5316SvBOTEB1Xm98IKfU2QH3zU1gE9xcMf6oHLC00CK+8P
hcEDRME0VnXBlmCEyTo8BtSPdBhehY2hQV6hhBYO4rfDSBJRjGgAd1RmRpg7hYfY
qXtgGclpWCSk0tgI1fDgOG2bS76bE/HJ1rjCE/Q7o1/vOQJqeE2tqovDD2XO6dpk
QkXFbKwmfoPJGLvtQd0giVxgdT42TF7qJbPI+8ToETvKedreM5flomBtKU+IxceV
jSYri1RFo6AHzmaOTuOE3TIJKaGQe+jmBct9713OoWQaqngFDkaffD/FdPAeUUq1
V1ILhDiniDwxqvSctTtN0Cn8rWwARrwugY4V9wAcaBdpLpt8P3ONMsOCm8KWdRIO
tWuvenkENO5gRFMox8vaYMd9TxLOzEjCOM3ItMwrxRZcC+W8lVls8+TR0nlYRgYl
tQbtqXFLmdoGFO1RqEOoja+dY9CZoU0fsQwAf6iAqkHp/Zp6W3mOd8CFpEAov7wD
/PhYTZV/ADfG+xeRgkxe2JE/ufCmN0DO5ocqtN+LB7CXXe3wcRBfNDt2LTuqxOwN
+z9dgNGVzSqUrv9VL3hxAOgHCyKXRzTqTpQP1Ws6KkW8EDFRokzj0GrW7sWTGbAS
998C1zYbnG14JPx88CjLgcstpFymeSDrcsR+3PFp8OMZNnFI8Wwyz85C9euwYH/Y
uWBoX/JM/i/SeFmt9qZUfMvaVV44hg2h4ELN7nXngn9+RlNTBHPa7GmmVDrYcGUu
3f/8Byw4MOyKouviM6wdlwGKLzBF9i5ibGgflaDdh272A+C4EJCaQyb2UXIg1o4B
iq943exbZ6JnQhADR8gwL2A9k1qX3MJdZrSn+3SS4UnPMlenvk1PC6rxrCAxVWRC
6lUOckV0K/WY/SCFhYQgAvPA+JC0L4SQeveMkYEJdoOsOTtrkQy20XxlVM5t+kDv
u638Ebx7T8qDmZzagIOH8/vuUqM5LCFqOBrrLlT0JwgRGnX3uilsOkre0WlyBzn+
MMDZ96s9hXP6U7eOjfB6A7RWJkgTO0sgFtC4e/Zgs+dj182aboSlA96ZYWD1QnVw
n2JDHuK2FhZ+WdCpVJHKGsDyg3oi5OIidP7oviM+c0vkoaH/N9nJql8YWHya2ubz
DErudWnmZrcMB5AqwNhCQgTjzqfJPjROpwjczsBNfT8hGNVIBy6ttv4IKb6kjkNq
9HEyd0IqdmSqxwhLlrd8AHUhkGcyVkQ/F/2I0KiA2JvSZ/Iasw0PKcCPJBwAGvK2
jWYYvBvmImyf5vbc2DufsCrU2LsDBv5Vr6bphLEhGvDdjss4cOLm3Ed9ofPts4UC
0wa6uGgUsuiDfdy6sk1BmoGBEn4KxSJlyJZ0pisI0P29LoYl0Jy/1zAYQ6NOJFsb
5oOKFEyUTrvdXf77HwmdoGuyQTY1yfiyq7its9BKdzppSpryPB825EnZzRnVp9Fa
`pragma protect end_protected
