// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L1scF9W8Y6oZWcfPbUNsZqIs3L7oiS7JzN1STsffzWGvoYCHi5Ye/g45dVopxfC0
+A4voY2DfFIp2WrAAybCLqO/8J44+lD4I8pfLYlPl8wT5vtMj9Y2OPgQHItacfWy
pHBuTXN0xA5i2Rj6HdzvliBQvqtY7qvIAY/ehNWhML0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58768)
h9Z3Lcx1wIxIKGEkRg5mF6lFirRdIsJCocHtMBTaY61zxcK+tUZ40iEFuEIzAwg1
aglqqeoSbthlSxsx+nugEtCBu5XdMpidjoRAHHF07igPWkFPs2KpnofUfN16ZEl3
CxWcaXBBteJGq/69qFT0OxumywBhhAsKIP8KHZF4Bcz042uhYy0qWHI8UpHisZTM
8evH2ziIsL7EXbrMdPOym2WzgyvjoSH/Rvk8fEadhTnF33q5plD6Cddm8yflOlmA
3eSTzgn4gQnUomIK9uRTmEG3CZuR4r2iSz5xUQ1B+KFKdTHlqHgWzDg4UUiqmyxw
dLnLwRFRiqRrZelPEYyaiN4D9P+JkWs1QsMNv+1lUNg6EDH1xZuxe94fCg5kG2RA
q2gAUPiZviQRQIX5hyMd1xBwRspENN1fX3dTZAShc8AxtXC68samSMxTwZYSoYx5
SCtUktl8q5w5YHAAkN9n3G00tfrOtQyCEChA60Uqw+oXgQ+pISQM/pxJ59j73LVc
TjT1bSD1g+rER7J1vPfYjI1xi6C/wO3AOJSwryUIT+EV+VzzzJIx6O3MuQI7DERG
L99JR+7K7HIiTMATREdz2RcPwuy/Ou7mDStAX4AYIiiJcYggGOsz6F0EVcfVrTuU
2F7h9wKyoMFM5tc1ZyZTTDEP+LRKXy56OZJ3B0jrtZJBblE7PoSvjKyoXr5V3vhm
IvDB2G621T5UnlixXyZdAF/iBogXhX1sIFSd9i2+bYfjfEA2Moyr0u2kfMf9PpLG
J9urCtjBvx2nWWooQGO0VwXjYKlnWzySQbYz0rGdUDPvxB9hCb6FZi5AOAr4NPMA
ZnCnuYdy7ivbLBr3fDDDtDe84MvlMhuC3uvmQhuXGTrQu7y6WbLvn20K68WcZxTJ
SoEgnKJuSbYRd4/Y5/600ez52D0MWSJm3bEMgGO87gFH0zztyYYlsS9hwghDsShr
hJZIV4aVEQzGRPQdkGUgIZdWp/dsedUqXTElqPyMop3Kb/sJi4SwtHZPGY2aug1J
+RC5IiyHV/gQMoTOTzcwY+BSdmc76fLpnlcGbrOSBHcVuFiaNd75LPT8FfBd0kXF
g4n4BJw4mDV7i97BiKHf2hMWaAp3yGgfY7DfTSNNxYc6QOmoubhBktCB8Z2ePDKc
tsZ+befh+Kt7bGSb64WDn10+kRklzAiFYCn3eRtVrGSxCHgZElJJ6di4w4hLwHnj
KfgRNWOEheHopFtwSn5/fiBe8QshRVt/yyddulpqXBV5CSlTa/4KMu3smQTa1bjH
8ZquKdg1rTrhvDJjbIuSacCFqbhRmg/HWYF6tSY+PCwSXXZklgLZRpnt55xylHKs
xQR6OAfA9u68rEmE5REW1s3U/HXHxgr1RXpbafcrJ2LaAKifTvWWeyWGZReGhsan
aOJ8R8LcgxuBEWzIuDUwC8+pBUkeurUCzhvjs4RTvtYX/haInxMiQjaaFqNV+tM5
hpR5GjCUNvGOjJD5/Vl/OkHIUyPzUIcA1sw+dVbFoqbnECkumyuq2SLvmpIULQdz
AZBkBJJdygQx96DwsGslA3MFE2bL0pCgTXINkEBD5QDucd025yEDTV67uXGZ5iEa
7jMVYTThWnOajtmRz+WK475857aEE3o89/VxynrcpPN+i4CQXlYho3XyzEors+rC
Pf1O3rN9p25MHyGwqYxOJmgRrAo34W5kiPRfo+smWPcR0Xx1yZVG8dn39avpRsin
XSn5E8ANksAh42olK59mPjQ1e7wSUSiYoAgGQqs7+vu3uuETcnoXc13XgoSP0+zF
jjj61vQA+JL76Bb856FmfNiBFtNGNKUsVRCayfItUO3300f6HPgNnpVFmIy4KGjF
YXiKYU1u5sC9/TQ1Kw6Vs9vpVkxpNJu4UaUFYkftapQoLJSxAKG0hf5Zje+4FkOW
WwRP9pVuuw569lk5Hr9BK6fEYQkG7m5CLFN/6ISrGmLUxToUrU1PlQ9/Qx2Gd3a7
Jlezf9POw0qBaFitRopLQSanfXMKwR6tz4G/fDPsNa/bXZp3koKPZdIAyhX/B26y
noD1gQLTIfT+eBFLihAKs0x+IDQR+zc8XKwYmR2Y/Vy8uPa/jj3hjgYNvgRQRXD2
7uhVqa2gt/UFH4auknZXPLidmlt5O/fLrFw1HqI13JG57hh7VBFHz9jUhFoqR7IU
wZy48P+OPmEsZhqajSu1o7toz4h+miUXGsgQiDYp/l42b7lQsder8wqpNCBriNRE
R3oGxp2lBey4GCaCegiNiDWtyRRr2LS2jSfGWBTZVp8mkpR70yrUkqJykHwnOgTt
oWaIkKo9N2CzwJqKOpI5mPb8tYcUBPLKYBBqPWWAp+2WvPqYj2y9FgcBXWecSm5D
l67ZhlPozZZSp/nt/L4S6E0E12SwktNSVbLJipudcKdFXwpBENQvIX5pnS7sAF7m
RT8MoqnaIEkn7xLXaMqBRhIDT65HBIL3MOIYV4F03oen3FnbWmgJJiJc+ChrU/Oz
SrzRPCWfiMYmvOtLI9RZp+eqOd4BmjnnJNqfJB5togaQM+RQoXlmyVaR77g8IhIn
veaBQBzv/phxw0vRSv51l6fxBxbbHyhob1R4gfbyx1vOinJmbPWiM1jnt2Yci3PB
NCg4HpCo/7jkGTdT5Dughkqt5XZim6TSJFblx9/a5PxxGZPNpfr2YgrKs9pegjDj
r9C/tqaE+zydzsDviY9EUgz36sFFhg2SP0+K4D+XLCXOk7XLFjrINvm6LkTTFJzq
2sL7NeFf1SMYbFJTrja5/itEwzcxQSJBRNj+bFd07iT58+xqTE9bQnW4j625wAQy
wMVQnpk7BOxefSjjbVInfAJimO74dDrdET+xXY4SYHuOAcThJxDPawLzP4tqZjjg
JH8VbDYG78Nh8k3LKWr49ME9bmK6kX81HqYOYPuU3/ZixPMN7376w4NEeNc3oala
a87ovwD8bGJB6Ww0+U5cuS7dXtFc2S7IwtS1jJtI8u8ydO00GzGhyqalagVNKajb
kVPQN621CwQXlPOZuMkMefXZO18yHojIFd5dNU2rneskJPlBHEGe7huZQt6AjmYF
l/j4RcfK0bibEwBLgmpopbQmg9Bw2NY2fAC4rbfApuFuhjh0GivaSflIS5K6cxHL
JpE9vIyx5Pt994kHFswrcXBw0rwu6pDNX0OgWNiPBMC1QWk8EFyV9H4dsUSbPG6v
py8mr5M0bZlt4Moxhld/q4oPDVqQdEG5wvqSmexznzOE61BhiQEeteykrSGCROTe
VHb1xq+EWsmtovglPXqu+AW1Pw6J09al4gGUmrpTYlDfvGOJX2iOzWElc6IhV2Vp
pLlTNquk5yA7/4T9Ir6HDcNiYQeJZQp/xQcchpJRj8jNwF9LntJAvUJ3FplSixJi
onOLGPZP2GbkZz2zXMb4NE+IFUC8qi4cmZpnEUctXbQ0PLDV0+AW6OncHe7LrJGm
89kTPlf7IffqAs7o1lj3b83Jc8IXd9rjfkq1Q00SrysUBl7ujTtTeEty5qfCoATs
2MsntlLbriTkn2EbDVoPDkHiRc9h5bUN/9JkBlWri5JOiRH3+DLorE21vjO0tTOC
eP2tfHfLEKTLTw9V+EP0Jtl1mwIby3Nce90w/geezsiBBfu6Sb6jVOwUvabCZDrR
MW+zjR7LQQTzWO4gn3r1aZkvXgF2EMEoa9QT2hLbVhqlMTF06ieKXXVvDL1gfKHB
IoY9qZwW6oCtSPiCbRKO4i8xJpb1xSu9lcXqZxsHx9UH/yIQV43opTM1tvOJlKkz
iceO7EHc1JV8ar8aJ1xZnGIyQPIqt9dgW9G87+iS3/QqDM1iAJd+oodQKLDcugLm
Qvod2Tvwbn/uIuaoxYxex4N7MPjrG3n2zpwiW5jpT8hfyRe7lM7CEN1YHORIfK8K
/ZAlNh5lZMWdKR7mQBRV/fPFwVbybOV6PHztrX6BjH3QnfFIiFC3cB9ekdKLhRI4
Bp1hjVdnPvns2rLDQgKJSfH6PG8AUMXuY4ULjD6/2Fhpf/8iQr/PbwDIaLcVchP+
eBMFmKZq33pwPMKmbABV9I3HfG0XA0hlC8EnP34J8aJ71lbRDNNBx2i1jKs4UD9r
YuOfL4qE+6XqN8Bq1h12DOjOvnCSz2ZOMGD4q1Sxv/pI/rWpzCR4w6/w4IJ9ujnI
z4Jc1oGFoYLk/+s4TnBIF0dwmJQ+Sg/LbPlsQtGPU1ZQQ6/C3QDb6MLRYrgEd2uf
aCLiESOSNJYQpiQde26xN31OXZzKwv5M1t6vSJNJRIjZtgxBTmubLaOuhiQBKdsm
kCSZbDp10i7u2R4j8pwCWVuZ07aDIL6P9iCutzl6stVTIjpGp+mvx16x7Nh7sveA
nq+JhgmwC+hWgZg9RDeJrJBSHsM8nj+E3enA5mH+Yy1Exf/TpQcJWPGRJkN0Cpaf
6Huauk8mNmfhG2gopX2GpfCCRdhi0pGVDU0uDRyR4d4drd1BRzrofPOWfhBwgheL
sVG5D+YqgZHhOgyC+9yt/42UstnChNfPqFShjevRt9vhO/flJKnQkmMi0vVrGhTZ
yg9RhxM1hjkwN0FlTE+hCM4abhoDEHKeb8OSHJe+CcL58C9f0+fJcIA/DPXYzPKx
Blyms3zJSk42JtWurZrAtj5MvRIrdRUnq6trKyIALm0TGsNTT03tIZnEEhRoqqUQ
zoVP2XNfN82XpeJwujWbMhy6+cEf8SX+EMZA6v4wujxznrRVInZzEDJGG+RdYry1
UeGeRwC99Ldy/J8nhbWhntkaV+Rz3hKit96cq4UBBTeikcR8r3vS343rfEXjoxwt
dNLqSIbHTq8Y+OSrJH+f9Aw/qkhScRq0ZKDxltQfJqlxeagoinEQ6bzvWr81J1Ed
yaQQ2gc64GGDaOXzCnwOrZ4ZD8q/EYXYjK/QBcnyb1XEe2xEaYSiEFLJnXn0WjWX
PcC4Joe+VcOEaTXvqfnd01JSvMxaySAxxon4HukYnR7Zw2wZs58lMbBvGYiJT1ua
+YLsAlH5o6wwrFE1LUnJ144JWIJkgyMPu/0fvWbKlntt1zXrSJlbFyJ8R5iZOxGA
NsY0Qfjrby2ps1vXpDWYZoUz2YsFLE67j98AJKc+bbC0NYTY1KVsD7n3OFZQTIZB
sFIB3czv6zt+5Ph9kFwXGCARqpfFuTPxtcUWRwU5uHs89wMlYNIKeuPCYgR3Y/CI
SsM/c05RSoWifuneNMXqiolBFF+ydjAz5p6+O24vDDU7M/KQ6AEX5DHI5RJZ1qio
AlYM/XoFhvosdpn3D6q6c0jBw7+HckGpBmTxhJSLNWAmQfOf2Y3mZNgsn0/LMszI
OCZeMP0H8PRXkoeiRAW/VTH7v+2cATf0vj7mgW2A4WcH4TyxSVEUB4xH89sYe6U9
uiGow1lYrMFmgTUZWHYbJikdYXau+qFXxfXUI+/KXUFeZKWD9MC2fzM3NnhrzcM6
rO3/F6SFkad8JURyo7o4r7MJZyqycjRWgFdEx0kQ8JoT0ceaoqLCSMItnn4NlQyO
/f0upsOXLcx581cZpfSrb7lI1qco5IjzjDzMMxKGn9+iMctVStjyzHHBLRAWFXV0
PczY/TkR0ut9bJjmgni8Y7n8rohXbxf7aI8sJacK7vV1YpTWgCgOPYDgVgQr1/7/
0O+18gBOZd3hHGvtdPir8O2CnOFGfx1K2pY+8q2fAWcBrCs46FXSlwK2eNBxXwM2
oHaMASaazBwaD+pLWKK5tTwMgbhXt2edAl6PGjVdkn8UwJxfBd8nhrecRMGaemY9
ZeyQmTiHAxZbsdf14GlKev0oE1CRcSjYBaG3whEVWmP6I/p6vGehDxMy9YHVxDTx
GLtdVuY20yom1+jysnhE7sDqPTun0cwbdD87m1Qi4XYrclJ0uFQ+bcIJMMrD6P/D
UB2m7/k/M55jWpDxZdGXS22hqDnT0iW+Cp6kjMn7PdXSK5Tp/JtZHhqvsmkC9ecR
lh8CjNtU0uh8omlV+i+LOPppq7+BrUQBIn5QJM/YI75a9Yh+cW9NedzFwTA9GE8Z
QWJ2DmIgH9pWBKcr+HKt9PHK0bFqCF4y/2MUT7SP2N3NSxgWuXwM73T6cvep9Acq
OuYZA/LLM6WCafFpxJmmhZImrjSsxROJjgK5mQxWcP1Xns3hhhkn/JIYIbpJYVX+
xF3La6qVz8O2GuxfwOV8sSKwZW92hMA5p+Ve8qGndBD7DhjsjP0bA8Hu1G6BuPaB
QSa3RD2g0Cs6G1pKE+oGpVdfSMT5pqoSil3yjF7KJ9Mnt/c2ZPHxBxwG+JkV+pwk
LYPteqTSPYUCcqzhIq1lqzyWKxAYs/Z+q/UnUpUr358DyYyI3cq/eZZ0XBSTROgN
tsWIjObkHemcDjFDmtXZMmRT68/7VkwETNdQz6EuZmfoQoh0lCXBBMDlmNR2PmRz
XGhrkvYWY5BhT/tCG9UI4AB8tPDqa96vhbLUOxJQ+QOHayRYQmXYEfLJt3c/4SB4
6ZkQWV+NI3bytjAQHdkg/Dyg3Tj7EIAfyBySb6XiP7GXMWGLqajMwdFKAA+fbGBM
DdOTkNgrl2y/F5dpmhaixbnRgtqLmP903OavPPpFqXGVEQG8qlFu5aiAeadXegtD
SXoFsi9LhRu+Mdf3UxYrTAgkzVDFTqEOrUkxl52ntAf0PPZIGgDPzLFtVQPJcpun
BaEObc0pSqRQTIfZSIW+oABmH+dwpX66O8LcBfLY4PwsPvwJOZklRJT8nsgxutiY
67QONjvXic70RMvzp+wcct/2T64c54qWacqvBgODhAyKXEX2JmB9MEWSe6qtHoFP
T2iWb05ZbsR/LkQKFZGwBvg6J3ir2TKTkJ/lQegGuNnApLTdRB0YoxOXKLft6tsc
ip3oyIwoCDTcDShKMTIz2NobfxwC3sZdoYgqJiko7qghIeSlh3AOTU9xsnw67Vzv
Ho7q9GhwDK08nSxQXo7lIfh1cF39/ykJHFhtbcWpilsS5F0/vJZsxHXeZnp+gTO1
5ZlOwEUAUL4BZcfgu5XGA+kG/ezq8M0pLVGB5iVbOZGug4h4tpPxKefXZ6QKZVdX
RicpFJCf/nfOhke+iAFwqo7jtTIJz2SvNMcdwTY32QDEeYBbKZ66xBbSumkTUoSm
o8dgARXXszfOW+37VDNyxK9zYK3tBhCil8AkzU5Oowlk4qhKEF36X6hHyN8OuxA8
iITOa6Dhg4cuHHSwmvuDB3Psjex7B6ctrf+U0LhDIG98WbLzryLOdn+Jd1c/uTGX
Z159mMZQyOg2uIhRQ6qBZ4flWyfxR+aStEPtLFi8m5NcbnLIq55y4L5wpZ2+ogUN
uzuSKfoZMUh8KhRfA7f6j7tOWA1GmbgJ0oYR6DO7a63rCPof2yu/PLw1k0jCQVjS
d60bZsJpQe6qw0dRm7FQM9YTguOo69JUVR3jJsJBOVVSVguNaI2IqUy3Q0Dh/yK6
6oiulvOiGDzY2fJFG3OyWWH6uti/MTwTVJia6TqLupHgS26/SJx01JnVj2zhz5CA
Mm4MRtyEdxKx9YNg2cC+FqUt9xVZa5bl15CBHbRbbXRFdXULw+eHEIkCZjOnvvU3
ize30zZDfG4fmWhY/3IGrr7LiQN74GY32MkMxv5D7xqkkJXIF8tZkXsDFRg/t7gR
hfxb8N0O6U40ju2rrBOEIR+gmVnRu3oeotHnRFbCFQGQ0X5lXqmgxcr6Z+MxVroD
KnIxmKTlVpYtd1bON3hEjkcL3whoe4oV20LfdW1/an75zRbpgjn4zVqlydThc/Nz
1mrD9OjwZg5mSi47Z6rt1gDzv9GsdDME96qOOoj9uyFDti3qLFN5KgN7AjgerTX4
lWNMsY5pjovuEEYyXf2sAqtu9vwxiROH546T2eFWnvx7ULVOPePh1zw3pv+46S7m
gchLr+kr4qAWGanUKx4IC/2XOzafVwn0S/a7ZVpeVxvoCYBA6p4fxcZBVG8vIWT6
cJTNu91fK+acziVeL0gsZMDKL4ePP9FZZdp3tAtNp6LP9zI+R7f8d6yTkc4WsyoE
7EPmGrs8Tr6PXgiP5kHHrcjeo+666D/c7z3mn1wvad0+M2ClHEICHQRrEmsW5qX0
UwnH2X/c6mYkLQySvbT5npCrFiNA9q61jHARDFieMe+33en2lQHR9bwHiZJfzBQF
xXOGuzn7I012eg+vYbNVWYfsH8qrEWioh2iGlap3V79GyRT7Qa26JonlySQVEt12
sP7W/CVBrYwclwaut6iaazjXKAOHXNQf0MwJtRv6npGLtzVDJAnciGkqdcK4fOl9
LYe4aH+rOoNZar9HIwrDeC2m3SYGY1fvXEFtIhr/Nk8J1IpCYBhuMlzGaulHe+si
d0tNqmgs5n0kA72yt4/ZjEQaMrmVJhYdl4t8DUXmpvOS0kANkYUeEAbmLLpEnxFj
gU1OV8ENQXH+bgeFbvvf6DEgjU+LC3j7FLgWAI3/8RSndYSWUbh1Htpv8J1TasEl
PvGtsVT9r29i/1am1NVxxkroMLPRkahZxAASiCRq0jGjMVTo5t9WVeA7p0megkGq
MFjO9Qy0Gtcha934Ps+m8NXV2l/qbb89lerUYMGAJKIYe9tPSCFy74Z+W1mCLy+t
0On8MFKpE9/CPzN8jqNxfKXpvo+5MoFgpMr5S88NVPInUUk2DONrMTOroC4KjY/n
cQMgNIIQ5jvyxnKcLWSoXbxliPZX+WXELRRbDJ7ei889uwPIX7i4e224C2NAr9xN
WjoYoM72IBBRDLQd2IjRbaA6+xRuJT6po6tWMi0z57AdPfhrfczDugXtAQwP1QSf
QzjzaoKB58uKHil/dRAutLKD9NdweNnYit+HGAOx5qOV5MQFkuo6bUfhkHh4jMaB
kWyQ5d15Ok0y2zpErfEk8MXieue7d+Dzl/WIlOeVVO2+Z2HbX1fxF9WG2Uyfnb5h
J9esaOgJq2ULq+MSh9ljPkSBrsjaurBoVMLANxFLO6KguW+5R3Zyi7quu3NycpSN
ki0q2Bwg6lSrYE56opfo7xeT3d7srIjcQGWOBDWktR5RK9dJsWVPVtGbiH1kztjd
cH/PJWlAbI+lwTIC9If6ZUUfOV243QZIgDjRqMUAdOYBcqF44JOfCT/bxEW+ampH
BNoVY5/zT86dmj0IZ20d4az0SrA7yRMVeiaJNJNM72I+k4TCFFMrImy49INUSeGM
qU5VnWRWw6RINOaXKad6v344Tl5wj8rvvtLoHQmNYlFqW/1BkVwp98VhF0cHhZqy
+P6CWVKYOqIRflS6rMeRj8hZ6oVRGAIqH5pil8iurhmDt1qLWn5oOwe+/H5++A9x
dWa88GblN/wWnCJRgElcHubk+e6YqrIpivkxGzkGq9IegIukbYzX3WUQFonh670r
BbmJmcUiLqo/J46v3JbvQJeaomMlvk+wEJsUc9AiMVmkC4MhwOPV/PiLDk+400T/
ERwZg3T4FNo942qKe2XYSFqgjEkTP1OA56wKEQviRXmhhgT2H59ODImgesjqJEtq
/Eg4bO3BconqoXf7cfvrdE49RuWdm0bVl0UDWPtj0z/gnZbZspGW4gqI/haraod8
kK01zRZM2Y1EweaMqET1e+yAeJZfuW8ty6K+1FOIjqZDFZNKOsWEjJK5vBpEuHVr
C/cSsdi834NFPVqKzFjeMQfvbAVg3am/ThFjZyPJ0394HuyZovc0tl1urjfQ3fX/
HxryYjzGE83LeJYEAcZQ5aYpJWvP3V8UCQ2S98t7nYqF1fdjj9HXh2Mvq0ii2Q6x
xNKiXXtJhWVALCbimsUVedHyD8zRY/S6BHRZJJU3IQZILqT8AFDy21V1IjvJ2lZ9
yaZH6jxiL9O4ROOjAgwbqG0Hd3E0qD3fyamXpdT5ZfI56RLy5p2A0hmFw3MshLsg
no6x7z986NC0Pvaq0xgJzvkuLYEmtnDpEd2I3GnRAJH+vqEqYGl47HK9civ4D0mG
uh8OTOtvpdSZsiqOexQG7BpBUjEYbT8zyuzYaPuOlrFA2kM6z+Bxc/WPs/XauESy
wsIo9dkETQpzJkIdrEMtTtCDlFPMdj+oU6CgqoOGzlMF+XNMtu9ubfbPyBensMAY
yAfyBJdo7tULFglypHAP9B3Uz6GaK2f96DuuRqmvktCeNyRF7v+enViCPKTQEp6k
tjqyz4MHX8J9HYCWYY6f/9NvK8cnpf/DozOmpSJnLjOPJQgStkJU/+HAZJsf7BG8
JsrrGO3QYoi6XOGu0n3qqtiP0V9oeteZu8f0w6sp/m5ij/13e65Pf960dDShf3Lb
ksIJDhW8MJDZ3lrtX/wqJIf1sl6L3EbcDDdLULMWAGR0ZOxoCPLiAdT96LB39/0Z
patEYWZh7Fv/J3pD/y1NQ+kEGDK68yDmVt1v7/YD0711MezPMomuJ+rJcraI4UKD
gUtOCdJ8NmDcanp5rmLyESF2kEfvV48SFCpNL07D0tbjyDlcdsYJOBHcH7ggCy33
s0pyxCRHto+IXzgPKkeT8BIWNFTYnQ6wufFT1TKL4Qv446S00Z5L11oUgY9959/K
12FDEmXh9ONC8VfOQWRR+hQOSr5JN2KOLZGoJPz8ar+B6odf9LVZqlZ+PT5xahbv
/weWkV7DwhLa+fREE59u8RUIk4XwMv9reg8i3dCLh4QChkMz5LAYBGWg6Can3yas
F8oMABxZA6VLEHCHOI2w9KK8PsmrwRRzsizqW6HFB/KoV5VqgLnxFECVjuQ2dATz
NlO1vRSxf4qj35RWp5gpFN1j3Z6wY2iltUNG7cGLKOotE46YYCWAQ5PL0tzRs91u
fm/4TDfRj+rxnTf64Vh81rwGXngpsDO2+Rhq729HE1Vj5iLUmOXjs2HCB+4YbYbq
i2Ks75r94o4t/9aV59SO+NIhznT7iIkcH8zJEqfk16s9jsHIuPLgOrE/qbQ05ZNc
+MMgRxASytezR6hW6ZhsGcKZ/w4mUvMhn7Bf1uiza+t9cJS9g5aVPdKQQhof6YiP
Y/sY4N1N8q3ZVErzNR0F4z+Ub6j6TIJwQ9tGGBOChqndj0JpHAhTTM35fSvnJbee
B980AwO3OXZjyHSOnhsCm4ZdD7ZGzjKKGS7FFVJvXY0pnk9vKLNUBReekhleLPeD
kV1byzXyBU7e6yUCGkCr2s/vfyUmrqdPlvNurrOvwwdfOJtWz3rAGEmIAGP9boot
qcLFrBhddqzOG+/WWUuJPz+Ld9Ju95eit4pR040NPxKrQO1iDk41bf2hSNnHq/qn
qOStSNXmTkM6UW+11oNshQXV59pw2hsendAhm6krrm3yauYQwWt78e5NMX8by113
qoHvMoVOpDUXy4WIOQhklCaqNLizcvZo1yqGWALwQQgyB1I2DL1o6QS5Fmt7or4t
022mOaNMnME1J2xhFfTApJWgfaXsVRandg/Uh3TrZXkCdq+m00DeJYmewi3x53HI
IzJnTfP/R6y9jBywRmiIcwCM0Dh0yXuXEq03apNkqdUEvxC/zzYrJVAhf91zCgiO
J30UICFJgsFBEQ8HGom9ICw5VxT/UFDcCGV/QgjnOEdfUXObkPNIiuWw5iyQqdU/
EHW8ajL5TNR/OUqb3h8UFKiiiLNDipKKM3pWvJNz/EciTRXe8igAeMc5TuA1x+Mf
oHz36T1gPyO+6pu+bVH6j1gdBwZAUBH+G2bzJyUJLaWjG1ad3FwqN+GMEg9uXrNF
e33Hq9GC21k4cNHG8rm4rVrpWACcTtaPVOod/EJ5px33RSGPfFUTIQRBWNwWGj5C
GIa+r/nGho9eSF2Ds3YAvJyZBuck+2IN3T00c+Osj3VESjABCCjFYSdR7DyV7hTZ
ZLmmA3NarFjWmlsEsXidEKypKc0g2Phled+jpMRRwnfDEdGA/Py1Vsj+AQ/HYB/O
ZAVG+gVb/H31LtjHhl7T4i3TNUvgHRoInfI4dmy6VqT9SjUxY8gcRzjaQ1iloaYZ
UHKI5djZFX9p/7bhe6eaCVmlNst51ugGvRpr+ETMQGAXZrwG+JBZai+kO82rAQUH
KeLFuMtivjO9XTJYjqvftjaQdSTBpXnjwtgj1qPzgc1S8H5QGF7N4oCJnV4crBp8
+ICbx2Rr9dddJ6UbYOUW0veTNa1WxJ5buMj0448jFxk8Tb4/rHby8jX0Q2I+VjkK
dVGNsm4Vy/Z8nJmgwFPWaUAWSws//ACdD+pZlPvKYU3pEVnfHReS2vjuTZvO6Jc+
/XEplYwd3DvHFyzft+kCh2EoGNeLZx1oqAkSymhZDxFeVdI1i8tY78Fy2Pg1OBM/
8rtO5AtPRM1TUzuUBzyL+hgm3iJcRLT2Rt1BSvyqsmvpawrYOGf49oeGEEbl7XIt
baQf/quwg+Szg1inAfO87wWB9kX25DbIuUdhAJj5jbMuJfYkovDaU89yg42bBmaT
/le2yo9XYWIgFzhJ2VK7gOOHSrwArokZiCs4Y49AVgU4foso4TBqRcyFs/Kw0pv9
0G+OOAqa+6ifv0qqSETkp1cubt9hlnboqa/f5u62xEMG49HvjFERBOdfG1BUgRG/
YTLL8NZyKbmDab1SCOs27HdBp2M+Ed14M38CSGKLhRDgtZRAbiiF1t76yzdQx87B
PICYsEhQywmEK9fXmDJTGefflOZxz/jiEDEvUNi1kr12rzFFpg7EopcXlYSy8wdD
DXMeM9CuYwa2yCqcKF7zN0068pX6zjyrpoKoKypqiOVFp2Sfp27+fBqnxFlO7K1F
xkXlWZ0qcOTzp+r9Ti939eaql+QvyJOtHbvjr0kxnVeF2S2WZURGxswH7nWaVVjR
Z5E41wGqJ6NsdQ5SNbdq1uhN4guLKi6DDaGoSBGiDKOocHDCSTTOBfNi5eJkEmDA
jBgQAngeEiAfSrHiYGndJ6RkMZObQoVG2wfBCQVPUS/wnmZB0rhaAQlOiTvUQWO+
oHh9rpiRUYo0OaXk5gX2Fkk/HTF0IyWBExhrUx+f2Hb2hi9kgRyJDfddy8Mmkgy8
Df6SnoDcMIpizpdkqgFqmFMtInAgD13bUebS8GDxIwU+gi8koPsNLTWKy2EokiOi
FXCP4xy3Z99QHYui24GPMyMqtMXORkRg4XE+N9smNGpbIXfRzvKvlV3vLXWjgk0P
QgweuFmm/ibM3l9VXNn6SA2kZ4w6OuGiouC/DfgDrIvGGMfni16GH9WzKr8f91f6
k5pwsAk0HCzHgU+MbDkBSDFyI5SVjiVSb7iUhXklelnGaQz4FGQ1u9v8jUvUmcY2
/zAMbcst6CACMe3Bm95w9oLi3n4HoaYee+x4zagPlT5memKw+N6WDQ0oDzOOmAJx
7Vxfmt18UTs73KAQ4YTC+BQrSZXzyqC0kazPOocNqigtI+7SJkXvozRHFioc5One
wO9pJ5wELdWlr9gcHINnuGoE1UlzShTzFMGeFFeADFaqeoEjtwZP7Z5jD5QKZ9a8
/q4nAGwxF976u5ZYCai7MddB8/mbq50BlCq16OB1OMb9fLvAvX6z13lGLHqz0+3P
0zhOd3mHLX8EyWcVONkI+FJ+5XJDR1Px06kNWvCwNGPQpbr7lhOvVstoZ5CwqAFI
I81T2AtXH+F8FVxDvYDjwiYnzd5TrV9TI+mTHQnfhtOlFjqL/8BDdSVFyokDcM7o
gU6a/tpkBjj935W1WdWUG7r3qupepJ1Il3Eql17YHYXucvmYvSs+saWfa4w/sCHp
2AJPQSt2a7dGm9FwzXoxqKqMh8aMPDZFtTQUsef/eJndiU4Jmn9q1uXdzbEzRLfA
kyt7zk5poT8D5pjUQIDBgzXNJrJBhxhlfi3N/iHyJDYtEbXnOeXIIw+49h9+1nCt
maxgoZx+luH9PcRIy3c6bhG9dCMo6wOsCm/o8HaU803nT4OjCqUWMw+XfgTKFobL
pXa98LdqH7BOHWcGttaWC3btHH1jnQeJkO9U/TUjQlA8SgrC02hkZENi9ntJAkew
qJLK8gy7cn6qpL1HUqxle6vnEe99ULr64PuYdsEeYG8z9tZP0m2z+rLUy1eIt9Ke
XKc54v5PgvAIjLMYklfFh/8c04R7HLTH1Emq0kvgDQmPH3KojnIVuKKWNxW7OnEM
uaMLoYxk9DepEVuwMk1MCDcYnKc02RH4iuZsOWkdQqode5br8yph+kNwHeYB1MqY
kHZnDiTfuqAbBjlBA3725QP/BBblnYFCApMCDbxU/DQWd7vY4hBfhCifRGso73kt
HU4cOTgbRarj9J23gIUMMv+kofApHoSg/cqxUUQPcALxq5JTPRtyPM3xMi8F2Mw/
GSJh4HVXba8RIGwO54V7UF8yFP0xyatWmfKPGgeej/LmgcNj03cizyGIKnftJQBe
NUOPbcxil190/FzEKhDNmg9W6bNyGMPsdu1Wq0alg5YwHU6bMBXrA/HuLDYMPXaI
ShIBMUavuAHDZXdt+hQD2RfD4YFWZjFR8LH6ABdL4B8cbEeM5UFX4zkAD1/xsZck
OYpegFauXJBYLvXlvaMwlHsAUD8bbBxiDXOrhfL7YrW/uV5n8NJhPUAXZYEIbFG6
0Bp3Tb10SQfjC/K79AReB+OX8wFXpEMAktRQLoxZ1D29hmbkeaKcoHYwlGiKbgfE
QPBHAC1/IJjuJaEx1P4A9khKu+6OG34f+9mRErJ2tLVadMIrFEaKGksqmIXPoTgy
ZsDoRYGleGpEOSK5xagbykHO+4b9KgWORjOOOEM83mmtmSIyxQflbdXIzEDVVbjX
De0ii8Lmru1UCbBhLb7HtibJ8zvfTBl9NhGllyjzJoW/iU8YCfhN5nCA8frs5a/u
NUdw73H+GrCuB2xB0uGcktAaIG7IuzdjJfBYooEBTeIiGWDXyUUcwY1OJyIs5BzJ
r0IH7NnuyzjhzSjgv8/bHSQ++JGIoV4Ppiu0GNA2ZuY7RHc0URvCuAG0JUfKl4bI
3fLkYEhmn2zQyRbdHVvC0zXivCDcXMaq/t7JU7EaDcW+eIISYbNgsLwrjZfPDcfP
yGTQHu2MX+ois7j4nHkvqOmqdS7fOiweoVNRwg7FqYKsx7HvYsLK/Wl6pG6HvL2T
no4bPkYAp4gcKSwvzuaPMPckBoueouWGeMzvFopDSewtAGHyW/rmIndZLJPrQzNq
QPmRgZ85UD+HpQ/Tlwvir3AAkT/2bxPUNcUz3j2CGUe9qzgBjQ7WU10xgJOLjm/t
J50dT9TtHxGxilxPFP1NL+iI+BfcmNAAzf+vU7xwkuh28IzZlFuAXdeoLS5jnu9p
UzOAqqNHwQDYDriJlDGB58oRQ/q5/ASpuXFluum5otxoBu1Apkk1vULfBLtE7nBP
sMfQPTTLRPgrWnooBAZNLu6GzkHYqDjrM7rkrRXeGcty4Kf3Ac/NfblD5+B904rN
7L5OQ/wcj8luQOpr6aECffhniqj7oB2kX/oh+e+GjRx8IPo9coTZdaW7fd/UWgEq
prb6B6zb+8ui27aZ1kJ6OizeVMWr6W0hFI2ARvW0Of5gc/Cfr333eT2wbLySL/uJ
70BIJMBGTVK54MmopGt3JNwIOk2NHKjd64XDBcUX3DnDWaG36/v1N+n5j90uDgZf
+ZeQU/pXCO/w1oUTyBXuadRiYYizimbuEHanpZBdVG5gE0GxGtGkKvI2BGLNaU/o
wCByqmOGdjVeDrXZAtlA8kshfcH6xEy4qjbXrADhTGaYySZNCMlWZYPOKE3i3f2z
9UPPy1ymofHFhlJmNxh/VU9wWg37DeDzc8+SdcVlYHKbFOABWe+4MnETk9cw3ENt
X7DgEHK3gFhlxcvc2YWTMT47udWhJiPZDxOohYZw6hoQs0YJGkrs26v6venIlh2C
0EDiDVzZoxtiengY6gLOpb5EW2RupGyz9k6byZufywbOlfTKDeKqEDqBZRpDCvEG
vHFHt1FYNO7AVneTh3MpGiiF7m2rVZBwQju/oxc8+p6zfhlvG4nKhCsEMM5sDtGj
rPgAuS/6OQGPU6D2BXJ4InFqIpqrrf9enKf8Lrvy2jZzVlv1sfLZBYSRFexGWWD1
5DAGKcLAr2vAro9FOoNT/05y0KdorUNuQjjfJl/v0N3x0PvqN2HEfYavRqlu7EYJ
d9t/xnL3K9yk62YaBIDZs+vDEu5yVUHV+WS2OMOy3yeHfmjOOgPO2PQQjvac/cBt
MQohORPOEwW2z6wlquTtwiSwXVCM/atX+a4S+0HmIPCv5owCSkK46zG1kQnDaNYM
hFaJxqtI2R2buAKYpM44sY1PVIdOWDeTc0V6oROAN121meUPh0bDwAo/Nb5wfkjl
/y+owhAKfSubgJTRGKp0XilBpFruqECKBHjTVIMyIMEwskgDdlUzEVV82br6heP3
HvW7D40EaDWwC+oMHmqcVM8ciZTSDkTQots6bhOUZUl9s67he/CnHw/uV61Ajju8
cAnUTgDfPlhon39uADSsDtEd7Zpx1y+hY+QeSSvLmvz8/5BKJk6hTSEw++qK4mTJ
Ckl3TWAmGGvRz+rMv/fksYDUjOIKrswLG54Al8fMkAfea0dtqU9IhKWMV0ABf/+l
9nDJQGF+JKwSm737WUSGYkzqmT37q8Rh7tU283z1ZnWhDUKLCXYDdlLG8MGga2QM
0XIq3wKE7wo3pfd0H7fw1u5K9+aA3svk14Kzeu+QErujOe+pwEJM9JJS+qj0BZvq
xyMUZMM5nZ4GUofBHHXVw3wkLg8Np4Rty1CtFL7oeLFDU3LFpCI7NRaqSVIfIZvi
Ay6oxOyu3560a93YHzelwuAFrI0s8qcb/AbR8eAz1ikDd1xr+31rR1/FZvmpUj6J
rZZhs8SOTU3xSoGuAxhf8msqwR5J5cv7JosICL82QEpavUUcKNb82d+zUrRTeg1K
JsJ0vAmlVGfaqeA2+8a0pbzpbfeVgRWlw4e3c+KDmPNXZsKG4KV2Mx1WLu+a32DL
gU0VJjMqBXKJBo6sCIbYid5F6PYaVRQviymyE2rNTwCo77sT3aSUm0lRG26YETw6
Ir1IHJq+dMq13jkZ08DRnwTc8tOdSkZ59Ukuqm0NQIQUbds0t7TY7K1KIVyuqTF6
bKLxWA5JpMIdHTanTE/d5Oj9EMWTASZ2DUGcVTFQFII+8y+5SIg+s8+TC6ntrv5a
Ax4wtSKTdUzUZldji4MmK9pvrsQQY9E0aSS9k0gz3karU7DnlJdf1aLzqLJHV+ym
chWcpRHxpPHlXzBVR0LjH41ComJwfMD2Z7+FsvzbsH9HL79VWnKna5e0Yntcowq7
PTt0A5u6zf+RsrjSCkhVra39a0jFTYSnietp+3WmdiAOsW1yQwb6lfF/Bs8PuK7o
JODv6ptx4TeVG9yl5dCwlJDtSNyWGPBX/cow1lvP2Na9xqRuWJr1Jzn3B4I4NuAw
BcGiIWnqheRPypHp8PpQmuihmaG7ToIu4+4GvVerkSlmsUmhyp74A70J/db1EW0A
lj1hLzKF6emypqcsrctYJ/tLb/hfAemMLToMmDbY6w3bfDUOH9KiNHMhPv7CQA5R
Au16IeLc6wzpFGy2DuKWt0bntXjB6XqbwqY3oDU2BM4iOKWcAPjEs5TbIjmM8dXC
MCEb5as76t2d398G07Dh/jTnzoxzfiRYo4HT+bvAfigjvd6P7BijrZ41qJzlEMJ9
7tkIIRaCPt/bQS8F4jc5877I+hUDwKF3kMRtvw5peWGxZz7Vrq68YSiz1a8cx5mi
UTvXDVTJcI1QDik1Yxha/pE+7G4sW123OENkaiOznI7v5mEKwjs4aosOrTDCKyVE
rK/JkbITNBc3rqgDlFQ81iMrVIJt1P0Ja49jx5DSjFqr4/FUSyfTdUFvpaQe1Bl3
/hIretH9I3xz6U7wGVAdFIknYlZ61wmUQYBQ8mTqKO9c59DZD1s0kKemTt26tVRI
KlDIZjZhH/3VJoAMkBopk5HXTsWvEByE/O+IJDZr3fgsylyp4Xm+6LUsjWBWykKb
ejWWJytQHBRDXGG4XjQqq8uY5H9Kj1P5AqE4l21Iet+KpGhiF2D23vwqJlkFs6yS
sNlCW4OpABYaEfojEwx9vD23bMiqYmOsywQwf34L5wNQW0T0o5g71pTI10V0IBjC
cB7vbUzD+1pustNze3ny4+6o4A5zN+5lxsNYOViUaA2MqRz52DFefq8aSq9KXjCX
N03/VIAgsW8Q/ZzeGcAAml4gXXsuEZ1VB8eFKO0+oKGNUcf/ZZVMYK6yE3s+/2gS
0Q1xnzsrUMWQVxR2VzQFMzZfxY0TwrNlEYGPYy+Uey1GMs+bQsruZWnlF2JRexlQ
YMuHq0GAsfnNCQqFJ25HKQ8IM2ZgbN9AkuP056hTyJaEYf0sb+xwlBlQqS1WkBUP
/poNQKBylIg6jwnJsLqhrIXgbQceNarxOXUZRi4g4O6zu9zXI6bEn+PIDgHXOXPh
+JOxW5OrcQeaHkXdcJmxVnkrBRCkC9JklZBMI/IeXtBzVsWF/1dtyipYiosxlAAa
vk2pu5lmlFF+ynya7DWzVTJWhtogjjeXwCmAov7+PQ2QUjE0xU4U3hjSHv6O7B/b
f9CWlflsVUDiY0GpRFO5UF4fAaPTPUHZYs0uTYMz1Wbloe8EkSoGoKEzllA5AMYS
mZElZFAYuOWBXhT9JHW7j/6injGWZzWG0Sx+nhc4zNVwJflSAp8sRLLopyX4qCC8
DuyGp/ViKe8jEXHkwGgf2I6uhT6rxlt49WTEgCCOUthRcdT1gQL/wF8DGB44LYAz
x/k4F1ZmYKJOHHhgOD/bEKr7s7079CDl212WyEqixg1c7YRmC3gUpm6DTCRpoNU/
Uzrvy7ZJAiAylbvsP3TWJ513G3aYOcTlI6HU/azNOqyrxAg2y4IdGkkUBhKdQb6t
xdVzuuTnZZIKC4XBWn1RMbYwmYnHB1MfuL6t/0WuVw69rm23+Ll/SQwTMmcNlYtm
2sAmn1A32JWhiaQsR3+W+8y3I+pSV3mY64l3pY6bSa6iLKNV6+S42WGsX6Vk7LXu
OQ9kvghaZlKGyP6gxt7aaz89XRgEdYQ2GilNgDSkKFcQAaAoE/po2k9IeRDlfVu0
/t6s7NhtKBY4ed5sSjKWCpvHcYQY5c/ma3ZAP1+mbB7Hfut/z9WoNnzudqwo07/R
xlSUSTDuuX1w/k36Qy0CyYv0xVrHYylQ4fLukpUkbKlxY5H4yCD0ElFMig78kZbP
LAuWlf4h2QxQAALQuPltMhcmC7bI1fPX5ZlmV/61i4W29/WNZqdvQfIgyqX6P3+R
is12LFgEG/ZQFKJjjpswEAtB2VyKSCjPpHPtajhyVR43ikcHmSzNpneQpHjA4NFL
aNb5QgewqVmcJO+98UFQhNxJBoCtm4PoDsIIfNUyS27Gm3yzdr6DTGI4eHL0IUxs
Vgm2CSWx9y8+ijiRQ431g5RtIuEUJaWkP++qALQnTUdL7ilSeyadOA4hk+oRWGxW
UfsGd5vNxyVo9q3+5Rcg2cShEEUEXnvZaPtrthdwfT4Ph/5gG6rcmLjboD3iBD23
PICtrbikek9RDb/ge6NDod+un9u5SIj1np/I2c4ic2g0Mnvj/+GtlIzRe5xxx+cZ
axJhBw4po6iJC/7RztH5ORUl4nKIQvDgeC+TxO5JBT5TBDtFEgI43ZdR6VxUgBWZ
cT/2Jwcpc85JqQNERBqETJHzTMWJ88s6aO42M3i/6HfEjx5hU4+vdnfk79XEAxQ4
l8zDcJ8YPnTb1crqxrDA5gNXwqWM//rLUFSm+iGoFMbDYSGZycYADvOGqnQQL2BA
c69HJpRzQEUMUj4CjX+sZ+Xa+RMleUdU7xC+yBSUZKwcOPkwLrXe+kjFrvNOagB3
fZiVJ9uQAGd74XcS1rXZVDJqfk4efqaNUok7PLGSkTBuQniiO7fCBsvkb3b87TNL
HLFDG1eievTP1KSUnG7nCEA1LE4f8GT2djBn9QXH/9aULzzDGJ3Z+GdL8vwEJOz3
qq6olCTSQfHvIPp+fs87FytXTrrMr3X/0dudKqQRKh1EPhY/gM7iZOprBxnphep5
ORrtcMNhEVg9k80gBWlbBWbB6HgShYA8fVEl8XHlm62S4plWOl4XtbKo1qdCpbMk
NaIcwlujm8160p7XHx6dAJUrmtCZpMXuEDmG46uUJyeJGSF0fY5ZlGGfgRO4rcqE
LPyoIo9rx/trn5zZOtED6ALfCZVIkk5ED37WL5C741yjedfkgWKNd7DDMYgIz9ck
BRLq4CT8e7w6lQyw/7nDmCVzxqfSOkC+SgYIS2ueJthZYQeBlzFgD0yo0BkH8LQL
T1BIanqQAmmjRfV0Lue3iJTXM9kJ4uPvhNzKVRsvPAp5V1Ul0tJYH6QbiYlx1E15
IWNmF2Q4I6c8x0bakLtXW3B7Ov5GtT4a2NTuYjJZ18zw2E0CwMDzpl4VopGoEJY1
67x8f9cQnAhA12rs7vilW316AM7mscqATGnYdRN+WaSlMX9LgdbZtZqUpP/PDrmH
qGaSi1eOfSjfap5+JlNYUXhSkSSG8wE8HBxnwr2WQrhd4/ry7lrHGDAHsiWcV9Xm
9uBPHSe4Zn5MJnwtNy7eVy8T/2BUhLfYVrcwFerVxvN39i8FvnIKpr11dzY403co
ZE8LShd1Nzo6u/dcReiv5TVG7bBvWq7GGEgOWUFcHfQASTeV8ZYzkD8F+DLjELZ0
bVVdpX8CRnYAF8xpd3w6yip+AhTx9+kGyK4GhVQREikaLK9puOOonJ9X6BjxVxSt
VH4iroevnvXP9rqUBsf+LJiKqlkRV5faUHhAWGI7Ox3+B0lNQ0aYfUH9ej5zr8Ul
pb5npTyye9/B08Yz5oi6KArUBkcEQaTMU/0Y8JCcCg6c/3mJUj/ZWyQx8boZ1tw5
ChlGTsQ/uu/BhfSbj4s/dMdxti4GsDQpNhWdQA06aaZSwSvoWdPiAYq8gx4P1Twk
4v/yJRvvlHVajqkFCs2eOwS29JsLLhwg6vBi8RWGvyRfuku2MaiBMxfKfeIgtQ5m
vexXx5hcHfjYOllEYsDiMRQyYVcdupO6Xi6z1cIRcaKOgxBGalAkmJ3YGPgT7PZO
2DgeXAZCkMYZGXGAghAUpQTmNXQhwdx91oGJYdptD/ztDwkbpTuu9h9pvrnQIiS6
Vd89Vd5ongNf/LgfjZFlTDmEDSOnechegFL9toHgi8ODwnZtXiSQXJGW+Srtv9UK
2lBuSYLcHpLLItaGmPtQdjJ7KWG2CvSPzHs8Hcoqno6ZVh+ypFRlex0EfKlA+GOU
PTSV5NrEWev69YH92PtUIMoPZYsRbc3V/oCqmDpc1EZaYWOtoIwPx+RU7zb4yVxa
mHEdQnKSeyOhe9l8k7TLJRGdt1Pf82zNPAWWeSeMrqmMfe6iLFNqLt/ocQOg0JLc
9iemR2dD7JTH/lpHNXK60gMqofo0wzdDOIh4V34L66Fc1O77Sgsj9TanqzuoK9BS
MYZ4p/RQb7xifQ27U7oV6xnuJznsZ1z5bfYg4UFBzfrGJwef12Q9PyxKjF8lFazb
TY96IFUFRbZq4aX4CPAK5kpHkcomSeC4jB+BBeksfmr0f3ZD9TSWNmDLGhJF2p4j
OKgu4cAC5xr89xsGHlua+uX8+Da8oJhYcWGI+60NRMtncDCZGAS253jCG9m5z59R
SosQejzCjO+bFgXeWmH7KYVDwEv23SRmCgSoRSEHY/kRnZHId2176t2USsTtMd43
KiLQYyKeU/N01Eno3ioA+iEmXvP6jsThlgQscuAn/wActlCFQ8jNfLTTHq/CrEsu
/CKlx/TH++0PrL1Nlv3CiB9UsrBcqcJihaqaWpClMpqwSMBLH2D8vyc1I1wPIwOj
bwqICSOIHCbk6tDcoVjk0j4o8BMBxlxlr8fl7WR+yFd/GLfqlRpqq2z5P5agfrtv
qS8R9jDWN5X69b5+TXlDwsy0L1mqNTkcvNSvRSplaUN/HOcAXy8qiVADccmj0tks
p7RiS+Q34C11m+WdVehKQbiXeinHsDZxYBPlXQyzWniK9woihKq8jbIQs8Hjq2XA
xQFB98IVGduDL+PwN1PjZlPiA8EhROa1qvxKqoX17W62IbB9TTihC33fbuvF1gPA
wzUCIi1wCp2qn+Kl1poV5htwPiKvjTZK9kYAnIyKOPp3HaJNMJrVethspyfrCFP3
4gvgmeVs6zy9lbe4ixr/ZDGSzAf2L7JNPW9ZT46CfLQUlSq0YmvmBXydHzpspW1m
J9Zq6hH7Pfk7r7tSmrmUGAaNyWZ1LalKaK2EVgdbKCkq6vVx4yICTqisxLYY0Qlb
QoNT4NZqCBIESjel0hklp/YpVse8fpJPiWR1pNSMX7mZwv7/GL3oaq+bBuIaJsY8
CgEl3PoMCLuSpTD738HDt0U6htmGmpEMy3oHhnlF5O0Pg/INs5nei749fyoWBZeX
vPdZYnynLnv5BVULSxmmkm4GHR7N0WftSDXGeR0b82IsbCUGh2INuUk/mJURaaRf
9lgDodgO4B8CyTTrLj6MZvjM6nu9+Dxn2AyppRcL7IKtKDyMBDPKhA4HIsUhXhrX
yfNPrwE5QN8wzzVpgeHKs7O01oJvrNemF13RIJo3W12sZzawNn9G+QrqOUpstouH
mRHv2WS1NN5d2XZ+jAgYJ/q6uG1KjmGnjMazrFG7Yfs2uQj+BNblCc/F2hv7Bod/
fwR+PC/S7g/hxYrRQXYe1kgpPR6SfpJpCLzi5/pFUI/VjRGUVbGFNTLdlBlUy19p
OkW8OL0qvttbgxbusne4jpBJYm2EF7blssCLE79vosViHDjJe+pBwnFIwpJVYTHe
oFXyK6c4w+OVXyWX7dwAhePx+coIjEbvqTaCsvLJadnTxCKVU5mQVe5FRlffOSAg
pB50FpeQRagOj53qLxKZe1FU8q1jLj4s557AeqWGxe3vPWef7xc+qqmNPwui7/XE
4sLJS/RPzgEF79Ubm446MkxGCkRGP1RxyM/L2EAv0WgXTeP4ydt6gcM4qqBmtwTu
v4NScbzI/NDLxmEoEsnDiiT7hKFB1FqMRI1GAtj+vaFsoxbnswF20JF6osS4rjFc
wo+DQngcGaR5Bfrv6NnB6eIWCMDkhdmTwYREeMOsedzA/7+JBNgKo41ZnQXvkulN
ViUwGVHtB3/EpJZte3xWANfaXWGYnlw/fYzvqFx3Mm7HC4lyBWXuAnlyj8zhI/Nb
ipUXh5/XFZv+ZrXvX9o3fC6PB0dJAo5VbTnCM0BtHeftc/zpfGRGgReXlmqdaAxq
XlfMrIfPq7svF7jYjQN+RozFUqcS2s7y0Ao3TPn2oN4bpL8OWhJ8OGIY5yS1+wZ8
sEfHo9U/YEJ/4X5vzO6os+nQzePl3OBP1s5nyioL6spry18wI9sqBWYLPGxYwxk1
NMUWFlTvI9dSm1KtbsySlXV0Tkm8ArQ/GXCZ5nG9P7sVWA3O8o8cm4q2eST1d4GG
9zuyTv1iRBEkDj1bOw/6Pw81JckvACOkno1iobHkcSQeew4xT1mXZ1Xo7wrnK94o
+JzqSOaOkc0GErIKmSxHYoWOm8GXsIZbo3PFHBJ0oUaJOxxx3bCExZ49OnAqbMnT
nPmIiuZ1T6jFtCEewqchVtkj7jEr+IwBe97W0kGM9EuXPf8je0QmIRgL1MJ5QDyc
LrL8xU+9GWFETqhXE7dV8UGHer+FC3AsjZfW3hQvjHHPCCULSBhi+jdEvjp0LS9p
7BFI6dW7toCDnCpnMG8R140tEgtbTqAA/CS3wsk8x6yuFHEZwEP/Vwtxnk62LoAi
cBpMP3xLBD/FgCRvKHJTJlsrQgoNQhc9IohkaPM9d0ociseE5x5xDnUlodjJegfY
nSvK51kUfSavQyWhIIxd4vvLqW7hgJKLhzPr8+iC82EGiltjerGOABXzWYas9qI+
fGRPme1njT2qi6v1WHd8+LBF4hI7L0AYkfoHvffAsbuo2ti3fyFskbABmlSUI/D9
wamm5LWhlgCklbyw1MdSZR98ivvNXaR94OaPiJOyPYZmH6uP3ub4z0cJRXTQIdcl
2EzyqeOKowad8y7twnn8UuNoyN3XI1AT8gvmFDEvVGYhDMP1uIIG3+/4FbZSHy+p
JJhB811WZdepbvyJRHet0tMn/vQEO+7GChXOuIsn5FW8dmmlXk1B+Svl/TQWga4E
qCZWWFN/90jOZxoNEQtTth9GjqvGzL1OMy+KMv8iQnGAFffNsQk0RG19KfpzWp7V
YYBpfohEewYebpS5+goitxo/yXilm0AvLrzwUBfj3v2Grs3oNKtRh7avII25S/35
2jq/6CcXyZ93Qmn/7AbzF8G5X2hypJOs9vIelu6qSnWaN0A3GvWggf793npNuuNQ
QLwclV7POivsGFtkoWPcmpXeO7qbgbar24uBJMWp83u3m0ekUAFUVOhIn9SdJBMg
Zm1JI9pAojO5ANRkW/a0pndmLGM+m84enARLa4W/5iQvcoQTVUR+2HhUTl5Yqitq
XLb3GUvk7LhXnSo5+e9cIJVnwxhl2LSzy4dk9sWKQgAbTiLLM1CudbJuMw1eXPRQ
DJwOsvjeP0y3tyTtnmPO18JOhYyX4xd9yiEgA7Q7NE79AK7gRa/34lzQXuJQeWFt
ALJUbMCQnhgl1CsWehSwpyca3WIHvzVsY8moBNJhWbx/CXtZcrDG+XsZvuTmnPnm
7aCEHIS8X3bbP7LjaiGAr3uMyjguYs9pce0MvEmXnx3WHrczemMpR+YM6O78cjwV
zXLR42EtVA2mkbgY+jUb9v21Rz7vOPQRg4qV5q7DyNvNsuJdaYUDA3DfW1wqSW/g
RbeGHsZxztPebhuj7f3Bty/k1NZmOcGAO8nwnMgkRZkCMoItdL6gWAbJZZuGL6Gv
RV8KC8cZ9aLNYFo7/sSaXqnKGLMxzB4SFaDSGEF3ItGWOfimeFqfLpswHuyvVG2l
MVcra+h0eRwN7AJtxHvUbqErz41/RRMgc6yUjDqfgR1/Va0smbgAfBqgqrC04EQx
TRQpzD9ct6oNHND3hqlZxL8Pvsoy2XYRgeJzqcuHJQDDZANm+rCblZtu+siwmuqC
4F8QoK6EktiDEqTgEQ4bLFN5PeL3FWuEICbe11IAdwDiJjWp5YXsQuUv8IkPLVAQ
huqtmnBXB96Mo1UqO1lBh3mJgtT7nGl8/88ORvlqvFYECZ31wdZ1ugTbCF17fN2O
GDqig+ksLTCZHSMnJ6vmpa+e4oGYo4SigghRWsnNobAIUfi83jBqxWQm8kQ7UWTP
wWkhP/wUEmvQrKlSnc0sRgV6bHart0XBvs213HG272C1ZRQD9/4H1TrGoQkL7LtU
VQCv71f4f27zN4TdiZaFRYiYaeRJ7K2RWuh6pVN5ttRr0KZPtTC6WkmzZERRgx02
ANc/1I7pV7OxoJLU8YQ2XdRa8DIb2JmJ/thsGLLxg3S2CTc6Q5IryUJIgnzXX6jV
8w7gvo6BrG6hFk9hjTL6Wqi/UVOe83WzU3519IyesPIGN4dHpl9eHuAuds2ouszy
m/rxQax5fkzmfhUB8ym3lRQF113VE3sL29Pcu+5UcAZglMF+rfS3mYGo4uip4BQs
WvTSH3tKQ5ED9uOqhYUeEFoXu/GVqosnsWv4FCTnnDfWFtVBOJDhJFaYjO3BcRkC
3u+v8QuX8XrP76D/ETZgS2XL4Wvcjx4yAtqxg/3ArxJeUITpBtVycv45NGAk4HnD
jJHOUHol2r5R03NrnbASoZHtwdS5pEapvzQsOedssyVWjS8kL6513NOkHFzIKaJP
R5TynFBOplGXq/eq1KUmRMfwZIiJ4KgmrwwIYyuFhtOq2XP6WSn6qAZrlQZ45Avr
jSO2bcP4Gf2bS0L4jaWfV2JvZ9zxeVeG7p+D6jye+KQ42CC3YeG00oGFlhdW1Aq7
PcRrfrqP3r/ajwRG+3FIDMpe5ZVOC4e7kHdWuVD4P/y0SmIfVPaLOq1UapELi7up
5yT8P5s4u7BCSDjdmhUBI6xqltaQXHc6stBsaMyAzHhUNu08YLeW/6bTCyyXmsyw
0PSYHVei2OF0uPS1AwTJzasFqMGRA7K7E2mglqIw2dw5DnsB2sc8kxzU3o6MfZ1M
+RdAdLa5HGB70kbocpSTmCAtc75E/eGySdfPiSX61v1D3KbWUOxrVuBrLVAwMnaL
v+xeiHAXnda2nhu6XvUfDOjBeXEz1RjFiAmJVQNxzwZN6NTG700BzY0BFtZZjBvt
36Vo3dUnr/uB4SkTR2RiBHXTU6h1o6r7/orYiBuKsVYUgfjNZ7f/0GRmOacti1h3
UKt3xMcuXweCyUIZAxx2sObnB64rSJ4M4H6FuhIaz8m0qtHdDDn4IGzqwHRWnghy
03kD8J3UgLSD6CSMQwwQO6FHmfR1DRzIW6JFksL4G/FKOVi8u8R2FRVE7sFmWG4j
eF4pAu16MUSQ3IqSdErwuKIRTFjeID1iJGmTemXkUJPUoZWKOz6PBk2tJdQtNe5h
6EinKHk6KPKjv8YjSwZq4hqsF/GjlYQuFEa47t0bytLMtrhjHAizVPrWNFHodJbc
mXFxtzpVwLHw/6MFcDvtsqfR66YHfumn7jTo/1lIWKxg09cji7dCY/RMBTX5CyWo
bCMEmMfrGAcubry3gScmDmFZrC9CGI6Y20WwQ6DIggXfXt6X9bap6Gwi+vVbncp4
wKvPKkm/cdoKvHVbgC2EraFgBMOmJa5U0aIoPSmRiWW0gHWPpJiIflFsa+sMUQ9I
B/cDbHbfvrJw8P4EgkgzP3wYfEhMaP9vQ49W6W32FwMU6Ptt/K57urZDn0KTJQZI
BAAG/n8VWCfH3bHLRbRH9LZDww0RyrY0UkZhzjl4+Z1Zf0fv++fe49I/KVmjv1tj
K8Mv95yFbvqwJywroo2xlCOt0wbkqZImQGwc6PYoPOoaVL8tsrymwcJBprF45krf
8CmcdNHueMHo+QYVA0Iu1SniET/mRoiaB8q5f4/3QKGtUbFSeBPNEGxjl4hceX0D
U5Nvl0myPQwN3u/s4fgOQ/XtLjJmWPWYzxjMIpqPrPzWQZOJbgWeUo8QdOsrQKmA
E/aikLUZjAEdf2dfLU4it6N4cQGiTdc/lMoiuG9vKXAnVqyQvWTWt3JDZXcRGvfc
7oioDutfhggkSEtOgrwyNuKnlam9Q0rxmMECMMQXH0odY+akV7SHdoxwEGisKjVi
8Mz7/VPpzy7vjhzbP7JTXJ7LicXksGoCgpP8GdV7xoSsIVuLKd7CUCcUeHFq061e
cFJslHQjMmHt8PCbIwl/xSMr8H2fTV6U3Qm1aaswtwThJ4/uJQqfjgFbQc2wQnPQ
YxMe7sSxVf4LzQICHv7iPKLGQj39Pn+rsZmgvxamTUV5760JkcEkBYTkkb5xRiHz
mIUDJGBTkgcOl5l1St92PxdB4t9nXhzm+79SNQPM/pqtUh9xbDL1rXpkfwp/yhpG
FwRrQVBDpngOZ2Kx9aSJ5DvrljAgpq52mKWFYGnYI9hGSIVsgV/lwkrNn4nYMB7x
4cq/vsGbKxYLu2kaR21VmyS0Kp1SihznBWkCWIBsoU5U1pF4LI5Fov4Y7i9g7P1z
wwDZylOsLpoQ7f38lGMGf9da9Fow0SgcbTmf+FwPaP2ei5laJKn5oEf9gMG13dz/
D1vg/v5Xz4nWfAeUTLkmAPfPjGuuO0o8qOj73kWBu7q6kXDloL+T7+SGuDtEy+1h
pHcC4d2gE5pake74b9Q81I4VKWT1fUSv0XlyKMd4r2825h3rBoyK9Ukhv8dHNIq3
nibzdeCVIACimHRzDMhhx87pG3+xrHFvlTR7iO93zByRwcBGab4/YvdN5gMyFwKb
6zxP+u7ghB6t3jIOWvJP6EQavdxI7nk0y5k9qKYVmMjkXwqX8rBFU9BlxyM9/gmF
8y2wlZ0aGW5yaELoFTdmfmqZLGF1EenQ0it+34tkpLzUJIlEeGmNjwA8tUnIJChF
Z0PmBFc1mvgibGaR+TPMc3+/WzFX1wSASSriSI8i928U9j2awexJEl89pq2e/Ecx
kKR2fdY7mxuw8LROPh2mpcct+wr47OWfIKQ3dgBKxXLkvFUttF8xT7BOoMm3GacN
MQBVbXkVg50KiaQA89rzm1K2cDmtkhW/4EZP/rI6x8C9coiRZ4Y7eg7/0bpndEkQ
GW16oVivgIffWdiDgOj1GC9xZMYUXqsOws3Gxc8TqEpwaLET1IpqwK9bglusQ/f1
S0JDUrgiC5oHuiSYXHO/HY9+nLFBhmT3bxGMzvBRh5fz7nn+E8Qz2dq4DatDnMhQ
biBMdNxPfppd6HU51/JIWQNyWbOEnZ8iE+RIOOMahsKtl65/qXTgz0wSsKnROgEY
vHKxOXbmK3Y4KW0hODaKUz4kHkh/esRcGDsM7lpuykO23/8CJxxPwHh94ChzUsEp
Tc/Tbq9NakroPEdpa/qwd9Sx5n+cDhs4YnEeF6QaClOivqbgJf1GsTOcux+JzTJ5
8TbXslI7G2IAw/yRy3d8gdOQVlZXDwvmRXbIiPxyDDFWPKVDzMfuAS+ALyPNCuwU
050+ZZ1HPdPLYPK9L0nfBD+GCIJcxXQTCUBMAGHn+lsA8gKeaSFqErq6yg8TPwtm
4fXUSXx6XA2+2ivZwn80/0tMHm2olzEcdNn7a1oTeWBnIb1BwEh8y+a0eFi6PbNr
cQmBmULrLq8XuJUA3OdNEXVVlqEW+ublQUb8u8FNkMdk9RQJ3w9VECezmpKQuM/M
E8n5pyv0aA3pfg6Ztp8YAqwi5EfS97dcBIK0dSBNTsSXdK/JXQAlXMhtysJn3W6q
586LY6sE/GbovB0IDszt32Otln9XCn0klt59faXEQqFDE6r0OePsAFbnLtXGaje7
TAT751nC2lBnOM49m2wIBbDLb1Q2qxYj8s28CEyZ+QYN400n6kG34SSMNEJlsNJO
PcfhdmJWu7GzhGXDvYpIPK0q/cYuKcMCjdSOB1ot5u+pwCXmFzGgqwbqExihSn03
UhswoHstPamwudqYWZZuNx6nlO3V6RjMmV16SpQhhIjyNYEGJuwhmHE48DbRrlTe
P3t4b/ea/peKCSMVhAXJjQDyDdMQvZTrUxKtNi6sEIsUQIZIRCFmB7y+YZysF6G9
jZO3yTbL8YsEJ2ir2zcd45/f47+4R47YoTVqltsTpMUyiZCoZmhczLh5Nq/GOF9o
FN6vEkr1+VFlaXjtKypkSmzifgz2IzVfR4kOIc7GRYHZzzR6lHATuXp0gloJJ6TR
aWWv/9k0Xwdl8rJo18myLlfdud0T67DY8dAEKcbsFS+8+4u35XqMJivhEDO3tibI
LkaZ/zX83d9DyY9PdaQixSR19aPlw6qbGzDw3X5H4k9XWJsGjZAK8d/TyHMhPL4k
CATiDH/ruZZtLIMSi3SyAXGPS1Vlr/I2y5HOq4GQJGeSivssMGeA6ATPLtsqzoh7
w124wk+ktH8tFMEjrxtKiOnJg4J4u6FuDEpHBIh+f61/JG4VOPdBTHAL70bP6Y+B
+9PTovpcPuQJjk1ukxnA5fChiNWisvuSRbKpY8xAJdVpBW8qMz7WrZTNMNmwkS8F
9Wr54lTuvRljuxWIxdLztFCqxp/FcImFrb4XF6aY5TPrdTVvsQDHpusGMYY8Y9D/
oVNoSZUsNRmfWefhihFoMfzO6vcAGmjqJHi4PkmQZpNOATMTAaGnaSNracxYceJN
+E48NGYAVsdVWCG9VotRX3GnG8kssYK8Q9Sinh+RYIv3IBYSrixA3v576DkLYi/k
IWDO5CKgXiuvQvN33sYSUhLuatLywM4xCyfVIgIehDpcFy3deeIcAmiH46P/foQe
SQbmr6eBgw80jNmCB+P2zonAFaq9cSqr5MC3jbqqB0kB6fHU9kPO1pvw0KSsh0UQ
Iw2lqr1bCUC2yvkzzohPn+dhD3MsQOUzzbduda7m75UAK92x8ffhwF2RLEhNfwac
9zWO2grcmwDStm0voqTIgRzc5/NXiqLIGXACduK9fUTZdLG9MVehB4sb01A5iora
nTuH7eYf0kOL7BQpjQuRKQetVVaAZzYNGTm81s3hYiz9Z4tIVkmXJEl+hY4drsvv
9E0ZIDNm+lBGvUvexsv7MnxiV1FXSC52b5dleG5FaLH6dZjHHNx+R+2wWMpfBOAU
dm/NkdUR3knc3Pj0QsABKLmt1MvLbGRHhLMENno9X04VXdRrXf2u9kDAbdfRyskH
Bi+xZO5mU9Q58c0ipQ13Ze1mSltKlWrO4xIN4epLVzjVtDtzISnU0y7wMFugxTb/
CYu8WeRY4qB86l7Z3s9NYDt1qXKlRgn0JBaG9i+BRgIuZpbfjV6EUcIoGWpptjjY
zKTY8wQsJrxxpRao5P37eiLh0j/xihQsoyjNHyh90wq6jCIpHn0DnRW8/HvOmwoj
s1zWzBcRACAgsth8aYScU3SUmS7yj8kAzBE7iSb/cLYmNu3HPYDIbvxO5d5lIprB
k1zFTSnOa7Gx7hkhrzvMoIys2ZfunYztll5uqJUAaaRtBHec1ZrY0OGxNOnnTtHk
vm2fbdyYqlt++AwNPRzH3sAjVz3u3l+Z43WWZXDJiZCZM5mgThS7RbsoxZDaiCqg
TxM3obB6CP6AOa9iCnWe7hKLgBCFKLjNifzAtOIsh1SOMe2x7taVW8qN2dXD6SG/
r4a6jNAQetTu+uHdrnLpvLGxxmQLoFZYc44qYmhc0PN28wQUQDt1xj89zblrguYA
hfK2UFZ9UVbNO20WuHYcg0s4q9a6DiEK4x1fud80YK8LaOXFLcDhF+14BUWY31xN
/U8Q+8kd0z+7WaNph0sN8b8hu4Q+AIgSbyQH4Gkkim4j1Hz57uSfFBTUlqFTnVyc
PVH1cQTAP2vVU+NMhickuZLVYMKsD1J05w/2G0i6UpES4WIOXgilG50wXzIagncu
ZmAN6NyH0it9CN3Pq1TgFJxic2SxAM1Nld0i3YgLENaVF2AiVouqdMOFqJ2PqtWK
RlkCAMl5/0vx66nkH9QY+RVDt497rgOh3P9TAjCtyuMm76IP7c5kYOkopJQrzxVw
Q6ZHcrO1dzpBq+zeKzgOhlac0xRPbWLe80/sNSJ6RsiSmmou/8eRFplaUCLYtqf/
uUCbxUNa19WcDnKBLhqQc3hENoQ3XZgr5W7XfBDpktBSLibDlc9M6wUlI3tWe42u
IH005zRWMy4B6pv/7DhpJ1FrMkRjYPxeP4n6Tk/9HVW2PKF7akBvcd6pwamAL1AZ
UR1bM7fuTwwO7I5qs4GT7HVI8nbgusqPNs9v9UzB93/qpRd1uFKl245HSWZ4m9cv
St7ePgPjF1SnZFrgVTHU6m+eQxRmOEDnGIZEm6FM5BUYsWqaYA9x9O41LJSq4OEW
mlZljykcgv/9bdy4QDQuvv6Bn1pY9/jCSmF7MghgnhoaBFG0Ln/J2ZocN70LbPnI
N4WFysxgN+GFbEJ/AsxhfPni7jCLmIF72/9NdRvugf+mIlIFJ2v6zAHcWquA+bIW
0Ya47E/RgFEft8ac/r16qn8atJ1iPCF7lthhHgntUDYWj9RnJ2WonfsyqCL8+k21
18o2jxEuFEr2h2KcQvC0txv7/RHLz4wnlQ4JbIyCi8hbTCDhOz0sQDzaOkuB1OpP
20Rn2CJZQNJaxpmHa9sRR36FZ8vyvLtbGBTSKFNQWYqTYp/tTIoN1E0nrXszuOdO
v0Jy7KhuwhEFhuoPIZMq26awKaHMBeasdlH38Wecv3WmYeKQx7pN/S64KMASctuE
4Ge5ldeP3RTzkrHhp8s+z+HnrYAKg3rKKbHaPUfQZhtxKDth+j7tLth1iPR2paE0
nWGvDsrvYOpv+hiBRonJPnt99xG3sNaELHMKzugN7m3woJCIkFPMvFAh1GRQsW08
Hlv1EL11cPkIA3h5VT/727DKGAs0GNoPE4D7v/4oJa8inatACWNQgQit2sR3+yOe
JS1FfxDFm3BtvWRsiPKG2TwYDjdPtyd9aj2JaFt18z9hgJSUsSQKZdYNr6gSSUF8
QRU2Mzx9Z0jg0K+3PBAT1nJCQpkXGyw5yxYybvDLn3nPnTBh7WXSVpP+j2VR9Cf6
AZ2UwNIbTTRki2mhlOUyeOxGgb2Gxr4e5JpQLBPZ3SLFQr3w3+RNmJyv1ZuKK/39
9kNILbYr0Pb2lPqoqx/9jDNsi2p6eg0QTsTyVKuWrXRp4kwIW9lwQIkCt6G306JD
fdrrCtVelxGjrlFf7pvmpeLv0VXwGSgnPOdWHmjTlXBNayqp/R9UA3j7pxkirE9A
fnfmu51jEhWRu0Kmp/SviaTVJYkXFtvXog6FuSfME4IxvdiSdOv8GBw+HN/NQdq3
/+AbYCAxMPqXCjybbs6R8IhQuFn4KjXLB8GWgOzvy4O+sKM0OPCgDru0bBUB6s89
FzSzx06LfUi33pdDX9Z4dHxzQXpsN6qDIFl+CAJF0Zk5cIx6Laov3v32MTltyRoi
jMxqp7awN/5GF85MSEU2i2Txvv7oAu8EnOD4YhaxFqDIKBi8Y0FX8XLFoVyVU5aX
cVv+B5R7vCCWaTFGOT5ZrKHwtv/lQZySTiPh4lU8KdNp7+SbadgI2mvqww09QmAo
X9rv0X8Eln2nLaTviXv35mWZHi6h1FAg9pi67XoYh552rwOLho1lYAU1GluWrnAt
B1MXjZ9DJz3xs4VWGe/2A0hoVkCw5zYmWqH47SfYj4qLzj51Gg5Utfmmm0gTeQP7
Gkgw4In7jopLOLay2k9ItU01oBXWB35EewaiUdbwrtEvGdegIoILjrNWCFNoTFZX
WBHXdv+Hym8yNJLVlRDFDQjD1VOTqf+PcgsCebqvCSUGK2Z3xIeLdKnplkNuKPy+
UcTQoETn86toE1581u+1SANlcqebIMID2puO7RudT3Nvw6xd/lT/L4HAZCzFZJhV
beUtEsga+cF35cyE5gC5w+bggW8mhOUiPNODxWXASK5dweYE+cOlMuIunZW7Xx9R
k2H8KmF3FCBnyADxviCYaUBgA6m/OayyvtV1o/YsARphuANRLPs47p/cxpddzRFI
Iy1SWzyPxcDQjMOhtumfyOwEnihfoSFsyv5gYkz2FUDSuGyRPeWKJJ9njpDgeUez
9GqEnrEIQxJQOGC8sP7ryQvV9MYRDRmQyQC3cUwSrdOZkL6O0QntSHk93zV5blWp
zrwQPH7pMufpFU+omkfz1yrG/JE4wctyJJ4b1ujAYUpe4mHBKALznjF+YD3VS4Ro
7LD5QR9n7pOkQNEsponJ9t7Lb4bqUnHUwteE6C126j0ji9UaUGkLsyW9Xrw4ZDKj
ZTxxGVrUU3/3TsORKI3PIU47WDtrF40Kevfuhuc72X+t08RalXwywcZsTgc3Lp2z
7+CSxEoCsvBGqJzhWkqgEu+J0Uszvb6bmNjrw17B/PXET+/vYcUs/icLtR4GhN8T
hTzXe2kl1IouXlMkx1bnP9caY7t+NFQ7Q4fzuUQYW3QoknYI9lzJD1BXfqDjIsP4
0tb/1PRFGcfyuzlkifPHSGxSE6+TAhR+i1bCeDqZ0QLv69jFdb0bZcWDr7gv87dL
szwtC/v8skLE19TOH9xut9vchokzWT0djIPiY4BoDr8Z5dIADDPEhQ2k03vQzhUl
wNDuW5Sjn2+ExRB1gmRpIlOp/TbBNkEAB9waUS3WZLcCeqggG3QWkPLp8nxEzzTX
91Psjshntp91qQB5iq+9KLDCtvZ4LKApwq0FzGbk7KBXJbSlXk5B07nF9Xdgi+rp
m0NkURTDsWC9X7BUy6gNfd27BbfwzmyPqwmEZCZAyBo99qPELBWDIDiPz59O+TZo
j5p6xGgsGDR0Y8nwBL0p6xSSG1e/K5LuCetzkbpnoWe4tHxWhs8bQ4l7e6XYQUfX
cSVIWlP3Teu+so+uXtKy9oK5g5+Wox1DsZYg2GzH2rZlmQxDi/ye/nLsZAh3iHff
tHFi3SaVwA51ptLnkGZbbSm3kMU0vtBnnBYncqBii+03edDWkgJor2SWon5OFtSr
p/Tl+C4tqT+H9R90uhaOwFAYrHnMdh3h801A8h56b8l+eOKIHAmuqdjJt3s4iF6+
Lp2A58RWgZJDkPwsO8KEUG0rv4TPKcG7ivMr7LKV4Z3OzEDdpUbUWEtGsYCxrlAS
yDzwc1IfcFxb1dnoorNMNMGTVj8QzJobLaZQIyG4w84jodhgZt5sPAm6y1fMkFhO
OEdNxA2vY2j9enA0JzMqyvdYM2GmD5PADDLH/75KdsXYFwHo7/9BV+Y2vD1bGcpK
jPJS4x0bd5VeaZ9Q/lbxyc2ArimWNRf9Ns9X/zROv9vOOdZfjFTSZ7zYSXlRdMXi
40Idj2ZnhFUilkjPF3WN+xojPOQSDNMyGWrrSq4dtnv5Z+rAZ7B43q3h5MnnhvRC
vAw6c65dDZN/QXwNoeNXv7xdl0RtE9rzPMVuvjHOlYpR9Ag5VnFPA2SA62VOn6PE
c9uwgvoMitZ4Gvbe16fX48RZZAGfCIdF91RUlxjmQdMjBOUHHdVljGL3YdbT0Vcz
AN14o6ewHbYwUu52Dk96rsu5Iok80PPeEs4j/7n4irByj9BJzf/ZpGV3jWJeqxav
jcF7nFwRAxYRxVzcP6BfLZTVcUxdHxcqXmFffVms0O7h418anVgsw31CV6H2BSzc
OoAmMUHvfvpKgYCYc3rL85ZiOWcvKGnLOve2AKpkEQELXQ70LG2bO8ysmtcTSgQJ
g0GVJ+lpoCNC5XYlLz1nyiPWSrPCHtxzaeQ8AfFDrEJyh2Sd6pe/Fr5ZP6tBbHKG
ycsZMh4QvgAI5EG/ohRzDMJRM/J7FhczVwVhXhl9P8yz10Rl7z4azlGcMz2dVfbv
DpdZbvtnPGA9eMbPm30NTXQJYLwttI8w/KBUcaIDxoC6MZCK9uc8HRW6mSGUaYZ2
cHy1iTtqXzjjyF/ChSyrCRDDEDfkveDUPPL8u3+86LyLcjGmgq9qTp1YUv69+wBs
vqEzWMdPyJ11Ltc1n9BqVUmZG4jeYRwItoSI5ifM0utzsStLOXWhYu+PTI4hk/fh
RqqOu0VviX8XQNJAAWo+1G8aUesy0nmGcQLUD9z8MyOr4cld5oM8Of5y8V6JoBxP
T3So1/1tN5SaCSRxWWjQbOGAtzOhtA6w3FcB4zHD/AM5skSy484fCLriYowaxvAD
E+so7uV7ECkr7Z6aiDgHVEHKM7px+XqulAD67Qtls3TucjKLkZwpzZTk02W10yoc
PsmO0DYB23/E1VFvkB09LV9aHt7IBKgMifx/PsVPSCikA9JbWT11psqVtuChFxwh
qi8Zfj4Lyz4AWLkRvGfFiS6IWs0jOybSw4bzklvKyk6luntg4Gjh9GpYFuZ5+wUc
/rLC5mf8Ljf/9uks6fldOxbS1Wqb0fZrceK1GlEFugj/01gyyAaKgZCdPw7DJbqi
sZF+kj3pzWN3xLj+RKMD/Rm9I85Msx/DLGvdrPYdao0DNYKEaYcgzgLftuSGWiMe
bU5/CdyG9tc1szGTl69nqKcPp8nGmDBzDTWezJXzvK2H3Yskhnz+nuUoRmbUPhss
XEUCCsUbOH9eMXWoj2yI9GgpulfiN6Xe3qkgCYVeUn6CkNUoJhfJV++lQBf3vcee
aXr7e/D+9/G/+b47E3x7zesq1iuZA6y58fRtOBflITItBlf0rM4qSuLg+SrC74qZ
7ZELxgz098KGyVhqImsjuSnkpV6Fa+aTSawUIYkLmDuf0KUo8YXM/kk+Rl8dUvIE
MbQVFkl4zd8h6PVEHr9F9vJ5Xz/PBmOZLdUY0mSjVbZJbTtdDF+1wLVp9S6V41WP
fW8H6075PG6FfM4gEW7ZfpYoYQgQ/lV+E+522RPzQ6hoqGFIowA010cNC+fLwGyb
DfcoxHWVrx0XZ2RAYU1t7Kw7a1FGnH1Pjf8ijdtRCKZBolCanPpuaAtfI3GIFiHw
gQeYQs1WGpLufjUzWQzjHM4XhU3H+TWY4cXSzJkEfTo8ryYzOAdW9llIrIy+uicH
YUDuXDFyZG/E+drKWXnHc/AiW0fzeKNtfYeAI3DyrybdQnhMEeni2RIGTZlaDZhq
ywVReBGBqcBU1JR93/DXFVlnCMggEZjqn3OcA9OQiBwhyVVNYuP9H9iPWuHGVD62
6ZxQEuPEsGJLtbbTDsx36VQeJ+vqVjE0LoI9be88QDPZU9RBVWnUQfu7Ea837HIk
ejk1rVGy7XdKmGMdlMMWl/gFl8sCd5UBpe2ry4x6aBzk3bSXaUbD9Q7gMeWI561A
/pnRhiMhElfebLT+5T9U2OYzC79xOUvEixdijpz1fRtRajwmoQS+9mov5s6/Z73q
ytProS9wMDY4PlVO1TcxghyYoayt1oaWok0b+6q0Y+xTiNK8IbRIRfJFcFJCrCy2
Mu6RJmP7k7W4Hn3Eoo0KWvBdHu86GtK6lkT7QxRtpf5FCdrAPkbKYNjss3mUSzH+
S750QaYuyHM+dQddK3cgQK+qE6BvPFlAZkfAzmRC7BgwCAFpNp0TFgEcXy/bjI/i
y66nWPl9IRg7VuX9mFTYowpj5IUsCYXmNo0cPLkvB82E91s3viDIXAhVFWKzJsPy
/rgye6dKt6QiDfLi+qiGMs1Yca588pj4S2zDhaG00SPBzUPo6nwBN1+Kw+55f2T0
AYgMmboZeYxV9NdPULF4m3RWV/DSFSDsU5svN3VSwK4Lw+GJ3/OLndnRbYo8erTI
7YDjjQ97MUVqoUg+aa1UNqec7+PJcBbLxDTlfTjAcbGvphwGVyvXWGobw5MdcQDE
FSvbXkST2nq0y0APmwCtNix4sJui3uKZbNLM+xG2gIUdd5qxyakYQUmXC5uM7Pyd
llY8MJQ90OLlev2xLyYfnIII8Vm/WgCYul27sn9coQKGCc9LEwNt8o+UOqXGwMvJ
VfRNQ8iuNYTt9hwupSRkt3qa1dK+8nOHPgvRtFj7STQRO59qLseDElofGcE2Md/V
/Cft4Apl0yvcxxopAtdUX/y9IPvpeqSuaF3wpjx+CeFNKwBsSUy6FZht6trCtAVs
+0g2tJLt53aiUSlgw37/ZihA9/F4WMiZ1JE7BDKX7JR9xiXIyYYwzdXUXbhc4KW6
rTYX/0d7Z5vkVYzRHtopZn1ZxbHrUHoLiHarvBwIfl3ofhZgS1VoDvtp+i0MzfLT
QIFMzMTfnpSjvsC2hkHaTX6sWOsm9tab7xD3DEeprFXqbu3vX10FMWJ7mCBsdA8c
/bvfp2whkGfPrQXQEc6LMd5oOaUiutpU1iPdc+Qs6Ush3M1LOWSbx/yGrluFu/bE
s+JyxiBu92IKbzUb/g56C4gyzCBb20WzhyG+2Hh/GMyjzmbTO7oyrzkLoEINbTT5
fuW6KD/xtpSB3eytqBQtncxHxHNDK6t9omB0G6fGknOWNpOMXqV3YT5htZ5eUw5w
B+0O1PfvrYTPwD6ZHEadHW1AkNWeYVjzHD6cqdp4f+VtrGBghOY4gu+ObLF2Jq94
bFi2rxpPuorhJb+p6idF4zhU6FaqeaLq7UP4WECw+UPjv6jU+l4tArLHfbmLvqK/
tQH11fdLxresuvFvIu9dx3tJMMq6zB3309Q+iFlNpRkkJ9CQwti89iKnybA5SNuc
ZMSk6Vp9g5Wz12Qg7gehdFNIjXMmtbDzfHPpYYHAGJTQSif2WlgQhB3lxVijOISp
XqRBpr3PVLcocWryQ3110jGIbNhYdCN01L1xKlJ6mfQumBxdlWCSSnKxz9sW6znX
v6zpvmNWIo4kXG1tlc8pMBWCksQSaG4JBYfoAcMMVL/ayUY7M37YXK0daepOZrwb
rurFadkTk7usINW/2DUWBQmD4X9lOOjkJix4szrEv6z3NcGLZDSuXGf8IVs/sTXM
b7eWqe7W65n3DIZObyeNfZjkZOIR3IzKJ5lnx4mmurAyWN0Y0Tm77hrUoodYV3KJ
hXLDqjh9Ini8vw5yqvM4gjaCDQfSOVfNVdg8Ghjhsh5xywTQZaU7yiKd7RR5GTB9
W93PFiycMPIxot5Gbz3pgMqiK7stF7e/lsIGrctEKig5nwjEqdwHfzhCAasIdIKn
CpWiEF0jgjxj5CR8+EMNqJeBBMO/P3m/EDrL5SQTGAzu+w9RzmlxD9qwA9ETD0uP
3b1jEN6fg4BF+KxuHGuxzBjlo5FQJv7jXpmJqekVdsVdljJRoaO6Y8bt8SwxjkSd
sojgMWuNhNHNIycGARrerPw6IafAH4ic+w37h194usgxWmkxPjMGaZPA05fh6bDV
Oo+uqs36iHAop+2e+MyCR6WO5PTB7kbDzASAIlClzsCm6ec2wd9YRTcvU1k/veF9
7AiLKq5iCH4A/ZkvyjCtJrnltHLU4velnME/9pDRCpoiE35MbkQ/E4bUBQJu0WEj
Po4aEb+uqqefxbXzoW2jlgkoJfabijnS5qx5VWjysVRDYoiiKyTBsWBxu2eZc17r
V+Asm8lh6BK2M//kwnt4g5Y6+Ctv1mQHeuJwF5YKYm0uOBWps9lGxgOHPsHXXipa
Bvq+lFqdygoFvQkQZ1nXhRtJ2PQO/tH7xz88wfKYjc0CqHbY9VuBYn+Fus2ByFaF
9yQIP6p7peFRSDuYVpaXQkETQf21Y/mycj8TzgQflThUIIMXBhqHCzapbRLFsCpt
gwVsuw3rK1rJIdf434iNxgIjF36VbifwSnttAkRk+N8ZEcpDrAhMt8EoG83qv3dG
6kS8mM+sr//yloptNggsGdPw2YnZ1Cdl0lpXFBQJ0ZEhRZmD/W67/YAlcV1iBBgd
B/o1v6oAw+kh4jOSIQrUB0Ngh5aOWTkeN4fEe55YwlY8JXoOMxQ1pewxwq6KQOf+
BQ7sn8f+OSkrYinHvUcwUGaRshiLngz8Q6+vt0qrD87P18T9Uq0scamLQon/vYk2
+gSZgLyFp9roWAK4DOx5RZVCUGjipFKEKHNmp/uwB7ootAVT2lifBBZMNF74Bdm9
fcr3g5WXmo/5UCbW7di9g3S7Syz8iG58bJXAEw/EUDBupOQ87+7Duds9DhE0MGwt
WjhdO7svOSqjjUxXvjo0I33WxQLhNwG4jHhczioKhCoacIy/kHZiPJ5jDJYQQ1zo
O4sBcRieU52GT1NqKbupEC+Xmb/JeZmYgwWuekiZ3Gr3cpAw35f+fkl9Qh4cfbqS
aFJdqWhrk5wTcXk7XaGVJEI/M2XonuyuB9tmidFITKKyFzUo2CqgmKkpkb3x0WIV
RlfQ7TZTGSvsIVYgpJlfFrSLs2ma6YuVLz1zsfsL0sfI8dcT0vz63GEj5uYwtcM4
hXuTIGxHvXU/t83m87YJbs7MzSaUPUdN+VG40KQYY/sx7TpnZX9YsUjXI1FGjR3Q
37Pmh8dzfA0MVkYNHBRS9IjVsCeClxjsx3OxBZ0iUKmpLBammYcf+CgdWFvYk5SW
lk6ELXj8AS+hzN4uZ9xriW0KAlY3lDwvi00HJ7/edZ0fR6lhSeW8oXLjws8iGz/p
3kBAUANBHjvlCcT/XMdZfWjp0N4jqvHrKsQyPrzoO2LPIrJwB6x+DHIiEfc9djaz
GxD6N/fDuIHwOn8dkD7NJUMtdA2UyCbmSY+e4w32xsiXa+N5/7yF4ZKVDjuFOhmX
tXamodjrsK/vPpvsXS7lGLVmluj63x0kEy56NMTzTiD/HYcrOb39dEifYPmHksP+
+jgB7QhSLt4l2eqgBSyWwUIYxyccYGaC+E0AU5v9B5DWK7Irs3W5u/oG5VHL0G9x
EUQgPjdIxxJ3m9BmgphI5pViCH9Sqwz1gngqOpcn/Lp2N+fYCycCwkGMWEJCliuG
BbCv4ovQfhNEHv2cfNwY2Xrs2k2HsH3kaEpQA0gMXj3emNZVgGD8HCb4LNh12vEs
/vUSX8v8T53lEPyGN16LFrurGumy/ojICGALW7WVVPyQG/2cBngf/JTiz2w51y7w
hvC8fOCzmNi1xpHTkh9JHQINMNMAujz5Fx6qudyMtUwxGzSdEG1hrre1+oiRB41X
WNyg8CVmf2XXps8FDILBeJoeHFX57DQiBFmXXgS2+aJdDrGzZprPC22muJz1sIbx
IVCFo95+PGZHccT8Dcdvu7vXxpGtvzBigTz2pLaxwypZmUa9QG0C28uzWjRX07No
Nr983zJNwnxpcimBTb7zz1pu6rdrIBHl9ZJBARoKibObzja1AbEln5y+TnEwaoB5
PGKqBEEH8hz2I43bsHNvpHbiqoO2ukDohhCCeKRAzZ/oXCzUA03PP5Eya83cKosC
zqmE0zKDNV8keiXxORqPMfM/PgIPev0QEj20Z3P0NdQQkgooDHTaU7aC/udt1BLZ
gttdlb8dDO6OgvCoEHw4HV1tvxVyUGMyoC1OeN9AgE9AVaDpqjQfCCAAH0HrtX5j
CY6tsnbfABtyt7nqk6EQVb9UXlbCOxH16LwQ9U74+dUPSooWeABu1u95uDQbmVkn
iGUyD87S/JGdrB0336G1XkjiC7Yp4b/JnFVLmaJJkMVoIWBynX1sEprVNLhKwyJM
/jnFmHrE1SxMgO0kFaWCYxoVx/9hiyen+hyGLyBCBRUIjdP9SVLid11RWmlxcZaX
VOQuNoyzIKJ+xLKsIWrYWFfI9WqC3BV7UF4knGSVArines2rWP6n8oLinwgSaq7y
zlWXA7WAw+oDdfgROA5UNIjLCetIHI77C1W8KuReyaKXOcnYNcXlhGHfkx4xVYYX
jGZdsathWRJMaEWBqfcObh+F3ai5/Q0W193S1mhvwn72sFky/sixiOtH843PjGNF
yHk/WpqVAE/yWAN73VzulUPh19vAGLJA5A8mZ4oi6SFqooqftgTi6JzHrZDJmjKN
tTMpxvLT32wpgY9ulvBO5NnLYUjf5pM0CUbJyhfoRTOBPMONBU2e7iceKj58srtT
w6DoG39435lAAasgGHVJ82Qlvg470YQqNLUiF82ruMB/OPFJV+/je1rnXIDvEOBq
bpLYPeGYGUJCT9OCjn12TlsKPCUqjpiXWhAnE9R/BCADWSkGgdNq292rZ5zdG8WU
qHUkOcqk209hB1LUAwD5b8YQxLNdBBfyPzNeMgtjhcWQHfeG3Ap7K9QiRsI3LNK1
4EkYNfq72xhgpnnARIfIWwHU3QuN5fdBJAsBkvRTaH6zIkatUsYKl4Fe64zXDgjw
dIPdLOeCoMzLbSTF9rezf5FrZgLhowghpYNX19H7eGwsRd7xaBr7YB9CPH9/euBa
vBue18jbQUBfyDj711jZgu7MFHoUzmA7im2GrP7PCTOYkp8BiSu6TsH6i08pb8bk
Vi9qZYCmhZoiDi3Z9+FrxR8zRMyRXxtrR01PI8HlV6BPYHhZ8+U3SfAuwsFHKcrF
BjNWxa/cZJRN49ynTJ1/tqiOpzYlNpW8N2iBmy+/bs3mjWM+mwusyw1C5UBMSraM
u1q0CdzEwFesn6wnP6ociGDkUWgUyYfBo/GHzCgbMj9Oac6zy+oQ9zDeGiKQNcRS
fK4FQ4/hvjeKbuiP2tWKWu1bl9hD5QW6qlGyu2/KLuZJUTqJB1o7uy0gkmXsDfMx
R84t3TMkrnJwfyNT3k17QqmTYNntltAaZM4gX94dyBJG9Rhrj/WCiZ29zSqMwTA3
HHj9NVLM1GuZx/QAbFKeQ96fIHArK5SjJcxg+24CPnX/dr8yU9L1C0AwossAgCZi
TZfEIVg9B67FJraucH7DZeXm7ycUFveMwJ4d45oAdYzELI03LBlnTIb12dAM0McC
iY17J20YfGWU23gz9/n1aOSvMpG+Sxe4/UokPpwT+nRSj6HaJezg8xdP69hPPMn7
Klki9hcFEvNjSbYHA7djVAq4u/qpqIvvztNVXnd87uGGDTwIdDlOPK2vTZWZfUZA
VevjPHzubVKXCdtpzG+AjIoC9t3ty/iQYOtRtKes2tbKw4krq9lQcGxvHBG6m/uL
QoxW1wsHTXScyoC9IPnB4dUuDXeibAR66jr2VYClKZn29h8ggOEbVlRK1UpFA9JR
bKun3GakckCzWHPiM5ZO+M68nHVCn3J4p0vF7sfJo3o8K6Pezsyd2e0A+awx4FDJ
R0LIkt6I/S2ghf30G2xbUuXmt4dtlTtGdsGzd431Y0Gy1JF191hfI/TUSX++df7i
U25kcWYnUkr8Epbt1xA9Y0UG6c9I75gkxC/ICwFhf4SFLZSZqVKhK2Le8bhuRHUj
+M91+EjXqy7K9DgISu88IgCUBSgWWkDhWUOoiVN45SwUtyZeUVEcJl6w4Ljw4+0F
WGETtasaZC9Kx91jVX9yoFSCQiTNUKSNp5vJchqvYqqzKjbCE3PvuKtFms+i1Qyd
lMnFm76ZlCxpGbULLUNW5nY8acbsq7+CEiuP9PGAsaTCfs4qPOGxU6bYm4RYqPSS
dX5IyccoufmnUI78ft4DnzRnNbt/lORSfy+9wAfeUpFhcXrI3U+MRGFw5pWsWnQW
IJin6iKV4b6FYsLrpjMYCduiBiDMMp1WMTbJmkkaNaA/7uJYmctvQ5NTO8t+rpiE
FgHZ40cSn9qEXp/8xgChotAwBbO446c9iQDVlLP9lftTkb7MZ4lpTyfKuVx34gaO
CYUH06sB3HLLvRrzkrCqVibTx/7NwV1wYd4IjZxUBB2m1hogpKduVF9KaB3x6sOw
tpkMHRGi59+bA6o0FvoePziKA8qiDHu8XOGzZGpWRPJ8FbQ4YlH61ZC6sRGRTsvi
x3djpI1apTwwmD21DicdVWgCo9wS0NlhMjQ69n2GQtQw4+/mr22BegN8oHwf/NOo
a6fZx0npwnNLBM9J3UJpi4UAjN6j8Nw70Lsc0mImHekEIsTPyN6UnjzcwCQnri64
PavUmmQYJQUqZPJtFsUMM6bWTlpEYLAXXgLdoyplFiF3/KhJRAm4/bxNhI10BIkH
YHEGbYC2bJUBGIMbbpUCw2yue5Rhe088mWyIPnaERN4iU16ALKQfGKmPVa/lZeTC
IUTAXHa94u+xVudOE6eLOclai6kH4Kq452vlkfU6iOFxcTZxtJ2uwwktti1vDKzJ
qrIYzhbKgL5XcaUudUXj18qvEYMTW+4AuQkc6TkqijXclbvR8DVMho8eZZc29miM
8Jl0bSI72uKZ7ZOVga0/yhZdKCi7uGzbGLXMng7AUau2ZIIHwzLXJXn5WMalRFhl
uWHAD/gkXKUPpwAWOE37dGS0rjNBTccNaZpKZq5NRJAnSg52FJ/UasHsPq4/OYYR
qSvKTCV3fLM8gU+1X8XArrzZwvftnZzj8n99JVw71HPxpB2HgWweGhWH1zrEK3Ll
RDe/2Kqdm26hZMenYnMRvrj/QQEzoXOHMF0ouMMqiX2Ad3knOmnVyVqhpgmBaGJF
JuFYT4ir3yilvACcxyrIuRGq80+MugnRvuTVkHchYcpg2NN9aR907UXfD+TI9GIp
ULAACsP8nQk9LZX43HOvS2l7C5MJbBJ2lB+rKR1l5Dkl9VyxJLPu3mVZbTHmw1ZX
H0CVKh6sFuvj7vbclGOu0Xc/toSkxntg5KmXePF1jr8Dl8kEGuP52J+G5KQ5y/ya
4vGmnfyG0QzLF4KFx8pNzw3tRMZDRT3FujIKsVRt0VCBgmJX4Hy6gy07F4XHehH5
peSYbNdZn1ksFtL5J3mooCd2bgW9G+bQrLbZLwrnfdvsnKXgSLqph0xV6tg7sqAI
aw5Uug9E1ewozfkQOMJJ0mJ6pp8r/PnkpsWdnB9BB8lOWzmqlUVVZbl5890B3Per
1i6uismcr0lYa0mczw35+aTd/8m70TvG0Wp73LgnZuNu07iTNMHi0OQ9ySfflTll
rjIYtd+KtnKc55CiivJ0+cYx0qrZSucWXDHj1EHLqCRZRtgGJgiVq5gJVYOVdWEM
1bmWwiL/RvLldPCGNPjQnX6/4JYVg5jCK3pAXglRM0dQrZRFfL8FQwSDQbNZ2zNn
kBeNFV/sbRk8HrXm2d2epBBK1tYJh+eXCIllmwvDO/k/g4IlPLPhSl3kW+bzy/vT
MZgnoi4bcvWKqLM0RVlLsGijY8bXIjTwxxTdZX3haH9lEI/yt8drM785+NSkGxvY
ZnsElQZeEBwe7drENvAJN2I8dBBNwkvSAHkaQ7G1s+0u/k0zjl3iD08fe1xk/hqN
tBIHsiRRdHZjb0yAjlRTq7IL2Ic39A4XJ/MAy3ZoPiZ3kLFGlJIMk3iLXo7WNHfS
pUAsuffJIHzyUZoyvUDUGLbcwqXLaFkNVWS4AtsRWppCziEFVzX/cLKXgfEKAQfP
m35agEawoG59+sGW/OTEr/i98PSBkc5Oe7ZoTkf1gxK+CjJLu9h+KGHzCxZ+Q14q
+yB9sPIgye5qCEJipuAc7o2Ub3RfIWrCAcxv7I4VUSLHNWnR5JGbS30baT5bFBFx
k6ODiMKTO9LLZ8EAFuxDu4HOkAsGcagIUZ92Jtqypm8C5lH2Sqa3jILHwbLISfCe
5ORplPfshy+V5Pc980+B3HMWw0tPsi8/2crer+J3WcnCzPY9h3WM7mfLcB9hcprb
zV1gWR4JqUs1fFm/NZqDc8H/gLknswqjjgSv6bnn6KtyEWE6M75yytzvrGTw91vP
2Ck48UGdoqh9FiMo6JLxUUrLr/7w33bMCbBIwTBK+SiEMtk8UpWPZs0uEJDwyKt3
6GaO+7lQgbngw00KmLakhOSi1LjfEA03peJ5/nC1cQ/Oz52APb46MX2Gxd43ijMo
8b12QPb/BlHVZwrrBBudmL/mr5BcDV9fOkVEfJp3Iclmt5bTKBtgorqXGfEzz8iG
W0tJKvZTz0dKh0JGBMSCLgvUHsvL0OhUGeZCI29AVWId/jHYKexvxmAYwkrXd8ti
SuB8sLhAvEuaAFI4SCufQ83FN21gn7OObkg29Mhvgc9w5j7uhuemGxqkTzK4zyl4
775Oy/7uPKVetp10uskvlVRDcyyhLulLvcrYIyPMdVCuXkQ4GyTrYjtmrhhAkPl5
X4GwZST+gTRh5c5Oasr9R3O0T/2LiGG2as6gxUGq75d9caU+seITmpUkHba/t4uR
w0QpP/LWHgzdd8GickSDtVnh+6KtIX/6LLlFLutQQC0hcaZM+uCuzWs0B/hvBpnT
0G2x/zq6FiWtsoVjrLKvFa7myMN9O46IdHsCgli78GTCM++3WvsFQYjOnxGZRQ5l
SkkRgGgjxvK/sROvoIUSdIvBbUdPL6XppKy5YzXQUaF0DJQBbgdliklInVEFQrKl
Jw578sDUdkTOq5/xVurae9tm8DKljJ3blB0JNDwj37oGXPpl8Ku8McuVkDpE9cbw
jND1LrJNxMsnA/bu3jSbEeDd7H6AV6itJKodDT6Fmw1wjsF0i4Y1QpfUzAjZZV4O
P8u6ZggZfQ9BqeUb3YGnszHY49iN/NEjcv/ChBWzxQfXsQm+sdpD93HJkWWcQuPV
BxNTzNaN9qEfMhG8herS/iaydgbW6Pqv8AIvcbbOjAnxF6rj5e/O7zkHA+qS/ljp
tFi2kRsI+ocf/gLTc7smRHjPi5qJlgGyfFUyGXsKpKatG1bdfTdL0AAU+kp+nqGE
CINkoITdSqOcc4rzXxYd1fQ3Z+pq1Un3lDVZwtx+FdsjdeJsOlXj+hNkLff0VtLy
JAQKS2UspPjQPvjCXCRtmiEYwUJqDc6f5mNSUVh9LjEP68EEDiPPmPQ42qYpRYSX
ZCnBcYECNOIY9sOpDuBJg+3MatK56Gtk1YlYDTHy1Bo3Homyh8MJUkxxqDkkcI4q
hzvVA7fDmdUix67cdaGVZXvJBAoOMFD/YYmJUuKYX4Lrt5EPOTyxmgeTa6uVlqii
ctEY9n+AMsqUVJxx7TRURLNfZzk8o8Lozo6+zK2B9CHvDk1m1ADlpNNQumBbDpWn
h0yuqde5sMf73N1tzqCltZEg/CsaGqNIeV4/IQxcHUHPPCD6AjxxtM09y9GUfqmR
Gbo8rqe7PCZh1JWsD8D+JG+ALhMc0Z0qFlXTDG9diwz8sw8NPRfRz7oJhLiGlRpg
pd7UQLdmAcuQt8NRcr2AfHcRpBOkloUkSle9vTbHWHuxFbWTYNcRCcLGhy2smIi+
xuhLEs3rW8XDEwh/PZ57T8rLbhdsnT4xqHUQ5kK6DvuARXp1rT5P43fgJzQ+LB0T
AwjzaYmGssNhCA7j0pXS78fx9tXwNEOoaPOvUoC/ogBb2O3hpMJzmID2J/h9voRL
WSK5v8UaXgZonVuOQHcmv2+9P82r00DjOZhUbTCarZyF3FYwDsxD+i0Hesc+adkR
fN8M1aqxizgbScChLsS1DoGt+dZyRrM5PxrkvR7ng+2Zpr9W+5UG272IH6Lw/II0
WgvgDFzHNxR35CtFKb8XI2IJ0mPsY01WfcY8IJRkY59owdV+kjziSz8wdySjm1uZ
fVohMSZW52D2koDZdsrGwgHTlhAlZJ67IwyP11F7qrAzUIVNKMGrm1Rb6gYC3gSR
HTqprpXJK/WIou8cRxmfEhevqoDGI9nriL7fJexSMu/twCA8NCGeTj/eaXE7h3p9
dMSjnEOUaC/C5mGp2j3/EHpUTsjhiIpZwmA38Enkyacy7vpOovCcgIeIkPsP5Bod
QYggluYy4Ud/rfBda2IYhmOpuOxWcnRNPR0rdRQ4GwTfj7tKUI6rWNHJ1pvZoziX
CnFEyxkGQM37e1zNxonQHi81GPNNzL9Xlce1maohFylOKYzNKDszIt0SEOo6vSee
eXyEQkuhHyf1/H5MopUCGT4oTDL4Ie5HKi2ynuy5ygZex0sdx5qa3J2/6KFR/DVX
hHB/AV908s8IOqR01ix8hMpsK0/vejR3t/pbYpNQS0yl0WukAlyOhO85hWOFQhK/
utfyVEkXxF/ALAECpglxev0Hsa2LA/HLExF7Q2q9ilqfIwLWA7NSmIzIDXV/LjJ6
pqDsEHC9oR19MrprWBjFYOw+bBgiEbnYbHwV3ucF8MnSnahSBdmdQ4eABu8C6ecG
nes5KM49VmEM58XWhRnEdr5D+aOjdH29rg/LVzyAMSol1ZnOFXMmnkiNhvvaSgl6
Owxrp1cvkL22y2XJ8ZcDhqb5KGh1n/HO9KyWb0NvrkdWYaIN8UQ4UdjrkjOpGlAg
oqyXqjPXXaLYo6FP/Aq0ZjNuV7pndhikPyEf0yHTriqvllkhPNFMi84eZnyBX6Rb
aAOjPnweAIjeT59udRdhcBWtrCTRiOaeiUBsBZwa0x4iuBTMna0PhW+LJeEbldv0
YUI5Ww81z4qkFp1/kVr3DTaIHbBbLNg4HIKpz8XONpAMtYxGQtL/YkNvpLd4YfsI
w540/PJeCrQ+vPMEgDAbhliS8uWxB+1TDRIZjVX5H8rZtq9GhncQ2rI6Yo4yHMW8
2Ed+/+5RY53babcD8lVaY8WMEainVATllZssW9WFpYf4jJGsH0+CL3BX9CdgXuBY
5Ubz9vc09ItmHv32JaHxYKW7hke5NFyrRvZwuvl5LLxEit8bhQh4aXDShNN+O86z
8HnbB1ykp1ujWC/qhKmrClMuAsKX5Aa+2MlFuX/xGnI7jxD4vUHZklQoD+qQxzaj
IVyzZuNm1fxr2we/GBycuRxADrxyoGtam7FouFd3KUx/ouuSTiGLZOi0kyLm0cnp
yFOLFA6hndfrV7DMeEw8GRxkhQxFW2/GARi0957pKnl3lo/erNtnmAISAmilC5zP
1xTC0oQ5Wo3xnbGSROyDVKyFFMX8dTbW5QfTJd1yaaJROD+rrI2YJXWLmydGevuO
tkyjYhoRHiK2vYgmdDp9NxxRClqG7saDSBDSq0vDKHPG9ByWUQleTLzMpxZsTVkt
X6oN/FJUlGSIaz4K4pviXKd+h/PQZsl2l+14dWHEsXBpDjA6bQ5YGs4IfylG7Eia
8Y6Ln6Mfp0tX3fDpxY9Id2iAzBRtulxzDTzr1fgPpwRbaIZAkaTY8JZy3GQu4zlk
EdHnwePFSvIQl6h+QNdyAEgxtODniYC8HiHuxk9Crdu+6AOxtoK2IrHsqPVJiO8k
vF0ZrGnjlT0PYO+6scy0jYPU0ixITSKN8Q6jrNlkgaziVcckT7xsOz0RWYa3PySy
9bIiNNsXGcq3Lpu4bpKRrjYH6k9uuEYgpryve+63OWUgqh0Awgzp7K8AyGwMS96h
LDlZK13k+VapyGNHwV1ftSEkPMGZdALMca9uxFqLA5nOMHCkUfo7t7HEB3SQjRlx
2ZJcUJSfs3Nmyx+pcNtuy/WiNX9+yDJGc8xvacbmg6soypMwKwotp1HP3L2Y6AEh
U9vI8AeMJnn4Vs8wn8ZGuQHEXQC1qqyO7dUpw69CuIiWqzx+zNHNK02FaURSpqwq
aIwekKh7XeY3sDjAHqzO9nH4nFRRAyjy9eAIJHwvPkTvRBNQ5eRVczhT7gv1d9Yg
ZC00JXR40W0RZ9Jz1Q6EQpNNjvmCxMbJYVP/ZtmnkzclxKqq0dpldf4Z9p/0SBtH
dlN0EVcg154Xq/0Yee+HxhQHF/tCWmjP+yxklU8ObrbRJO1FY/lf7EjH2xL0fTgL
jiIPAf1XVG1ZObD6tC8nn5Wf13eoEdxuyXPirHjHBZkuu3CdQEHRYJoOia7Uvr9n
QLQoU3Zk1kIEuswhZXkgZnetbcJMobG3AUW7pqaBEcXFUjo6YQLUYyyH5T0oUCCo
kcoSZXjcNVYKnHBuGvPr6THZ9TDXv4NBzMWgBYctPmZMypdRj/nOXJHqEEuemfOx
h9iUrLtD2vQg3uukAqmElDDINEuUZul9q6+BQ3S1SZpY5/vupjq2b30CTc2MPznM
7cu2Di13qq3LfMm+SWxww2JH438Q8Sq9JO03otVp28Fhc8SnPWsxynW3xFA/6hlU
S3NKHaDkYwZiqRp+OkDIHyh2sleqEGvFjW/XdI/AKznvCwljND+If7+EDVK4A1p9
nKGpFBlEZcIqOPn0UvxKGYca6lDRYko/YM2swXuuOmnIndjumGQk+lZQMDWHTr2X
P9V2CIDaqpflhQTRgoZvEkqsGtEdwANpyJ1EbyfVfmwBWKlJ2FjlvsN3s3tWcpJY
nbaSMA5Hx7DJz5M+DXKsvZZorvCgLrNlvwfLOARMwOIyVG5nGBWtSWR68GHvNKmY
adEx+nXgGIX4QcTQBeuJH1GHwKzh89DNk7rtznoVgQJLJK/2ermxnLa6pb49iRgC
N4JWp2i0k+PEvPgrJg0S0hcoOydCs0m+M30i9P6zQPNKoJjUvUrp0VmgBhu9Xt98
2zHKlugYxG+Rb5vL4z89yMt+TVVhYvlNWLCQhK0MfjnbfjG8K+eH9w3tyrQ1aJmU
Noki/W1ms3NatVBJC7GrKpZvnmoi8d/vPiE4kKDxUmbUCCt0Is8cLJoBdH/lYU44
LTMArZC34atE+NYE9XgfN+of1CR5m8JKd/l77/vptD8jh6/R9d2q1XyEm/PXZ2DX
PSMEoVJb1oSa2+h3I1/xrLJc58dFCx9dxn9+xSqAt9e48TpYkOfbRTdrXZD0Vkmk
6O0sNCUmMtvRQQXeU3taYTB+vGpKDnwV0IY2DmIjfi0K4EN0gKILWALE4orfFq0S
xwV870PuZihf8kfjjUTG8jJaXxpk+yd5j6U+vA3S6xV63f6K9GP4pZZUgk2Z6+Q+
hocjyo6Mc+kfq+VJ20goBfAAXOj8kKNrbdmOJkCg85Tck1S9SrxcHWKTf3qfOLmo
+OmaVcwLNbfHsuzqfHCcGHZl5Tctm4DfoZPOV45BzgZ2WQetGuDx+Vb4u8JBkYZV
lLVTPW4fnZy6SOygTjcZ+lAGC4apjcwIl6Bd1LhXykS/M+LFIX+MDraOn5ANc/pk
otRjixXhV0p0KyK8ugIGxPlnlx1q2+aU+Gd8XJp+0n43ZtM0K85TVJkn02/DLNje
s4aNFmWtBlRC7Mgdn6p6i/BKD5iT4UqMvhnCYMOtQCUtb1VTaTepnTPZmfOiYVIU
yjIwIm7A7qU0D2D8ztBfgGJ4Vpef9hC9QZBz6R0xCqRNs3lH1MS7k5lediNwcpTD
CnIPBfWdmELTJD7MvwPn6cJmB/pwfBJRfYoGH8xzWp4WKcJC75XKfUkAX/F5yPp4
1TW+UoYS/ac9XWu8jF+gD+PEcL6JUsw7bSIq5Htn6qtjO7YdFlEdC/A6pTZf7On2
kQ/0VBmbs7OszlN0TFJSzktgMKnuuLHpSxy/mxff3n0mxuaLWJN1neC+z4x7Dc7R
BOu64dCtv0Ecvewe925DwLPH5TZ7P9eCxIKOvO387QTvfHEKVm9UZCHcTeY0I1Kr
DkbedFOG+LBTfOP+quScAQdwaLRXhN+CS1fDIgDrtotI7LBOG5ZpStT0KBoYOAGp
uwtJbfGvOXkMd9zs+VVx3RUf8GIQl22QuVA9hh+D5+q6Z1iX4MQXPO5n0yYq9y+T
z7FpAjjMPtQZY3JKn460KgfvHaMiPcvAfB4Lfb0Lc9b8ta6yEpUidPrg38SetaQj
SRatt10jLM9M57KdZnSrMMFCZEtEovgEWUllTu4nU8R/AgDfyYgY7ma+qbTW3Vke
O5OxTrMmdkHzVe3tv9rYcDdGdSMyFV+KRYHTYoW+4BCq0hMkArOzan6n2L7oyrzM
V6vtjVrluw+Zo271+YIiYiu8fU+M1M/O9Zd1j5PUaotfmx+TUhvS+3ryAXOfP0ZR
Sv60nmXNkzEOJKLDGxsCNWOHoaIcQYSc4TNQQmG4mSgWArVC+C8lgvnMi0cyu3GK
SF+hd5PChFOzHBWvNjKJCKD24JxWUhw5P1pE4WTgBXll1vS3Gvt2bncMRZwtK5Q1
9uidXxTk+usppfJJX9yWyMtotLD76SWljhRozY5dzmQ82HKtacdT2GwzFQwcdGfd
06w1QEW9e01ptQ2yFGce5gQtmPiUJx/9OtYIXNTjkfRcn1mBitAzqR1GgmIzVGqp
kSfPQfLMBnic9avnDXwqsw5etzMUZ8dmsWDoZJldGARvB5LfocMlej+zUAw0gqKV
2aaafccrtZIPp9xKKCjK8cjQ4jO+u5u+4OKSM/2LeCYBnLCbwDAwUM8cCk1Mr7Np
4SaquX9evKt5YCJAb+p7+9iNB87VD4PAicrWZNPSkyrq4E0eyWM/H1bJAYYhof0+
7L4JkZZZVL/O+Xn5uwIGkHtg99pdPKyBVignKP1ElYmjJXoKwooTRuew1yG9whTN
uYVQIcDoEezSkUxKcck9urcSMrR8XaCencDJD0YuSInLt3f7O6wuhqkmaTL0uzOQ
79yCviic8420TucP5mMGWxKVmBiEac65KmQRyTJ4kQX9sra9icp/LbVs642LjnNU
87ab79GRuYku0tDWBbwjjd/6EQhEu+2rkjH6y7+aZdvnW8wjuxch4psaD+MfQef2
uqCl74dcabwwPm4/L3DONxBMlYZKslMzkmEvHRnioDZGput2yaEDYm6kCWM2hVb3
anuzDxdQFaI0qyLEO2zMl8rSZxgo9ob+NNMprFlSQRnFe+sRKQkagSFsS9Ask9JZ
I3NL/pPBMFCS1rO7Uy/89j+NABFvFjkatjqBJE/GlOpNVlpbTWF7xZHWO5g+CC06
q4jf3DiJF90UMynCVX9InZVcB/cKKXtQd3O9ILnDeyAch0OeLms7nnx3hon55ECK
9BL0y7Z98qdL0TJEVctIi+yw6DguK+pqjAvFEAfrqKFcOARIYTlj7TxBf0o4HHR4
w6yLx0hlyGIWEDDhF9Su+9NwMi/N+X0XhUTjKeMN5cVyO/+H5qtkAw9aEpN0QBbD
myh+byDl8fx0k3m6Ga/Jl1w7bVgdhzVEWIP+NQbUBZ3a1ATK/gDwOpaC91AFoUiJ
V8o7S6/yQLCkTjbAA9ikQGdyD0QbtIBfmccV6/xLz9171CNFDa/9k6Xk9DVvggD1
hKLzx32Ury5vd2o1mBZp1tTJEK00do6fHh6KBqkcdH5WsHw2PSY5qTw5JZq67sJz
+vRCyzML42NKCc2a+lNDQZdIpSTIXv4hpTC9BRhpaP4EEPhfhVCd4sgRd5NleMXs
/nTXcQ5UGvdC0dX0wC+KM9zv1ruNFpdi+UYgusqttyFpDRbFImC5UYvNA9nxiFjb
49Yu1tEQRa5pjnd79dv1y5yrGLeIa+yJREPu/C9FxlmgNMFNWRDwZYjmjumKxNV3
1FQRRYp/SGxkuz528WDUEVMX/vtDvDrAQf9C9bg6C07oGCi0cxp7Y62DNKexuORF
6I1O9Phi36GFVCNlLMOti2OL5C8tRahFId6bn3ZCNXIwKsHlTfxXJDaKKUj4qLYS
HU3gIck9zl1oBlOZSscQDt9rX2o2im5bEq+uEdHI3H5M+vHwdA6UcMtCIkdsvgm5
RV8urVi6PqmA1EzYncF5NrvUK3QAahcUf3lvgR+0eeMsw7Xvtbb32c5dz9XjgCdg
ZD6YnJtpggCgk8Ns4XAeL/mLCmUpzOjFp/A3yIdNkNoz169CeFHy1/IYVkfGIV/j
DbA7E27aerNqE8hvxE9rYDWGAckETyICw7FVKJSSahjz3e9ruKvFUyZenizOC1p1
2k6x/Bu4wncH5fnB/CUKFyzfE7gDZ4jAB2fxoTIXLIhU8gyqVNz/PmsgBh+CSUFx
8iEly+I+1vRRsExHQquDkjq9ZiZIf9T4SGq8W0CSDhEKtCa5E2aCgOSl393iVgBh
f1Y3fRVGbw2EZnzcotkr/gu7FDFAv4Nj+NVZ+cycNAbZ/mQ66kgu5nvxTRr+0wHT
dDx+YW62s1qUTxoEH3z9vbh/KBs5IkhTc28YrVoApZD5cSw96NJqmKbo/EvSH73L
2u6oKzT9p48bpTOrKnkkGUADDGMwaBdK+7okhfSAzRL3ttuYIYhi1Bk/0fg8R5AH
onTa0L55FRgDRKbBEuPYfwAW+n577GjxbuRH0iGoG7WIMZQjHHRxrc+ZYSgj/h4+
pGTxcdKHCPxhYvSioLWsNWmIls4C10lROgzS8aHzxci0e85o/k6NUwtnSBHlA8AL
VfYAQZ0H3RE0Q9EN2r6zOcU5DoA0q1bAuUtE945I625GQPWnTfbeJ443kSfHI8sS
frbRkrOR+EZSSsDt1kBl/Ytjl+hZq+OeXEp7E+PMoN88gztCOgWR4AhziNsqAgbW
+opOZgYDNdb8Ty4Sy4lzfJo2KisyCclsQbBhLhOC0bVEATg2MTGtiJwa0qROanN/
sGvV2Q/A6uO8h20oamVS5+quGryFdpxBH3uo+5shpGkw8B4xvIealIpvzaxjdinc
dK0FPkuONRueYHJl0TVsjTzXAyyfvp7OXYa4dsZno/iyxp8RLsLHrzcEC8PdVo23
/jkzG5MKMy0USPszu26D6a6fO8TyIFcMNH/T6VaVZ2/fzWdwJQM4J0Wxhn5TN9Z7
K0PzpE8rVZolckLUCcRK536w93ExCbel7ULYaCEZ9skO7Xt9SZZE3r5gV6Hhty4I
CE3JAs+wrJ/mimUeTYvY982Cb4iCR7Zfa4ZsGPiCVYDDfwKg0Yk72xjat6+o5AX+
4M+4gXXarf9Dc9/vCNjICsfjhuv1P6nDgG2nsGsyEWcgeQRCgr1jZOgkJQE6ZlzI
TIAOdG4SfiWgSGUmEvj7YA/jGLNo7DeyF7ahqJRo+swAV4TKywFaHROrzArWbcuH
Xc65lMeyWo+Lqg7aMEj6weNZzhcyx5aeQ6LvZKa0FD8FnvjKvNpQvh2xrBaPg8fO
8V9co2ZTHP9AB5w1RvNYMegYBCU1qUfDSv9oRtvu/4EtYGbOhnze+owAH4L1aWGF
lbqKj92FBpU86V8gC8VKgCi1o/V7CoYLOo6K8B2xrYMW0bH4QmhSsFlDenojSZXv
a0uWCf1RggRrZcNz7WzTejhBVYYioLFC1Vgj638lyJDmBR59J1zkjwcu33TA+SGU
wsTIa3uEXdmkuVKZtn/crGyGE7E7PDTBmrXl9rMVuQl2HLk/h+g0+rGUIJkxMtFP
YysFsANagMJYz6hC8cE6eks39thhwPKamLvgpVpzmQR7CWX37auuyHulFeP9IQaY
9cKhT8dyqFWGcD+wWA3aYlGPIcGzIC9PKJ4AQBFE30/cIrY5iaubFFbOQ45wk9Fo
DhJ8HydpRJ2yTEDAzcv77aMeT2frst/hcFlJ49JXKIkDCn0sLVrrvh7Ji0xP2cC4
oTkM0LwampSTQz86FHqZPoJMWfgyNRDbYIeTK0PH+1A9hM6mxF9snzYB0rRxRRK+
HRscBGkruJaM+MbaVI/JGma63GrhL7ukAWeDNE+unWI9VWagjE1l3AXexGIjNCp8
1sPp4a7tLQ87SGRB8Y21ITy8pUm0eVje1mpJTKd08IZ7ExQYimtMmzti/8XmfFeg
Bjl35RXX5achobhlWJtHGG6uA2vJbGPgefk214M9KJ6oDSPNM+ZQIf2x6Dk+3KhX
BivryANhz1dMHGXjIgFUy5OUWh0PczN4aMbOEoQOC9pY3c8FVEQ/jtvO61qPb4SN
hLXtJxgxUs2kBZSqvwZwJt7aHOrTqXaEZXKIZuUQv0ipwopsH59s1+3wy+1HguwQ
kJFTUkYejO6j47qyHoDP96S0w/JJbhD294CtiCLmvUViP/oioP9fi+XlKqZ4vD0+
Hqogrb1+9xwAmy26UZErYHidbq9t9os76XJQLvS2TdDz2wlbkvGod1sOZZuObgB7
XyipBkOXgEclVUVsQkdBRES+G5ySSxcQoEo088nal72L/VQDwpLyqRv1TE+7IGPk
bogciT6v8V5zHTIOiJ8IgHIg0hoKhe3eHGf1iKGQ6ZibBJZ0umnv/c+HPf44huu9
zAI0ksbDVhneT6UEccT4TZ1TfnF+w0cA3H7cBM21QmUiToyBjDBekJqiUrEEC2FT
5h3um+W0UX6MPAnwXw2ASpi9AFLcodNnTPZ2N1CNgpuJoq6VXTDGqxDBeALkJl6n
qp6TPMdwbYywU2FWopUhXHIsf9JkTLNrAd2TKxr+u3gFHxFu1QqheyvbdYuzVnC5
eVEgNr1Nk2fIeTcNGvqI1JkkkW9prqXQCjVvHo/TP2nBbEwXzVgoBhvXt5D6tkMO
C7PJbwT9aH0w9/sWixNuZGRcd9loK9qx+VwTvCljsXqGL29evC637Ted5nvMH3Z3
mXGMZSA/GXkSMKg4ms4Y55Khgc7bncSLxvtKTmwaSwA1YZcoZqbtnIiyYTAXCJXc
f6lQpaAddPk2ah50WzVudcUFjq27xdlHJuLNrB0uO5ZpQb/Z7YKdWrRURa8IczLH
c1mF7fAVGSHjiPr2oPnn24oDxYk79z2xDIhUzgsFCFsZecf4PSUb7/qkxlQjyKxt
1yxqQ56MdIR5CgMrOceGnsdRZ2Lp/PgURgxitzVjwlzGbT/ZnjTIfkqyLVJZ3uuq
zmmoDkHCUzPnODDxL5Mpn740GnfA63XAD5GN2P16OFwNKOf610bKKAwBztJ01l2K
NlXotiLi4HVQSm/28M803cEOmbIXp++KxNw6zCsC0qPXsRBU0ZU1Y1ldp4fZ005p
7wnFcQWAGrUBQ4PVaIRbLXbRVRR0NLNakAqav9fQ+nRT39ZXN0tmZn2lpJezS1Ld
zUS7UYlanau5tH2eu/JLd7nV1CLMeXDAnerkmAwItS0s8HTOD9vIPbZM9vmhyhzD
ihF2f/F5lS700UUjylEQzBoSzvmeYnB4RRTRRLJ8FN/xQKDjeBKHJPncLeg4Q8jt
Oq6VVHFUjA2jk5VPGEYG56zKyqwQZ8v4nDD2Gp5HyqrucyxtDedI+Kuq2V3NIeGA
BLobUypLrdsArZkbPtlMRYIpIMhDGc5Uf2fp6IL0i+CcQE/NA/8xP03TPEw18a1L
DIu3eVBKYV3J50ZjFwcMK1hLaUVlpImMyRmsoM0oR4TE6AQtithdlHpcFj0liTH5
Hgz94dMmENmTJS8v/B/bNy8kPkhQ3NfdDj5lfESVMYtwxmz8m90Km8bGyyEW72ZY
hs0YHCVXYbSkg0ul0MWEb/GbGC4H2ZUnHmGTvZx5JSvtPjLsUp2EbbLW23PviVot
jZDsRzLNE8m+EpABGg3O/cZk5zisqWy77+O0tV+znl+ti0Ftopt9HeZfAPeGPxPR
34htEEaJPKb9ivFQhF3Y+Rg9QXUjMeoPaiwIkt39Np3AfREk4cefMUZ2ALFBJbSh
CpCGWQkUnjRIvj8L03MvX6Wjmeich+sm/SSYzPksMeXptFDGtrLq20McHi+lHxWx
9RYZGx6RMZ7QG4bKZtf8Tt0X+U7T+y6WEtkwI3/iVdS0zP5ripl7U8WNCB7uRjb1
HO9tmcaB+apHoWRY83JYr6rBBTDpEuUmRasC6aPgteNm8N4O1GoFYBlJUZ2FECZn
pQUiaegRN2iAefF3u+fd0xbC1tvuK9qPw11kAplvLXJY5KacMlB32MBMIxe1qUlk
Ov1vcQadiyFzunwKq86lLKkJApuh2aXShPuSmeuYoV/PTxB4c+CHiJF2c+R2t/6h
QQpLovaw5SxO2m7N9+mYWPvPp655wqsffGnT8oyip3Ksu7Fs7N4TTProVu789fBo
d2HMFJdzltpDDHaIuy1rEWrCiSpsZsM+C1FZJL5s+s2VjKsy5F4gO/68wNuy/rfp
eaWP0iJgx/GCyWZteuLyG15HvoVhHbB10q1AZl3jgwvQZ7CazyvMIb0yNYzWMf6P
tcNiZA4KUeWgYj84G6v/v4UcIuBhTHfL3v4zAgAgVcWiVUfxPKMWd+ZxFRDS9Sr7
Oyou/LC8kWJdE5H6wE7b5/9ceemqAb7BCxw+FMzOT/4UQrcwSCAkr3VvNYNbDfay
aWQ5MQs0fvkjyU+pAMAoB9cAEAuRfUqg0WIA8UNPrCKHtwEn3T8aNtGVZCgk/rty
tj1DbIPGfzd5+fmEyQyL97/cMmf3x0ABDUuY+827simi0ZyNiDI9tWFcMKGFX1Tm
uuKuKiSITv/cMOSLJYyyfOC0/VNh1DncAc8xD9qdkjPIMIxFBogWYJ7ux2I6GjPZ
4YXqHCjY5boENeKGjc8dkgCeyXk7UTDo0M0SgdZvKhK9EPpENa48b7Bkbe1QEvBo
ZD/kM/HcZ+I2+ANnIFR3IkHbnXyceSCstI9BDWod2CfmiF3MT259zXOsmV07ytn0
dfJPymSIL9EIqHtOEEFR7hbShZGdioXTCKtjg0WMw2AzXUCrQfgS6770w6ZpjLJr
b7/CydnrcDLrYrhrd/uJCm2vHoXK/Vo2BVo/AlZbAZ0a0DKW9bT0nwHAd8Ha3XqG
B3fb4mHJXzLY5F/v2ih0YhycM5XEP1HfrS7oRDSDRNB+FKdw9+AhY1ZJ6zMctewt
88FGAbRX4Sb4JzQxo5wwONIaw9LftEmDB4AJ0tWDongrHlIjpd3AJ2xlEDygL9U2
caLU04yhCQnSR4I7hwOoR7Yq9AEKhH4Ehli046p78Pbkp+b+AA0Zir2bb4WpiEAc
zvoQFZaiaTfL71vDgvrpTPOOpSqq5ezXC8nqxZRuDlhk6RKS3GLunYG0orXaALTc
cpXjjoB08L0VCyOCF9N2L6ZRQUotQtSOgDSUQce0eiXLdQfODrGUo8r9RQ7VQurk
3xs0nAucyKqWXMO0ocYr89DtwOOqXU/6CvLAf+BZ0nUqJ9mC1Qt4NGv61bITPOBX
6ZFKpkLAKOpmyBVzS9TTsYb49vDb9ObmVirWCQU/NYD9juuyeKtGJndn7q+uF4r8
jPNr0O5VQAUCaKFO4AUG7kNESonv8S9apM9A6xNxqfJQMvDPdo+73p5t8K9NKs6+
wZDw4lazDYnisq9cVqsm+fO5qqI5G3blvhqOBygJcPL1G7U8WaORb73DzCEVSgkI
4hyq/X8M+fk/AsnjDkURh63qMsXA4uoku/bq8qEG1gIvGjx7EJXcXyjFN/hec+3l
+u/Ig2J254nI/5gwFmviP17mFDSwVvopqpbZrolfLIN3yiSOYvN8SytmVq0+HENX
QwSLZ0Ok8CRWWVZWBdEyuGprbVi+Y3FlsBtIV5zXlItT5HAykQH8xVhiEU9FfFgu
H61fDRxuddWqxzhCeaM4y4wP2G4bau+8Nb8I21jRFzD/tOnjkQ8B5tlCZj4Ftqen
/bhvcliwFdUyi0q1CJ5r0M65z4R4HQEFZNJD7T2zVGQUrIrjKAHTmBJz+tSCnNuj
umtY+XgfpSjCMPv/sOKwey6SaHHcAgqjOwk2t/W9aDUAZnxflKw2Mf4Xn4lOsikN
qE0Se7ixnIspcADHT6U8w0Q1Nz9yYqnL2vjSynMRKzjM1JD8cKMoxrmO8F1tji7R
ZOmjoe+2rkjER+EA0BgdNOyqBRZ5/7BdnekYtot2p0HCf/idj24yh5i9ASf6/r46
jDEhuOR3g+Mg+zLtNbNMp1uCQc2aEgLeyXrcm4G2cF0x6OwcCZboV7+NYD9laIZu
bfrE0f01QFi9Fp+IoG1h40aAwYmrLazNqZ4cPmcuzKAD6ZF22v0rEQfH/C8C9Jjd
Kx6MuIOh/69VotGFYW72bZBTJPcQ6amv3RUy2z9Qm+tz5PAoFOJ0ZwxdosF2alen
SLQNadcU2U5aNd34ievYqF28RFFoSmh87ouZRPXGOD21uKi9RaO7ksjeMhyzNovs
Yb3Y9ZT1DTo2niWoOJKOfgO0ZDQUz7ecyzoawvkMLb8eLbFsJ6uWiR/n4+jcjXqC
9FQC65pVPMXU4h/wj8fDMbp93rZUYnZWkvpvSBDscTj4CDkz7we3TrXJPVW+ne9x
T1Thy3ZErF780pvWaTkrf+8c1lh8X3p45Y9HycfPRsFqApCH+z5RUIZ6aTh0UMau
2rSJVxuTKoldxDkOJlfwsBjYFvN7wTRyZZp3htKm6lQjg8nDLFo02ZC6GaOBgPky
uPQTYR9GgjR2F7Z9CHuFmG5jOpJysPbvyD2PM5Yo5lle9/NtZIJc2NlSkI7lfjs6
PzGcGAt5jSy5mUOdaJYKESEtxnPxOhs3qvZBXCgMPIU4ojojsF0Bqt6R0VsaplUe
mxuUvY/m4BfGNyLf7H7FSuT4wnBfvdI6OzLyXOMQvi6dNV69TbD7su5nxMp4lOb7
PA6HOojPCjL/1UM24L9r2Uw+nsEx+SnrSjSOxNxXxKt23jNP93F9h5GjUP6F2XOX
fVCEIM1ELaSqmboi74ozaN/Dg6814yQHFjNs/aIxmJiox9yUhieaRkxezGQjcSlf
ajS5YP00yfgzYFmgj1nNmxkUUGLm4ukOcC5jW/RC2stutIqdpAiaT9V2/5UC5mQO
dBwSokx8fXNN6syBe2Mo5eOL3CtLJxZIcuaVmkGGfqki53aJEosLECqywQS4dLZ7
8a3OTxR7NazR2zZ7UFVQx/d4tCYqL4UME15hji7tk7l48tp/ei5WbSfGBdnF41Ox
CinoxFq4i2rw8A8VCdjgY/yj7GBhaEke23cgIot5mspgeGoR7pMPCSLJlfRWKHua
T/dMdTVhYoDfTWHrhfLf5zz5vEgS7bJPzp0GRlDZbrXs3via0LyeGsePT5Lau6IV
0czzgOgP5VPHq/hTkQ2Kkn//S1T3SuukQHFOgyBxhwqcf39FrEdQ5JgABjvkqhoV
PK0M73eIPrI2RT0wxWDnQEoaLkCfN9uNJ8YPaPhM1uaNHKUJDTuJ8vahY9zwHbBG
VU1RswbFfaC0DnhXWwRE5bb9Ytqbl6QOXfPPJ9XkfizS0P4zepcigiuIYR55AcZ5
JBXE1hS2x+7OW0s8gOuzJFFTuELgz2ABtjNTWzvpo9u4b/js9q4PAUEgdpZZvuY3
ZovTDE/5e9Xn328IIiVtZoDk6lPUGA9gjUFbE1eBLhxSRcREb0kj3vohLYyxsUjS
63ZQ9RkxWqjfsgRbInEg86U81SwXxo+BGLofjiHvSSJ898tDkAMh3W4zA2ScdRVn
E7kMDoJjdYEgZ+eWeflnpJflvOIqU3yNG8UTG2YU1wCUqzyL/NlcSbEw6mfYvmgf
eXsp/XfyDD0ACLnbK6xudih8keOPo0IrtEyaZ2PzMfZv0uuRhsUjgc+V23TB409x
bG0dWyUCacARh/mjw5PnfAis6VqygUmVwj0WiR2g4ZwsXMZsOHyp8niJWj+pVU5e
Xe3/K+xDKfagtA0vRhUX2QYJ0C7t6d58NEVotbp+tGQrrfBzAxVJK5sDuHTIIUXw
ICl8Ed3yiCrWg/8qQG5xHvG5+Bp+oyQ5aCF3aW4WOtWD0xVkkSVtHGrfUPUMj47E
BPgiOihXVIbvFwMhRy4T1RIDIXsLt7fvzZD6qGZZyMSkZLxBUc0SLcFVT0LBhyQp
DtM9O3O/5Ub0dHIUwLM9hLVCjjD9auMPoXiOEQaX179xbQxIPizvBC0Qzy4i860p
Jghipr6Vt6ddyomoQojBSu/SSaeAuIHpyQus8lZzTswRtbplJEP5sxS0eclMaN7Q
f55VdH558JV4hbRNrGULRIqILnXXtZL56tyK5S+mFAb1K84zQaCFB349re69X4ui
vDSmZOJvIrSPazN5k2Bc0r+MM3uSUeRz6GOYPeKFlhp7WZ2zUc50UqTQxXpLp1Uy
B55egiBd0M+hcqK6/z2rwibsn6uJxWAYlqAvGz13CfCcUWlSwBDlrQ1/VxtVtzAU
ViC5uHnQYokGQTXOkhFzf7zrDp/urV6xX8n4Cj+ubfXSr14cgfVeGWJsR+T9bbIf
AO7p9vQWmA8RHls2SItS6ilmLcVUpqyTxn/l6YkrEb1ydIbLl+fC1j59t2f2nwtm
I4CaAoVNUiOjlP5J5fhMlH/jav1sVydRsXNYFwIe5rc1UgkoiUR7JjD/6QkcYIhf
WI39dpMHOFR91A9BdaW4meoeDMusD1HaLRAaWa/I1As9TORvi8YlIw1tutOvl58n
X6bO0GWGHuNe5/HTsSBUZI6l/Yil+sejqRNN+UzKANMTfaGWUnsJ5/dCcHYBPGDQ
ukntjFXIMuXWmDlzWKNrveo2JfTs3FfB6MHzjneXHO6yIp+KhoL668xgRyd086M9
9OvJE5xMssJTGVgZf/EY/BDt58IM68PjSHvBXFjk43oIpsD0j22WLnT++ekVMy8I
cRe74QVb8trigpJe9bhzVteRSrsyjz+0B/C9eGoD/FnI0U5yAljvqC1ToV+SBnQY
bhIjc7wdELrpRMWrj44UjYZDRr4xhSsuL/aK8q8xshppEvmgNQC63KBkCvYkCZby
eOVrro6zHU/Lu30YXpL3XLBAIucZF/Ls7uQuU7Rtocb4KosIsTGF21xAkhNQfZ7v
sp6lkAKI3psL5IvO2lxnu07+IvhKSbInaas2eRjONAHnV12BRIhctcimxT1qpo63
LUnTTXDA514JIDu2t3trrZKvO2GZALFra9by4ELZ6GuaUjWPV1pvGJnUxznanvxN
lBsbet4WAjcZb1rpzTSpfjFLNjykIUB+61E3BUhccB88TBT3a3xCnH5hLP69UhGK
V08pApupDAPR0F6i1lLBllnpOVKntX5OhlCmvRunPPOp/vebR7HwkcW2+BnDaP4O
YYMJjQ03RwALnZCjqHkhjeqkaruktfUvmLaVKvcj18839R4UwXLOcjHB4YuWmXMQ
s4LicFXlpoVTDPFKL0BteOHy4ddZR0wHAG5ZGZ9mQnq21N0H+I2EeYZc07Tp/509
ghvcd2UzL6A5YOhCRT01435uZBZIEli/NdfWxFVD8T7+WPxdGAkdNvzwvw7SCHXp
//bAupFGZm2+zxAxaHw9oMg6EfONqAG1trSjbGOtB4d/bfZ0SI7fI0w6nXo+iizE
aUbs/UCWXDKT+0Krq61rFg84M4+C9h5zPdNcPpHi781d4l2FDgca28g7XD4gH+/H
cJWvv6r8Tm95HV4G/ikwPiQwtIFq3pwqWcNw0WVbDYTTsSHznp8y6GWNbyQfHCBB
j+9gf/Mo6j0FdrtAAhXU2tg8Zb/zzGBeHSnk+GFy8Z4VBQzA0EH7+Zh2BNQFhnSL
WVCFxfi13o2HupmeVHl7cDNXkQsGoHp77LN89MYIHkGs3i9GdH/SCgZRt9+Z9cxU
w/nMhLNFzjW8EnkG+Q+XqNH8RMJMQ4nzDqaCEIEN30QMJgkkbzMyr/RsujDmTpKo
TQd/SbLyTV+I7BtdF6cMOVSny4mQE7TjBOD9q7aTEe16gNZ247WtE26okxJ74+EH
KCzooFzNPn1pn5i94pr+JNPnLDlUYBRz8OjLq6LCWpt71tQ4wQjpilEkhJFNEpO4
H8b/OepHCjZpiKkeWHSSEpT2yu8D3TEdp500Mi3H5l7U6dakODy8pgVaIdaI3dfc
wbrOOo4G5Ipb5Ct6tNHmZebc05z8MotDePmVBGn4lA8ADdAD/bqA/lYMk45kBgpX
PM6WKQ6rqpshHSS8hdXtx68Ryogw9nzOHxUb7fVLjVTfZF/ANkPUNnhJdnf+Telc
exXyV+huIWD1KFTL3q/jCP4Dt/cFwH+FBq9IhKnTd4uA7fTWt4NMk+ATaDWmQx1R
TT+mfr/vNOynKdCcvzvo44UYWEvuPqSIuD+YGeIHxQnm2lDESPWLhveu+qgfrChJ
5v3OHTR6QcaG61TrbpeEB+oKKUfOcjV76ONqtP0c72534Wx6gi18Fu3vgwukJiB5
gf4fzoGOLN5JdC5M0635iNDwi63Lw2Hq5fZt7mBM/SNG9nzEhn1XkZb6FanaBBtn
t/+zn2V7UxHdjhlUFFBkIGZ8qK86nvINlesE6xiI1d4wwWS8/JbNYe7uSfGgydve
gJeAa34CLlRBeVUHIV4uuGPu38W9eGOi5MHxUCkmYVqcGv66WnqXD3MWCtzBOmmW
IFEtSHRODcpZwQIvotyUsFOw1/Mu7M0TF5kCbRiUv7xht1iYNhNxlXhlnLbzn62q
VtQSLjGRzRq93BQpmuCxpOS6CU87NHI017jczr/rbZCUfGhXsXqCUG+OMdVAFKsM
Zog6ksUxICNtHwGiSRipPSHJW8HiyTxRHpIaO7BNvCGZDGUDQaDN8OExmw8hT4Ga
S4PDNe2ZC2osyaFSsz2/qZkJuq9Jy4m/KgbWh0zj5dtwssXq3NgQti7THQ+HEQCd
Dd6YA0De/noYw3manqE5c7UTqUQRjmwmWLR+PrI6617mlCqxPWj3KXPx2V/EMF5m
PQu3ROnOWuWWn6Ce12E4lCZi2smOndQieiK3/qSJ6t2V+0QaKxYUWYD7bHUzbJdp
oAh518/kwPFpkwKH7SQqSrCiJ5sQMKXGV+Kfv+Vnv94saorvgRiH6pFOZC7Jr9Bf
F2921aeoMMtZjM4/s4Kd0m5MOA1T+4M15rE1Ph7C3JzXJ05pmgbFqW4AXJ2767zO
E2IVEIlrLtfMvALu0zNtHvS2MFBC8mZsIiBPMpY+pTaebySIJUfQeIY1a6fILETe
2UMnc1iyhodKbIAaiwtMY24LmWAxI7zLx67pSTwjteIcsR56t4lfXpz0IfLfWEtc
cpEw1fV4YJYLyGGljuEEVcmPkbOyNMeU5HqMMciqwdGfO0cSzaN4EL/pTiShTFH/
gpkN9XP8kPRKPRy1lYQ0dHpNI0VJEpbg1i/mZ2RG4+ztD7CvcyOav+N75iMgAMR5
Qj0mk6d2X3ZrcO1hwsWv2SSlg2QZKJWldXzkfDOSYHYf1kpPB3Fuxvyrxv6kcG96
ou8Xgw2DGaKt2cgAqT52ODmKP2IrboHC1xCQjm1ppD/qiwn0ro8OuaPHiHT1fkYR
B+2nYQGI3RpzmAydhvkKTVEKDZtgHq5N9wyPxGj54RI1syDgpymRx8jTBE+TcMdC
wvSAOYnGTDTFfmMUMAy6R5o4+LSpMhEz+VsPLqhnv5OEkrig66nEKolliDDaqMch
Vb80PJV4a4pFlX/tkORLPt1h9fBKsBIyBCyyugQhYqMjemlemNmotfstPSQDrzad
1n/Rm30NLpIlYG7goCF+TOCb865f7iZ34GixMrmzk/Eun8pLVo8rB3cSZ3aSqX24
uw4R3H0yq/49G891hlp7a6Ju5EdxZjwy2wD57pKTmuTAk332TtiYUrC8K26/MS6E
qbPKpkSeKbjEMHkivltNAo6+HVmd8I0o4Bdv6Lvv9OD4s11JvXH7xoDsEUfeNqIa
/4sZtgWL9/p04d7C4KOQEmMiOYooaxOY1veLV6k2HFAUWM4y81iOT05NRoZ9mYRk
fdzC76kIrILNxPJGaLUY5iZnpCeQTZZwzIwURJc+FoMmVbFeO0y+rjKr41h0nJfW
+GG+A1l1+p7QEnbtm4c4bxrjxsYstXDw5jpifPOvA8WIjV4/TADff6vDxvtUni1l
bA1ezNhbUsHu4uGLsOfOpVSZfTnJ2vod3WLSREWPXvDwdc66nuY8abtivuQbMGNB
BQCf3JiUonL2QfTUtF7oMs8g0D7L9PLUU3bNtFrJk5W9xfqEf9npcAyIdH+O5epL
DrxbWbBQ/RIJq+e9a904VBYb20pLrMgNLCx7xqOb6D0T5Hc//V1zUGS2akGpO2oQ
Kkw7vEEJkb25OFYTatYyGnw29lA39vREFQWjyINhfbPNtd3mdpeCs86LhBiDYsOO
u8c6lPyCiNO7bB1VjpwU82TTRg6wZzC9hw/DrPc1Hu1p9dQ4ECpcdoAYNLDdF5Dg
3sLaGrVmCjq40lS3oiFuPugvxgdeP2qkU6G62WQH3/XsXxD8vZvLrfWD0zHUA/7V
Gu211W+53IVUsd8ZacwLlPsB75j8DbmBwrSVHUiHy60NKoLxyhNsdL5DPf4U0nIi
zijFnyDsV6F3F1miHY9FubLU6u6Dna0Bz04erhrmvgNR7LdPA961vBB2IPxWohDT
lTNxlHuxgdNw2ihpyg2K4BdwLaKUPKXsF9VsBvFqoLkBlNzZCoxTAaIcHA/SNDqO
X/XaUoap59WxiUQgLGxT2EzaivA9O77KUlQaYFjqjZ/LoA4TdttiVydmObIUnpQP
PXpsGcdrxKZ905eRRSs/H1pJ3B4VETLHwMoaA+U5uymG8ocz4BXlgcjAJyOjihwU
czyxb8UNtffdPvX2rIhhrw2ci4yVUeyWd4qIpdp0q/oeBcw8N2LKZb+/DXS9IXgf
WDOctxUhzjpqKPLqzKbyajRwP4TInLpJhxUkVFUuZtb01aS7LkdgRsIIaUcTJlQH
U/8JQGzEqWJ0bNqIAoAuf65V21El3/qy2zPil67+Lc81iL1wef1E5t//KPxAjDGH
ZL43E0VJ52LEYl5c5w+hHYM3LR/ykt/i0r43aGUIWt91K7Z2PF1vLlZQVRpPHwUL
JiPxGufUlAv1QErJfqxt0qL3VL5EJ2hT+oaN30+GAp4//51sXLGg6pb+3dl5p7da
mRBwYwOKXzVltzcH+vir5enGR7wSH0e1QFkkZHlhdMbTuywyZ6YIY7lGI+x7HZWx
R0U1/6X5jreYx45R+oKVQS528XqEnTob9lyNhntOSYsuADt2Rfn1RGBvtdwEnX2W
enK4X2dXGsC50jLGVew0Ono7U6C+zGS/LUSzXjYD6PBkuRF/rDUwTo2umHGGsd3X
Wg0yj/WgknCWvaqq02AeBXEvzuIBMpbRL8dYuCCgbMz6qr5zcMj4SWeSWyTJE/Z2
wv0Kuifqp4+QYgpNB1Kjarodv/gLjhg5F2lgAlHU2aWoYgGsBF9VXIamN48Gjp79
6ka3eNIvGYG7Z+GBMANbuQYhVGJLLuN4NGkeU52dZaeffmGPgVb/OT+JVUGtbDH2
Ci7s/JMWhCCdNhpM5Tu5anP2u+Rlf2PqTeAOJZvYptU+MlXYkRj8WC7hsvdfzNRk
F1kVEO/iIPD9ooy3dIABQ0oH3e8MYIXYnOz18a46/aNmcHm8EgprQp0SfFXQ2Rt5
QhVXjy4X+ki+/CEsdDowVYdLcJDtMBTAnOXYFttRy8zV/AT92vJ7K5kvmud7ms6U
4408gOC6qNFNzzvoaO1VzbTZKqhTYzNyp+XfPijx2sMY6SudCCRvbWUe14qUMV8r
3NxB+SVTvrdlTKhrFX+qFkA/FtON5JTNM11wNisXtPXL4VAofLNfYUt2R7TVrCu/
xAn0uT3gzEIE0cm266rHv3h4H3HAirYgCNmdDvLwEdT0Co0mbl1XjSl5jDB4yj8q
ytmO/OaAxPVkN0XbLwrqG49HjHNol6hM5S7JU5OpFuxiwmzxXQMTBGq7djIv0Mss
I+G6VCv7UZgAjhfNnyGf8sOh7UPyNe1AwVNobiinIQGa22W0rjDLrVXxWT4k8/c0
TKqmZO9+h/yYuvxRT/H2zZA6viXOfbwaaBKNdF4/Ve/787JJIHZzHFlIHu0D10qg
NbMZVwFnfQ67uPoL+DO8sNWj0KESXKUkwBU8nOrmQkeBGOJVrNIm6igfr41C+SjC
fH5RITv2jAGjmx2fm5AZnLZZWsYTmerHGTAd5pyKRC7AVRl0coA7Ck8alMt8LlpI
JL6moUa79dTTNazN5b4Nzu9Jua9+Q/4HajGHwdq8IyMBAwYx4p/jC4e0DUGsH/Pz
aij9Wg2fVSE7r+MGYWT0njycdU9MCwoDaJrVVeWBLA4C1BZdADZVa3+FLVFP8elc
peRzZ4AaZiS1Fj6B09Nzik2wD3GvDzUWkAmOosYtrf0wBKCQAzPqGFFJ/n8/RaY4
qVDVVZeMKrdAlQc+Apls1BcZdU+PNhk9WUhRHc9cf+dmDsq4HVpoX1Z802j+6nR2
UqElRLLXqV8inQcsK1Lv9kBUbN4Sq/u24pxDWLn5Y8KRU572L7njJMrJy+SYCu8L
UyG+goyXU1bFIG7OSjAQnD8cok+mvj+cRbhzt6CSHd8UA8zxWjowNr9L2Aw3028J
2nF3Ket8llkXt5RqhZfkt4l4dYJm9FywZ7y3iOyE36dqi+Y12G/8w5MXrkVCzP24
PSyKjL8ZfJcnLuj8UpZxfKAwnFkBxHC1ERddizfVswVOCTs2qMosLXnR1P3rIvZx
MTE7C/sby6Qp83PL7YHEL0iXEVE2Iziyi0RTHJkMvj//VqH3aGNdDgmezzcmFZaw
t1HKGMDoaXPZHbqgpcjH36nQdoKtyk7uRwALjUGL0cyTSbIhykuELKKoYjQHiAZo
QvNDcelGMyw5BNU2zDcoCq7QDDG5pi4jkA92snm/uQoYFwcDAT+fRt9V87I7mT9O
CGm2ecMNxuHZSJHdUiiglO5F7PtR/s+0L7g3O2zMQ6LIAcVAmy/k+xbb5sHzVwJo
jGzEJzmQ/D2S+8GAxJ4I0JVR1uSrxr9Mg3gxH4YlFqiuOY8BMf0+yp82402qu3Er
C/OpXndIb+dOAmpGTfJNKrMPTh4qW6pvlDhB6HiBt0ZNDHSCos7KKGWxOfmXoAQz
gGxG3zbSQJcWoAUkRaAsezJ3OBjkUUCLZIRyBctjfKA7uBsbJPN2mHabzayIYyfC
E562ByNKUX4dIA37r7b9hMWGCpJtlnKO92SKM2PUKxRt3SuavzfTgLZqJqX6UEaK
M7YGDe3FueNJrNPGJJOb12s7X2gww6yhStt73x/XsZjFL63bx9R5AFulFljG/Ddq
v1bOTJw6ei+9sqpNH6uanKTv9dG/J8vOiU07uyn/vl1RyKeJkM4YLWT6rJZPTQdb
8Yh1ByDHZbeFIWumAaD2SghPfhay4LsfsYe0yamKvEutXdzRqi8w46OhO/i4AfgY
Oq4V7DsBpmqJrXNRxr1Nj0PfGwda+Q8d/NA7eiullJPs45LEXsgyxzLVkBMNr5Qw
xP75Q6DqR7vS1nBt/Uu7uyISJAX/w8wDoDzfIPSUdUGYJAxSGe4+lFWkxKGVRJDJ
oFbTSaClb48u7z91zstQaR6FajN+dgw+Bg4N3B8+snJjDukXpP7srLwZ8QgNwXOo
FYvcaVUGzURP04uA6gu/WcpEuhDRZAb+/Mk0yIJkJWJx4WkhGk9o1ype8jZT/fEK
x/3B9EctU+2s2daOwufqbnss1EMKofLXfBprvsCz9CkGa12GPBUP9bSanHBnsZrV
leyFmYiwbAt2et2xl39G0NFGVrgsGvtAu4Du8r7+K+EZIQilu9dR8pIY1dgWfNzg
P3M8voQT7NTT7Hv/NQzt0v2GGY+RRRIDfqpWe0zQPqIqha1v0N1T79E2esJM94l9
PRT38WfADEMRRkRAUhsggguCvVB90E4FiQBPiy6hV2dMyufowiW1mvzSgz6Oujzu
vVcDban4g2U6pMfmk0/cqs34UT+YQwBhMTn0W6X5t4jYMNpRuEI9/vXPdr1O+Emr
2VawPcOq2RN2812AxCxcp2l19xbYZ7bJaUZE9PTtNgHWx710wquAVhIVY6tygdd8
MHbidUXEta3pcBEDPz4x3gUSWqj3okXDbUQI3vX4zP17sKu48Xa+oG/pozT6sDGo
BCMFlAqm7Ya8WFc2guxzIkfmQq4K7OFVRHkXHkv/RuZ3Ztd9acgv8rqOv5iPY+nt
/bSUYmtT0ulJ15Dpm4SjU/joMzAr2rLbQeLFzab8TLp4I8ZO21SOWPyadAtRuMC+
/W21c4wTiJteRTjjUtSGzIjMtovChD5dDa09XxutWZtsgpEhioDmyaU5O/4WFVFZ
wqPaVW7d/Fj/fXp4xypYttLC97a5lWe5o8VKN+SrdXF4PRE+9BNtjQ1SBJcFV5NR
T3m9wzDvumh63+l7C93/PJwCtWEwXU9QquM0D7LbLlrgpcq7tMPVESqdKcxN/kx0
DhTxqnfUZdldrRZLVCe5IRUJXAlktboXZL7LfAFcvtF1GXXw91ZOtUb74Ye+0vd8
K0DCJL2VjCx/X+vZ1+HLRKple0Yh0NEv5l/nuOGbFbFO33w5Wb/5kTd8yEGmeDMK
iDEAkrhI4nWdDzumH6K4ykVta2UJmjyz61dFcAfM7Bc5oWRSshIX2hEsOUm+Ribg
F2Pz2cgrHPkixJZjNeHubyJRk3wGw2A6KPHQdA9UYy4hlfplZONuh/TRjHOSIbLM
jWGbrq5lNlVxITBhrgzABHcbTO0WCebU0uJtP+7dWl2LEDfcC/0ntoHzwQy8qEN3
vBEWROg/dkKFXG/SXN4otj1J7ZJOJjElQffIXsu2qMhD9kWdoXFj7KRIygVDfxlZ
+D005DBtolRa6fA+tcAHLcuTwwf+TrI8ddlsVctIYDc9cbb/Rvp0V3TQABq+0BMs
qnQVY6A3JnYiycLGX6bcvi+dUcwOKMFT0p1H7MeirClXrQndbn4BsZqhH/dpVkwu
84peZitlxiU497NNxlYIsLitEedgLT394HzlnPTyve82hllD7tMXt444VNlhfsGG
RB8SCuMZuW4gd/9OgJ/gNcb2Z0cQ8ZkhEyKX4NlHy2DAcvPD+SDAa2MloFJPH8NN
gQ073UAByyKAisohXXy6b7kYi/nuYrCjkEDKA5J5RbvuRq1PGrp85GWN/wN1kxe9
My3g7xOqnCEwQKXBNUol77+P4jgjwUWogMAp3NnjRTESFlx98IyJHiX0UH35ABbn
4AeyYbqCF8rtgq6bXHqECJw4qDZsZaHI52CgfuUbZHe6B1f/XsrQa1rNSTI0R5xP
nvr1TkfePEAmUS12P24IvthbwfaRyF6cQSNQsxxuZxQmBJ4otzKGV1GWnSlMvpZ6
+TJIwvUReXv82VCybfjunGY5Pg91gDO8kWhe+NwjOyOKGPDOCuzIC5IBPuaPFCvC
rKcuVOaBNRCyOUvDoctTmxv7fU33xpuEh+tfSiigy7hv790pAwLFgLrBIGspmHPU
TXIq3fv0h7Ta9QpeZmrF2GJWTwegE27wgHUuH2FHXbphFyqgAE3avLOxEyiMHZse
W+Pc2CCT7K9U4aImOzMt4q2LzAiXRN9wB/GZpcY4gNcGBDLpwmvkOejxF2k4qSaQ
+9sjqvWci0ARYg6ryDb3YiOR2tMtqW3SsaxEV8/DTQgoD9xz9QZLWNgyZO/d//kE
uhLNjPqVQ4HJ7RzQ9bpvOr11y168mpbrB45GYLYs35gTFTgmhEF5CDJmgrCm7c57
gvFP8qiSxK1nBNoar06WSeqxOJIzaEhp+Dg0LtcMblKa35QXNbduQJKD1W+DHBWM
iN7H3NYAfpbGr5FNvus16ZJLCumQLHl1uzwTas3pK03pxoRw9up2Q/xaptq715gN
SxgcOGlQePkwWvCyFKP5WgZnUZ/dnEgUfBseeyhpmS9ZQUDezpRtLEm5/rK29EVX
2opjrrWFlnyHtV8npbycYn52dridz9bkRVr2LLvOaSdXwMW8S7hWprCazruU/WjJ
nm/UjY+yoEmsY9Z+7SlE3ItFMFtVRRYohh6s9i5ezjNmYOZsYhl55PP2ArVQjibO
slRlFGES56CaNWYHnviuAR5fkQUncqYzeLFDs3EWTdDFPh34eoxZDx417OgVPUKO
if2f/tTYl7nbSEV0f9zqCNePJLfT92/eOCm5TUkckCO4Y3DJdRtE2ODCeb2fmQoE
sog34yzNswW3KNNa25BrBl+Xl2j+UOokJQco3BpSVuEKSUFBgFdiy6NlvL5+80AJ
dMgm+v4rCJW2SfnnPiP9BAV5ARZZXgVhv5To0lQSIIjBnPgArU3On7RQIrE3lYzH
x61r9JrHtZE6x59bUTV3G2zIfnWtRP5uZVvhfpK+qwDQZT38aTBs+X6BeIhS4mxO
97FVUIcv/ZqZKtqcYkieVKJQB441XwZ0HAUU9CQKHlFhIHzQcswqgNJ346P3caPN
frdv8XCktYp60tJ26Yy+pBcZKkbX0o5WxNba67dhMb+WBVWXex/1TowBdfh2FxmG
TYcVsbanOggrlnIq/IUk9RRa0MOXC5t0oOCuR2CRcn2tfCQ0HQkeTsvz1kGK8I2Y
d9yWUxW98AfKSqHDgtDEb2oQ49/20mKbprl7z0D0Tz06+AjaFIrzLVgq2hVoAhR6
IpBkbrEVoOGNnEuLbhbgNdnZmkC6EgItyC6lA61lGKRkuDP5Dp4rKsyd3DCetlcl
27a9b/Ey9O5+U0qpTbjU9nGuPMuf51sCHzz7wGSJNzXXvUYYyuiOT9U/Dn5CL+tg
722/X7qlfrZFXh62USb7I0kYEHJoNaAsQVrnwuoQhbUoXA8NDGJZQlXn0j3dnyi8
44C3t7MohnaVsPHNlalc0fAl+sNhhqi4WgxEp9smUCoQfV//XhyQM6Rn2gMh3vh2
liV3rL8mV3e5Bvbmog0Hc7EyX8K1JWoWcii2uVOi4DdDDj4Eog5uCzC7MMdu2Fzm
mdp6Dd34oy6krsnctQHuwNSTTCJleRZfpPh89tSHQwMlXE8Ea0dFJzlE3Ul7aYVk
alEpQja4jjv2/9GEdXKsELYcLD8qO4IYline+rVEolXADYb/WDqDf8WG4E+r2+jv
QthXjdCXOW99qN5FOVos6Wnal5uqwLyfIVBsv6q720hq4WZFDznHouJrf2AMcnwE
7Z9yuBVUxUFZj6LsRMq/VjzjL+2xeVeDqomM/qcAE3lZCst75+RMQNUJatTdxfpP
xEvGZ9SbuiNvsxl6oLpRcPLp2CnXuCWsgjjFYVfh5HmnaYmSYDtrYt4+3tIETw6k
MjHlnqKAtvMf7J1n/lG4PkOFD19EpAr2TYpt98LblvjsLnJfQ98pjbhEmrI1x8DJ
Wl/zQFNae96xazrDU5NRwkkHyHEig24XM2jcYp5Ew/3u67UatX4rgQkiQR11M98e
u1tAz7UC0JKBSUdDe8Bo5X+ffumhvmFJiWYBTySFdvacRudHoqVaR3L0TYtP5YuJ
bN2hXZNn3iwZsHupsMZ7fdiNoRh4bXi6IAmre93TEcJuiPntBVmFpsZtHo4fPwYZ
D66vjc/2oQn8t1ek5MLIwkqRwFdFWShYAqf4wSnz9RbxsfCV36cP3IeFssCYboRK
/xf6tKjS9+xHc+OWJVucWC4Im8rQ+fFYP40kxoMhyWFx4NVZ38eODnd8qSg8YnBY
mXirQ8TsF1N18aNFXclF8zlt6LHQvceX7/OyUYpkogNu6azpZHEPWzZBtVcC5pxn
RVlRGqh0yjYZWs9GadYgy9Rz30vnMUexcoXC0vF7aCn2xPK6zNRfG54IKlg8pTds
9INLSHruEzABH53OgZEfws+iHMA7GIRg2Jf9/bgm/s9C1R9RLiG+JRGHgRiI85Pe
9Jhvsf8Asg4U2HmfQW5LlYJOtwHY9Fj73AwI4cYrNItck5jFa7R4x9UBq0w7aK0H
87mhL4kgpwrVm6iYScxeDipMpUE/sAkJOf4Iz9ZoaDk+XaFqE86oGCmDApidqkgz
1wkDJKsz075S6CHK9+P0aXUTCkybNW5V8eiFRyt2xbe0Dz+eheTh6I35eDSElVrP
j1OBsH0dgKMxBbQp79H6lJbkwREpk5XWu6hHVZ2frXmAjNU+ebvjIFGcOUTGOgQS
/+q5tVaYnIw8gHZlD76YASz3xw2/NJpnWwQGD6pShXMo076vhKhNXPK/CpFuFepw
PGR9SxuVTjUVsKElFlRrEPsObqhV+eaJkmzNhqKidatKnQ53Mk9EcAyTOZPZxX9h
/Kb24+EUG0/UnPlMITTHUkdCn2mVYs7CEoaSHm5xckhZMMASdjeq9dJ0CXiM64+8
QraZm+aktAfRTkA2gwBS73G5gHyxL7kghP7JYwAS38ZpyGkngwq5MqiA9IuXEjmB
ueejGq8Diw3xiYcthVAptBQhjtQQTiVxiHUZ/wvvnmMw69o8TreoHk1LfkhUJiUn
ez2z81LVUzA52X+YOMlfi1v16Z4cPYMZFsBkQ5Zmso5lEjeIDvAVxQG0+aEYWb9y
1RrHNu/GRP53jEhtGd2n9AIPTYZCLo3ga7HKoDKjmg+whmTNfpJpm/ejcMEC4gBm
uNPbL81ujk1KbTVZ8/v7uzK4siT4gJ47fpfAyFo9Tby8PXQeFehE4Wyqij6uTmmZ
8kv+iG9YeLSAlOjdSqpnr0CgPyz9iHpXv+lKyNMFtgaQU6EnOgZJjyylUIoQI0uG
AmWOK39foY6ewURHy4feGyZpnul8UXiNdgXqHweE+/QdI4ak52gxzy+K13Fg9AS2
SYYBbg3OGzXmeUHfpMifww9cmTWNLFSb+dV/MDWd5NhNFlOYyuzv0WdoVkp6H6zk
1JcsIiVVgfnA6z3/Ph6XmflPYer9dLexfRrkJ3/3VL2fCssrHt4ZMp7DZLFa1CPZ
frlM1HvL3kf0VHtFucvaWtX8wHUYC7slRWiphftRCWHuaWJH1GYdYPvBr1YV9UXQ
ZodBphdUG9BaNSGJlHurkLCdV3k2xV9J9mMzS2FDZzjvHPLbJoGhs/1QdA8tH6y/
ZUXCHnodkI76erpQsX0bS7NhgAkOt8VpI6qHio9dWacAeUgqXJeU0eulNqDUN57B
euirpqwElNnSIyfXJoOEbtH4fMkbGyS3u6jdwa82i3/8MsB1IhsajbENQgglLzxO
6hQV7DCw/TpboxFgaZlSeO6G1FvKkPTs+lBWtDQ81URQESblNfpiM7Dw7dy2Rx7f
8yEnQ30omSwjUjByPKpUO4cEe1NZYfGwXJPojxhjFTuhvOrBXWyqq+eHWE/zIMYM
PmqKa9mNXolIjqpeAJA4A4C64nnnP3vqWVAcW4I1Qt61NySALctbVFgnePB/7lHP
XuvgudN5dXATrYBMH+8xrzLzR3tY6UXO/7PzHom8FdRIYD9nq7OeWEXRTEZZCPJ4
/CI6TUg+/vo4UK0OJPCCplWWKNRYwhENLXleEFj6Tb7W2yIZERYzo4FQ6LljBVIc
Os4idIy0q0/uWCKm5KiInc+G7M1KulSJjmz6POyD5JVODR503muHPSULs6DWlfmL
/VhegbyISrHIrk5MhH2xIV6SLJAOyuJRsXnxggv1P5mi0S87HYOBB5HxRTSTlysZ
sHoKMfeDB+jA+tqJ2IsXVSvptql2bhuz0HAzDzeqqp5qBt8rvND3SaeK9tXdAhSz
d8+zmzCJS8UEaJgZqXsbjjvCY7mX3zdCzY3vPCL1aUbuG7rFXhPtT0opHWIWojrY
XIBVPjqR6l+UIO+DW9qmm8I+mxbCyHwwM3gf1B5qqvFM33GB1lt1d3tUbcIvBWnU
0JM+HWPmqseF+p6Ms3mc5IvXkhomAi8q3dKY7qIbLSfjMQOraL65a4ATKsAkWkv3
v88HN8VudThG/wV2FuggWwv1iBBXx+bmGRvLWAyP/TnUZIbCvfpg8nHxPfuqLkbj
NdO065f3IMQP3vuUQozwRK4R0+S/F94jgdBmiHP7ijQhZMdgfJ2v400mjn6knojh
qcPOwpfieANU5U2cKiwftgHe6FVP1NTswxCA4mHLWh1UxuBQ2st/jmi5q1U2LHyk
D9GNY/u523U+d80uQ1GqGAloZW9dRSDreJx3rzyh1ckVhfu6BM6GLypJad3/qGUH
1uviCkF5UvMAJxDOC5KK0bzGjSrhT6qarUZt1xkuUm5G4vb+6mOPt7eCNpspEbXt
O53Qq3UTDuSV+B0Ah6Ir+oxS/o5kkWvss1RFuYq1nPWDHLbGsVgQxZP2oO5wV1fr
w2pXHT6W5YdDWlzbn0tLlG2vIcWxtrjEC9mOVz1O9Gho+6gqsw1YcTcpi1tK4drS
vbegMLkWpIAFqQZLHDxv1w/ofOs55VJSCBEXj5kwDQWAaYsN3mfH71o1T80rkXXq
jL6gWIvoX8M9CiBi083a6OAmm2ZyIXf+Bs7NIAKnbx3Wl6SNH79ydmXn9/jM9alb
Ttq1XEaNm5XwMk8f7bJbAtveAvwTvLE87vGn3rwXDrRt1RJYk8Ac7yJOiNtJb5Gu
akZL20TGXsfmRgeh5ry3Z3XcuUH+13aoW+lUkynB4j1g0SOWc+jS6p14apErBmcb
+xfVGMrZxxLfZyECepmLAK4mvWB0081niNIcgIMLu9h3E1RR7av7HgU6fN/L+pFr
bIqNwIL29/Tfy54e3vbBnsZnFUjmMlo5Er0EGvJJ3U9LRgkQsUxTnrPHnVo8vVg6
rwYmZIcE3dzxelnwmrfah0w0YlM6gT8hau6qoL1QdUr5TH5+NlnIFa3t0K6mArn3
7tjdPrBr4/7ogTPsrUA5pOxKlWmb6/5Z87gXMSDymM1C5DI8esDCEOYC8OB1Zkwz
nrsZgqnfMF+wkPDfSHlDaex4Nu4EEqAGXLQNFW3M+03V+7ZMwRJd4xi4YsGXNRgU
6AdCKQuM2c+PI/noSbuT0fAFfS/5RkIGWdpUoua4UGGsPxCFt6Pi+ONX0cHabr2Q
N4J6/+5RA3kAs2J/HL1O9KWQ5OjwlzKpF3fQFln+dGbNwFd47x6H/Hg8gB8WImgr
eeNjpkYe0x0OBeMkNuG5CcDoQJvaMXzZ9xsDhwW4vCnFNXkX1LYy2vgOXPwzzdPJ
mfv2/Xe1gA5dIip45+zqCziXUqhILeN7ulK+dLXkIixI0vCWHS5WtARqVz4Xk8SE
cRPm0OnJCIUQ6SseOKe+ha6LBo6sMKy4fzhddr1FWwswFRcg147ti7Sam0BDpVlB
vLWGuORYOlK4CZoy5mFPzsT3oSxHaXvFHyE+JvhCPdmHL+xTm7O96NRdZVB3hYCV
53gYdvbEMhwf+CHTaUDGi/o7xdgU55QH21RXCNjYh59RRwu1oiIC+CxBKjUOuqmj
fARgwBoNtCJh4E9OgbXTpNZedcmN2KMjpc0Cyh0R0NQ7MvoE7J6yQlV1bawS6+vA
8FrBUJAQNJHWabpqLtDbVP4VkUXOGW/8wzUKvLjDhohRTAC86kocbsIbGfFO/QWO
u7XaMSh5O7ZjAFwzNivHFO5MTYNIhekzDEFsVE0PJ7XLj1irdsFf2pl2XZc2llSo
EFJHPUa//4xU11x0S/YQ3z47Yh6ioBQ6vhWUpZdvSyHZKn9qtpyIw5+nFGJtOEDM
L/iW0CIUsBP38Hw78Bv82/18wzJs/Dov3pgpewcGJSPoBhwS57uICg2FGs64M41T
3oL/gPbD6/fCh+qjCKuxN5PSoiwG7UPPhOVImpT1fFVeGJq51rW8PZdJkcPEW07K
7YASNjXmthUgRLC6saqPzxVIgfwRIc8iMLxmcTv6EV13or76Qp2O9KvIqHisYo1N
+J+YxYgsV6Y8ysm2claCywS+zz5bX5ty39lCI9V5JWlbSrTtpUsX8Ux8e566PPtF
QOaltsYk/BQwbMel5vG44S47x+TAWzwubCRlWTonDI8H93DFqHi1HRlDd4id14X1
HXu+KoIjnzmGFWmtywv+TwQRkp8uWwAbfJPZQ2jMPvAz+xU4WlWd18kyKOJ6P6TA
DU5zpmUbNZ+s/mqVLamIg9QIDGFxURCpGDiw4qf0U6cZV04WI+QBRfwS49ra+xe4
EPlylpATuZbWmYWYTiKHdApqE0gt8lxGeRpvX5Zx6EvxqXWuhBtkF6tO0bEq0uCf
tyMegT4MbGWZMz64FgylH3ayGcG2esFpuoR8gjGezRyQdGq/a2FA1KLb2xjFe6H8
31giLZ9iCeJa2qNjHX6ZJT2oM5Am+nRjGsInVxyZF9UakgylvZhQLvAufINU4ZKI
R2k5vxt+4BNhXgN00/c9X6hRxwRPsmVau+Sufm+rot1iiU+X6TuU015K0HI4hr2o
3HjD9fKAgpK71u/j6Uq9rr9uqE92x+5K2yIXkRSAsSmOsmb3Q4RcjqpffAHEU6J3
CtcFHCKU2aGKuCN0hb+HLVjrtbxsj6cpW2V0dhUqHiwrfqVE4nQ+th2UtYHO4x4u
tRyzDCDapaCGkKKXV3SpavDfXLw42hCmWSqhjUku/oS+IEsjklogfEg+cjelIX0S
CBw1fW98HKaLxwlCpyh+npSQumcbpJY2AsiaSLIgQJMmlTukpHIxnvwploF/1vwf
RijyZGvzpYSG0wPlx84hkdkqVrXWV7PfVeTKiCWk+laQzVJMs9ascKeZBxWO1PKO
R23bcq6/O3b4uDDpen9o/4KFdFGvTla8pm3aPZ+D4KC1Lwj4z3tlwK0Fj0+5Vz14
o3625DLZe6bMyF7v0ZhMfYEDcbHpfAlFPkKrHm8Pfgg/YuvXcDSor5dHZypA6WsC
T+lTj0pTfWjpgrSZKGfPKKX03j7wJk8khxVfE+GudE+b90zymqZVpfq/UcSG4W5E
hstVKxQxCPdojPZQDyvoT9uWNQqtQTFTx/ThMN1TDCh+wSh7HOMES/O2X2iNtIZL
wH89SjsYnDtNcOdeUDJ0XHZd5bHGWNzHc61CHwXjriXqvUZJ7KA3m8BJGPnZNCdf
BILjYHsOaL83+TCSMpnZvGEhAISniqiHKFKZxsKmVrY1lNh6ZykLoJTJUUAxedHO
7iancYfZi8XmxKBpfwMT6VtnPkqEAmIMOgeMnI1EDFjxze0Q1ySO7LiywKOXXS7Q
eOLOVJTlCOw3Um+lgf4mwpB6sOk/sC0X/DpqgllTdhzosAK7T8BEuCrCEHr8mHdq
57PkjIOq4nUHvbWE6VcYvSUOU0hD64CFoIFgsj+CvQXpGj51TTD5HxZP5g/rpM+I
MWFap7yFAzhUhyMOc/pc80iX+28K4n/RukhZaGU1zTVHKpvQEgvQNs+clqu033k9
efLH1IwgHEnCQJU+DDhVL1h8XwPo3/eHkUiQ10HoVL0DM1O7XCnZ99hWZ45OdTyB
wlJ4aG0alsBgVpvtZHV2hD0pI9lt/FdEZPuHDQC8cGLpWETRX6hUugiSCek2LwsG
U4ieHklwx+z2mZvfrsWPHoEsJPnlvwzoE0+ObS8/EC9hzMmTtQJvWxC30qWqinSV
2XBJb/w8LNCWB9X+h96JUiiDv3oYjD1xxY6jCJeBNePw09BdLHbreszAWApQpSj+
f1Olszq+aW6R+2waNxCqdL/YAW6x9U27M83V6V2U7S6EgU8WmHNwhC8Pdl6vicgz
dOl1+djrL7lpzL7TyJ2cREBMSL9PEIogitJdTp06RU6z1xwdNMtzwtYRULmslkhQ
8lxfAG0TY5kwNwGnvSrLQM1MoqLLCQUa0oMhbJQ+pGnItq9nbrAFhayzb7FRbtY5
pC3q0pbI2UWIi4pd/5uMPcj4QC1haoFHEGBN7scA7bHDGPPheEoza/qKYLaDL9NN
M0AfdHCX7AeTgFLcb6cR3M2ku/Bp+ift8IcrYHAtS0mkiAMowdeg9m8opSTEpHW/
KZ+EGcNxDSR5sv4afw5hG5N6J06sckgkx3U/Cfk6Si8d6WHO+KUIOyhMXS4Asvl9
a9R6jNCPOGsS5bxRFBOPAbevs8yfCokCPAC6wg8S902D7TYNyieP8NscXc6zCR+E
J2l3cMfBhaEPlV08yBhUt7lVhk+FMEIUtczCVIHSrNTS/uE8GYD++oL4vMKlCZC/
0t8CUwv0HF7OIMZDZNWHQ+E+kyB3ZmV1Fxvw2eep8raC9eLeKjm1GtLlTjmMdzeJ
E7dnrMEmYEVPy6TqEYwM0HbGdC9FBVyATRyKxXjmhyzs0eocXqdrIhric9ouj2Ud
db5av2NBJ/6nZ54ZgcWjY3Lt/IkmOkh65UXP/zk7bLCNui/TkXERd7W8Ynk50HAT
9Vc1UFuAwDJUnbXITYue2WcTbmvcml3/BFgMNWZn6HPuJ0IqaplkuhnmKIei4iqT
wBwvx0PDtqqilK32DAb3OpwPDOWSXdmDJhVUlkXAYwfxrixEloGahIuWWMIonuFM
Gi73iOaeI0aEMt9kzRTNBT2/RLr2/rOqYEMBI3GDbSwLLIX0BeGx8Yr2fqbpvDYb
gEARdvHK3V+ZOGT5ApAbl/KyhdA6k0AUwvbMU7w6nUGEJAOMZMFnt+rLz6Ncoeyy
pHcR6ilG4lleso5TtYyF35iXA5hjXmjdY6GNIpc4afI3fQvZLbob2QuEbcX5TSg/
bbSh+jIHdUykKe1VG1epBaixyID+DJZzYnmjGeUWEZ+l1ZXFRI+tKDz2PD5a16fj
OfX+lJqImWINiSoAy7RGJXZ+LO1P3X9I8H7ImQQSGM25ydYIBMQbVxA8I4FuWLoj
bJUn7k23vPWSaCHSGz8VAA==
`pragma protect end_protected
