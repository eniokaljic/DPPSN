// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:35 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fKbtCT+AYf0nxp0cbj1OMxhT2c/SAbh8mUrq/vCgF0r52UJZHK75u2+ReKaM74x7
dQmieBJK5TZ9v8FAuFoZw+37k8QrADyco1mVz5U/Om8wIAYKUmMhPylJRd6xqDph
R5IKFGD5BkakL3DkobQobENneVM1RVF0YYxg6FyJ0Ik=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 135008)
FD4IRHkNoVkd7fwD/aFjCJEOoYAtV9L9jtQc9W4wVMSLssxNRDpcWjtoHDTP3HqA
dVI4zMnEczFgryN3qvOU292bLef/qIKklEXtb1O4IPAmRqWu805r1S5xGp9r5hlY
bUtXxJxZ1Cg1bFydzSVZjMixINGtfIorVJP3aovjMkzvTO6FczwoRWoJG+/9zvgZ
/3Nv1LWWUExHXzbyO23C0Mmuor4E/+4RMNAK85qCu83WGw2lY395k9f8jLwY700+
btlHVS3nFEIDUlXkxAcqcHMPSeH1fgjJaJ4ecOTri/Jm5gsZBX+czXLof3hn9mkI
RACIumwjPNBiGkOSHMjJy/rTsK4g0f6GjLDUHmoCSKwWAu1iDaQGdk5QCS8r3wNu
5DBxBKw0Wf/ojDgUjqHJ5O9OUvdZvx5frlN2BF4rh1RuVeuCmMQISAliEfhdCs0B
8FxuBVCEYHpmT8a3kpl6Bm1KR7y2NLSgb1pZHiEaH2oDdfbhnP43pBz6MF1Po5h/
r1SeWNJk+fIM1am+QqjsoHesdrcYLqkip0Gevo7KskZXaizlbs2mhtuJ0WdQ5a4g
Tx55daU95iO3FrZFH1EBxAHVSgXqCdL4fdq6VCQHFgqxZo0FqAwiua1jUnvz0JEe
4N4FXNtRH1H1aQvvS/P26DhPFWSiz5M1fJLOgTYLbBkWY/thLSu7WAHmO2AuUK9S
yPT8v2yDwz3mSTdg2uZvbaG3pZuKSgVeLti9CU2iDV/WNoNrfTubdfma9pogzWBK
2u6oPkLAKTVH5xxd4Xjv1JUp62aiR5A/aw0ng5dGX8Sd6ZTMxl9ThuEr2GZOYJx+
khD+pPSxFfiGEKQEHh1ydUNuW7EuM2zQNB34yIq0e3oTDfAMRIRVj5kw01Cwv8VR
1uWtioYjvMDvx0hMItJY5IONkIklmIEurdMN2oibgYmFwhUDp8aRhfuMkv0Z1ZWT
zDssuvweLgoolBOTNKKcJ4bmOfebPDSfEtQSxfEyVQfoE5CIgD5ypGfQTyKrjyUF
lIY3iiu69tRMl4lL1RSkQCvpgZQuFGq3f+hhcHa7Gg/CIOF8jzM4eqVrwmstwHWY
RvoyWbOcODcOHkNKhWu/b9901O6SBWS7bFNyZauUYo7r0daeRyDZDg+OGg84/HEI
5Myqjw9+jKo18mSC6eF/CR+pWs4He+AhwkQLMCZVvy8COPTZi7WmQHRndCURxbJY
yb+5iiqbL5AIXrTMecAzscGhKlAMtNBfqU2JEp+SxcZJSILEwrTUzFM5XUikeRki
mvaIawC41P6ACQDdlqsjEoFNnNvo2q2VjYegZDXUFM7Dap/kqZLlJfg2+9xQuvXe
JZZQEnVT+zK441Vy1f7XosxgA4X6/xAR0GZKJpKupRxIvoKztUvJiT60FvbgtulP
XmkpEJxya6GMADfutaQuto+lrmWmBGKwe+vLTt6BYPVXneOcoQUR4mm8ZVSU5XC4
H/F2fMjg4kjlQ+68NFIX80Wobk3PQwvKI0hyNW/WAZlUzK6YcQ3dhZllcywzbQ7Q
qWLEBoqqZNubOVPUquOeu6NnkkvW6rS39OAZ5vfD/o65bnAtdN5xxYQLneQ9D8Fi
U3hEQ+lDjIJJTvI5aaUdnsK3kbzdctiHbhIs+Zykbxgq+qs2xmpArlhZbYkeQrfM
/848PzH/rrGoPP4tK/2Yx9OOqD/+qgqiyDh674cnjPxGCQSHAdox5C3Qh70zMSyl
TWwEpaLYCsCE+2WQ3Zwho+AS8oVax8SumGQ0rocWCWOeTW4Ydcumkrspp2sxtF62
S2Hk1gylE5qpEmQGiZMwfH1e99DCrU5xvXzabZuMQbaujROlNPzosEjxqA/vRrlY
vEhnQgguDCoSupA9gGSA/a4Av94tnBPwOPaC6ZSzS2+QEJyhIK/wgvZibjTi4cXh
ddwGdpefu/kURSpcIDBQfn8lSTJ5woDtzk5nX6pkdEpeQ1Z2yFbxRegHC5eH4D18
lvyotWsKXaLaK42BCGfpmlam4nBvz6YFoRxAHoezhgsIVgzf23a2X5xz47HDQmKU
Hup7Q/MAXOy8wKurpOiPp7IySE+gECOu4X6lTHrmtlOWxchHO15NJHaqHLp8rTjE
nmLWLRuc7pYFcXS8PfPCRXilq4Ps7+mFr25YXdI/DpAnOpNqojU04VqKj5YIrGsy
8WOyKO/j1iKR9gy0fxFxBqBspa7NvV6VZ7SPQ92y3a0iIZ7ctsly/+69uoco1wix
+niW1uQtnIh2/kJdKGpXYZa3M1WOhqa/hHQBrZDgIxd68mdvp2pDIXKNFtMW+Klx
Bgqbr4ddmt7rCYYBwwws7nx/0qCEIxVnzJF2g4aUqo2xYZ36LYxwXHiApa4ZBlnM
chWzB/HZl19FWRD4A4ttr4fhA2CJwQDWQ47rVMGkOiiHItAPBNG7nK5xbsriHS8+
niICcc5ds9TmrAXNwuduvqAm78R1dXQh32qjrftpgpnYBBtYi4reRGTFUvHdqqvA
C8hTzACLoQT2L262LChU2UlENAzUa4SzkyLXe6uAujT581shXs4NoH/TLTuXPkO0
WiBwuADNSYgBdBbj4cwk6vvpwbkI+3tHmqGZ9t4LTsG3sVF5DGr9BsgBGtdoJyQX
Dqu5JSbKnsRQBM1EWc1SjY5u71WSxDlt67rT5gVxh4vLdljE2NnNmtinfiJZVJDL
2PQybs4qU94Q6gQEuaLHisulTBWHbSpRgStqMaw6Mww3phmA9mhe6h0D8AMDQRdQ
kWpFI+8pK+owzyqeZxzpmaiBqyUXZm6gRw6dG6PFjqfLPKiIOzTghQQw548nYd2t
8APgC6Y9mXO6HtDLz7lfRUNR5zeQ3q7XfI5XLWgo2vkpas6IaYB35HZ7wpoQRl5m
DgYC7HPFy/MwmND/y8jpH5d5q+Pum1vCJuvS+YgpWrq4Mv6bcww9Karmkgo95cRn
/pV5n1j6fipv8W6KDTBUdyfdmxrXtEe42XYSP7jHTkyZiKBUKEGp1RyL/WhJOUkS
4g95qrQE1DaZYctWeOQimZyAvgL6vqJXHwQYlZg1Ejk2pHKFHQCJArfKlJJ3FNje
WBOeVu59vZVFOQNQ3SjDusFshzxi9KI+SRfoQEa4Fb5bczAYrClFFum1ZjMhEl/h
EJAKNMiUrCG2mn/sEdMQ1zp1Q/QOLTmbuZpShuEr7dV4Ogyru9quzn5+4TuxN6J5
4KDHLOL3vxEnpRyyc2c6xZy7s5OsB0jscvyduLNl6nfgRxHn/HVHBUlTZ0oh+VWH
NFa6X6Ema/RPosqnFZv6Po6Hmgov4XGt9q/1U+ruqVK1W3aTCmiKjpU/ymBzXf94
vA7mqKnu6LYFxqED1wa+3ej5ySL0TxDP05wpl9xvsRL7+nj1eKdvVppEhPISFtQk
b9ydtz3YQooBrfMHjx6c3T5vubuz8vFKV9tJicN8nx48N1e71NafNVQjcHXhpgoa
LON4B/X5FEhVuqWheZWO6IpoA+9MUlz2tFCYENO5JcNVUmF9VfbHi3ca1IyNSdsg
0wGDXAitEEVdu9/EAz3FVLuABTcyVUM1Tswj69fEqow2p2TwJsKN8qb2ADXQGguf
B/HeBeSvf0zAltuzWSqdfV0GahPcctggSXnXt0Q8zHEYpe9ydwGAs0XiFt5ep2g5
zoICZU04DPlDvJhXLuD7sMavfLenkt6va6duukM49JbKR3Cuta4DGqcnE9w4S1Ll
FJ4UE7TbJD+r/Sypm8EpO+gBiKA0o7EvOj101sh6LGg1JI5LjwEy5Z1/zHZb+osX
+oo6uqIYLJlXBp/gPeIoM2tQK57nHiQUf15/p7TfRkQp3uy17/+XQgw+gmGqAl7D
QCiHpoKebskSZwiJHcRLK1w3vZztcLs1rfRfULwAjNTnyI9s31GJtqfGjAxx0b1/
wbXm4oPKlLzzWbVjXvd24NT1DRB7r2IuLChdRs2Cu/c2MkRW3qzPP1OiW697nAuD
29qZCIAMv+eCXbUNv6UR/KY4mtyFSfoQyhCfxpp0+fZA3xc+WJSyjE7Rm4DgSGoe
XyCs22zGmYe6di424zkfO3a+3sEy/RXFK6KOZQRai8ulHyvOeDI+w6BRFGDf5orW
IQvXyXHDI/5m7tZ/4wHQIayiATu67UP0Ms74jZioRk+RAIp3geW1wUKMPS2BXGbs
AaaXGflvs9YWq89i3JSDH8cHKKPv8PsChzvFxvGWJsuJOu901xVd+p9pJTHc9dVg
JSE/yWlaq+GW1EDXOLTCmKty9SwZJz+FoOp5q1CIdNccZ1e4dvoADB417z13lJ+H
4Vkiy5/oaS0Y8m+Fubs4EIRdtUW7zLUte2NysD4zpzH6zTpp475Cez4RnJDVTB4S
p6wMkFS9+sLC/EiqfSjPKNln5IhEu9vK9HWPeoK5N3mJqQqFUdMY7tgbTegrVtcS
NGXk15esnrBj8Feebg0CDbG+gE1Beq50ucVEGP+j+WufBsNDk+xqaYe/Ls7lUNIK
LTt96ZMoy1O6KTRq/S3yG+jA08W56HQjfjUdOLt419n0nelBARlj2x65C+ncueB7
Bs7ofBOFdqYgTLKrLP+cwDkl81gQomamtJJwB7gDIqQ4MkvV/qWW62NFRYnWEn2h
+efq1MlbaLke9VebUZzzORI0Tuq29jAssWGuZa862QL1dvjwqVcSItrMrdyIJweN
XwkHLr8t95hxRYvpr5+O+/h8+4G2Xgi6PnxTbaMF3xnxRhSyOseCKGxP9uPZvD3i
iSJSj4BkLZGAuzkVIOPrF9+f+5o69XALELumJ89OV6O+NmBeOlE7i4OeM550Ni2r
qBDFUnyHa5jIjDtVXMt+XxVNLfnHPUp3V+0yeFC2gmtXwPRBalCnjzzGESlkQ5f4
dKyeGbym5HpcKF/08U85huPoc8+Xsv9WPfbBV/pBsex4yMeJBC4LepXSACSEyeyW
Y+2dZFAludbrXzyt8o+k2aJcN09D1l1aoO+hTSzpUF5slqXoVJcc/g0fbjRnMsmf
+tv+2XCUZY6bJH5uIxwVbr1LDt6zlexyqqIuh/AetLcoMTrL2ciP9XZFQgetJyz2
EzqVBklUf7fgbLPVlvNles9fH5A8MrVIl+zwKuDvSC9kn4x3F26h4OOWQoIbqZWX
ZX2jcGFBWlb2apoeFBS0c2TdO8/wjW7LcNlLdBkxleW6qwX2SKX7YCdezsHkKOzR
g/Led1iZor7ZpGptDoPL8wZWda6rdlBVlj2nJmdGjPquYZoGvv+e9SeDQLD5zjp4
EwcxfX17dOcxU3EmNKUVORAqZ5ArDlqyAtaCMXiuyFlPXOeDESrSkThyCKtcPRPM
BCEy2UC81J7NdVuC3kcee2vnwOMjpH6dzl+hOrWSJ32zGDQ8VlImG2+khBHICA64
IKifiE4CTdoTyYUsicjw0PIOm1XoH4h9Z4W4tSiAHdLooOiq8DhSYU3K3r/TRhv5
p3isTkRfXF90igd/lQhsqxRTtNnFGFkay2ZlBXVTwW73h/vGM4HCDTmPS0IhGORX
LpZexxFY9Mb2GyktntkAxdjaVHIuBxl3UvrQGPwWgEwhJc+dtMupUDg0u1JdtD2R
xe4vB+DUz0wazeaZ/mqFaYHwKETXhjP9p8i4npa5gE+bu1uCL4/o4u8VHYcnK7sC
jH8wRfOtznoGk2wmj4y+31VmqhjZ7hxISIm7CDHKpV2Q6GxZyw+feP8P3HduAdhc
YW0S1VQOlpxo1eD5VVQMoJQFddrpJewfRxXOQILuwiRT+LL5UDKWFPnIRHdvcCrx
aHjxc/M5BoXTruZ51i9M0ZdrasJPtitniuI3Z9ZxJEzsXe5tg4XThwtANTt6WTp2
TnmBW1pRvAAqITT0WJba67Q8nmWgXbX2LXRdKZMJemW2Z2JOxLrn9xwKJ8jCsUvM
gaomLw2QBnXA716FxTxceUxv9c2ZTtXqVoRYTLnXMsnRquE8R7x3m50ceNZG3eYw
nIIeuT+FDR9jtkTfoPZistAda3XY+rlD9lYk2DUxahrcRPdj0+8L+MHrjqYpLA96
lJA8gbSXYnf8i4IQtPbP+aZd0IypzeQHQQ2HsF8C2c8NWja4IzklCtxny3Xpiins
sspLLz9Omwl9CjhFt7zzZ5PYgDhZ6dD+0mMsvrkkqiXmIAb6wTgKuvrB7MbjIU97
2OurTwFHZnfUuBJR7aPSpJqDqoJkn1uscZ8A9tEJbNJtArZpE8/MOoFAYiSeY2q0
bqKtphrpl8o59el0jxZZgCjpxmYMQPihh0KP9MNTsT64ObsbYPCcPFr+Cc95hobF
tqseH5t4+pDZV6q2m7Wgam0U7/OHeMXkaONQ8R5gOvfDYzrRK74n+oKm4psW1+We
axsH/5x+gbcZ37JaRvXGWsTYV2OdzQLM01ayGxH5elV46ZsKard3ullQp9Hrs16W
tbMgQbI8os5KexQKRlFuWw9szZn25gLzHl57TcvQdwRqgyGwSkbz4Aa+9pOSG+S4
GZwZkeeMMUupxaKhcPNEhEALlKF68Acv9irJXN2giyC1lq9yPmXMvVFmHnytNeiM
9mH3i43libB5rRqTZBhIJ/+oiH5/ovLccAF2hE/gC2Wr4wmvh3/fHCLxWdCOK+I+
qs9DhmxYoTEBce8qboHaJ106H60Tt7j6L9C/YO3WMgejrc4W0z8GkhfXJQaNdGyd
AcCS1vcx7lrhS5YRK/48265kd/GznWpFDHcbyGN74ZuQ6ui6z2brMOLScxLuIUmm
Km27AoTZ60W0rl28r2kUg1f8/TPJT5Tr41zzNwR3egDiB0ErK8juz9+1xWgkjopo
uc7N+ueyy3yfaJEd/YE/Etb+eS+6tlOLmFPB0Z/SSgAIt+tqgw5b8RLTg67kSUB5
J4gQ8BJxtd3ix7HpferLaW1dx7sUVBxkw65aI+nFxC0CM+UXxqKXeixgpeM9yaYs
iO+8YuLOsHuYo7iUTG6LRpP4AzhwIqGC0v5DU4PR7iKMflNr25GAK0IVwRijRLYx
8f1DBtSAMtUNwoAgtcdEJqpiJLBxnod91fLgT5OJ5GUH4Ipz0VMpESzolZncj5nE
bxScB2TkuM/89p9xZKOz3xck5hC/yTGNFoaAoxygwrwnoAAdXfQF/tSG41Keht7j
Vphph+NNHz7e2gdNRZjZE2KQmO2LvxL241hLVuNgq4oxpEH76mF5mwLriziekNBL
RlfHYzvWEXtiCQrVrBxqu3uNRPtkI9ZdFSdwDrV1j8g94Ube4Ged21RdodWFY6KA
dC2/famQXIo7Ps3VUWJwFOyEpGKNWh1TMeckWkzt0cYkSgL0KXPhqlIT8lLRxG7O
klJJDqZsF/Yvvy2FGPOG7or7CYvzTTfFFNisp9x84j1P32xSQTFXj6rGaad8tFsg
Kcl26vq6iQo8wo+jxKoCELXc4x2zagaJOeFK58f4cFcDITV45iQivxCw+jdpwdEQ
K6fQbC2vytNfLN23r7luD82oegnMwtLGv2zO6+zTb+mK5TglxdfyaDie01XrD2K5
AHyk9w4/6JYszq+krbKUZ5UrfajJzoPUTdBa/UfwMd05Casm8t4PV2vFyjIoaBqj
IOyS6A+k9vk8V8MW4ZhqdnAWyU9fOoPWoOqK1tiH2j/Uc5i5UQuwTFT25gxJgxFN
Mtk8BxPTsubRz1iklGWsUZxgvzzvbVidSIdXe+/FaM0e/xaYd2dIWlkorctPUxIm
pnYqJVUHwz2ytZ3ctI/UBMNr3bmXQt0FzG3gAzKxkLGSoQs0nYjc7nLDKUaoLNXc
zJn51R3mQpsa8E1v5/5WMuBC45lyGIqdWt8lXbAeVmbeU5KhM3P9n3yYEXvKASZD
chwhWeR0ryLH3IIgiBseNRJLiY+/a6Iy6pP2RqrsNPsl9gJavNisxQ39pEZA/yCK
M8TWmFYvup3oCVX1uiFClHPC8wgb/YPnCiRtyNFVRbzl9+SkGNGmFQ0g+6AOnjd9
oxFn1xnIl0d4JUGA+0M1RmJES7q3uUTny43H+ctsuQTlDaOcz0scD+x/ZPcf2RC+
EwxGF9pfehTx1gj2wqq/nI32BnX9bwLmLtRUSgygzNyQqT8Q/3yqe3bvnEPhpRP+
7uw3cONc4ykv9jlspJGtGmGn7eoe70AaAybrMo9nSZ4K+dDxVk0v55SuZqHwBZQv
DZBJIdpm3nS1mX0d733rn60I8b902Pq8g0nzFcmxfaplzGn9ZhJ/XCEAV56v2ZgD
0fDAJKkete7RJ+VBSGx3qvF5tn6GLARKSwxUufqyTCk0M5UXF9FZRTIF06fIXSVZ
zja8LUc0+HGYYxnVlaz4nrUcuqxdONS89Myo61+K8PD395TqPz1qi26EJfybrdDz
Nq3k1f0ZiLZ2oZrQ6LPygiJLkKRpqpHkyvh2xQor/KYOYgVngkSWZLGNO2apwMRS
7lBJFoyDt3bqy2TiR3f0DqH4gL4hJGubjtdU5BPfm4pR+fahGYqFyzNetPgSIQER
tGWQeUhwivtSnCpst79wLif+mzYzX/qXzovvmgx8/unXCIaXatB59pgqy+S7BCwN
w/LKRkXI4P6jIDE8zS+9T9WIrUuhxGN4aJts+XLgExLQp3vmdnMwWCPcgaZan9TD
oBpAGBOT2oeyJJICyRxbHm562MnXVTObNuoGYYKvzJXmhVtMv7Ubwx7+DlebIXGn
gUu6mDssaDn3BfGLsIiBEKQW6a+48RKXfFXYan3spA69AkGSV2xkNAeXzipzhequ
nUVN5agmmQ91ePg2LHweBW9mlTeTkUDrpIncZp1FTf1Nw0ZFVwAOdRZACn1IaPKe
Q4yg0nxndegfv8bsSisWy9FCjvq6WGsEVXp9MuqcMsN8M+HHknbeX+SZWcg6u5sI
IL/miwLzrZjOSGyei7BzhdtfIiM0D/PAqFR2RQVcYH4Hnca9dLmBEcUceeNo0esA
NmtSDVqGcx4CUynIqI/IeQb5mz42DUm5QEA+UCmtlFkpalDcgBKND01Sfh8qUSPV
iXMluLdiiYljudXDVb0UDpr9d6Zz/78+gXGTo3yy99HDiMgUj8zMD1LVTzHS4dAt
c4r2MPHtanLg7LhIPD70XDwpVZzj6Euvc56G9me7tc1fiKcrhQo2G4A1t7ZXle5g
0CA7/6KDGlPdkbWOtH++zDGiP4iKWn1v+1Q+MQxby5I32eCDp9f+1u8/HIV/oH6n
as2QPWEfwkCtA2os5G8HVWIkpI4ORyn5qHdrHy38JP/TlzyjqFN56Q42cKS93EZE
tqkSfIb1iNWDgOvbsFlvgDtp6G3xaxqdP3iCXpEDR8+aDLmVTaS5iIihxy0VRRg+
eq0aGuMXkkBxwXc+K91R6fVTNppYds8Trzc9Q3uXu1U2eFIukgw2zUAZZsN/4hNm
TcXDeGhpNMDIwmN6CxmEA/2gYGfBUzo3QD0nQyiAdGsq4GnsrU1TSs/QRdSRvOIw
rR0Krsy2JPZPrs9KFlcye/U51sBnRNxL7S/AhB8IIK2KSpk8Yq4/voIe7o06tjN1
0nJ2DLzM+SPowbD0WvOxqgOA2fMj8CNtuYg35DOnK50+0ZStI8HLeuPY+IMJOc98
uUA7PHj6eA/sbgj7dNI7lb/Cev/IBAIa816Wui8coX7nF+yE2pKlak2QlMWmoaCi
MGzuneVvrCzg1Vy9UHXy5dNO2lBdc19pSKxD1jxwF4+g6Azak0SDg3+R+TepMPQB
JdJs7HssBmwyaZt2oOmPJFZuXiGLIYoDfXtzrY8flRC141B+xUC4ZrOcmM9Gmekq
ANE/xYsjyazIJRhu1tYgf9xKeQQLEyXFUpx4todu48fmKMpYP+pn56OVrLmpLxXt
Ode0YyNQNuWh2Aw8+D46auLG7b7hqcKUCJdoxOZQ7JiSJpxXeLTIAqc4SspFYnAm
+bJlzme4oyUy33CWYBAxFDgrtc/Sa6H9wIzokoZ9SbDJEdJfIoHjNZOjzh2TSI82
dZHBKBxLBmNAxy04uqBa8Wn9t/8trxNCxE7krsFo+AmFILBlyWCwCTnfdziLT/5w
AeUn+i6SqBkkVJZldB81TY99SrHOLfa7IJRfwIeBTjVsEO24sJAASRN/7wkSV0JM
NnS/sheiLUIJresTiMvnWf1L44mCWHEDM/J35sVUXT5tSmQiAF2dnRGHgXUUazGR
w/yC8M6Nu6LooRnwGnimkZI8koHtbjcPxjhlaYyltKMIU2RbDw1UAmcxeRSrWPU3
HfYC8w1LkdFC2evrkNbfw4J1dwK1qnlnU7/O2eEBEapWBpwO3BomG6O24L9GRck+
+2GhdUoiqV3o//A9dd6Ys3DQ0enfdZzU//iGm1TJDeJDo5Qu0ip32InhN4eHs6p9
mO8WMcSx4mxsQcFeYzys+Rrnlhvp9RsQHi202/bZyj3nH0TpOBzcryX77v8U0Ir6
kHE/VulS/zaN/sTySRrHWlOgw1iGYP4xz4F1U4oxYnuzNc1ubbxFQEdJH5X2uO2P
BXZSm23Yd3tgOrBBjUApDGFtPR3m+0TrnNLu+jSQFh1xtMSXWb6vGiQU1yDxgT0G
Ax6mfrgnG3HAskYHqeNKXPq3Eb2WuQEFfd1OpfUs2CJ+kcVIiZJJxylfyA9MLI0b
xFi9JsCa3iqNPqat4k5sKIIF0gcJDexdA/gds+d/XbLdVNsQAaePI8xmeXRkokae
DuApIYRShC5I6faOUoTvsDKt0VSlX1hex4ELCKC9F7IiKcHTFodms3EmDcKSRFkS
alw1kUgFs9cBxOjWujkCaiJWOMyb2yund/bl2CYjdPPqR7tCE0loQ4Wg3zJAWKVf
i3fCFdoRM7BDjR8lZ4+38qntk4Fr1kSOyS06b8lnS2RQx3WhygkLPCl2lFvJxsTs
OFCLWBMoq2wQy4XdxnKq9pp0BBFyPqqOyS3ke7LqGFc/I9GZpHmGRjKZpUyIgX+U
xBq3BhTZh7aQZE63kyTiOMBi8KuvUoV5G/cKmagg537iKn/DvjWaNJxpZJ3WQn/e
RIfsoR0sk9J+Br2dqHwrISQoWPl71TIQeDbPi25HANKb6uAWfq3ap2vZfisAOpjN
28MwIS+9oGVVrOzBF5Uml1+cbEM6T66Rg9dYnh1iRGEDzEAPc/Xe1bkuUYxneHsX
23MYazoMRtc2yMOllHRn4tvSMO9QLCd64Py0gEg/BUSZuOtK1tZA0BTR2PWg9IaM
aCXfn09bopbRjmzUiAEg1ezf+MTJ3xdcXEJHlO6qBekS6p5vb4D7me7HFwgRW/dj
wcqqs23U0jc/wnuesBCZHeNsyAHl256u003BWIYJyji6qEElFGMaAlWVJx0EdJhd
sxs5g3WOcLVaXU/imz80JjNAIP9pi0ltD/J/QHXuPSisi7IPQdT7GxdUPqKXDju1
n1/zzb15YB/PbRsF4tbPwAZeKJQX1VKZwCDFHJtZL8pUHAzOJsrhpzax/AS+Dbxc
OHk7jA0jQFj/ooeWuXsYehbc7yXuth5ycSF780gNURXG98dBoSHFwX9ElqPvEFWH
WfoPvyNY4pz22ydVwFTVtvhpCnJMUdNzmk2110h5eSevfBPicLT8N8BMF0JwvStj
at9+b2wS9ahyLAALE1TqVpij9x/RsHjTqFjEFf21sPBIJtyIatIqJyr1L7RbJ8XQ
YW4MvgtT1K7zL8ejkj+FgMMQ/JM7DqFNhTl0DdSbp4c1E6kQNQ8TCZpIHiJSzv7h
LnGznSyhSIyx5cqEjBifzHubYcxB0EiMJDmLkAfKeT2xuuZ55clCGwnTPk6zKz29
N4R7rTLxD9BUivsd8wKs1N+stvTX3WlmPzlIwrvbOA/bxxLPLVG7XeP3qVLK8khT
klLFpAtN04Ym/FOqI/Xpel2djqENQ+oRqans6t28fGTEgpZbvKCSdGBfvuraHd/7
l/6MlQmpnK1Zl+5bVU/21ubC8Enm7JQgmXV7sPUFdzUh2eGyiOFCAMWVFPYbzvGo
tNiDQr2RWXbZ+PnOKlHfhcyoM+x3VANzYfO9J5m8ukvMBehu3IoMatIu13KlWhMC
gBj/D5kpdzqXqLDBUNZMy6mDKFhR/IakA3XZtsOLJFWftel67rMYEIaJG+KbK2RD
4WS7sd5+m0vFzNMJsEb8zc+PUqx8UWqqfsMv6UEypFRXHgv4ZXgGu5/cHwmz1Oam
9etnKRJpny3Ri+obiAlacrxk48AbkAId+R8Z9TgbpImNG2wWCPKyPHon1NKQBuzG
9D4QFu6GwOPH0mTtBZgAKvIndP8Yse64E1/N4Esce1QJH4cD10s1Qb4ZAFMPd164
TXWmrLksyN8u3k+zDATPOtj4fTMQyqDs+cQDJTpyi/Nv0dfZq7Eg5HGfgCVrNEBy
P5S5SMMSYlq88pzehRtIQaYsvys+4jXYyT13V2Dw/VXk80SwlrntT4yVcYVBwwxJ
/M4Jbn/X8z9wHQ3D8572KynHcJg7OfgWgsb59Cq9xPDGLKYcsDAml/fTKw6+o5fp
zlBypclU2sHMt3UodE9qREGciGfRspKug4/GOd2rjd+h0CD5KlVAKv77okDMFV2z
9pkhncgXlCxdukAaL34KGRdSj2F5m1ejrpWwDHzPyskaMwM9QtP/mBiIlA35WSrs
7ySmycEpOtg+6oLmJtXfPN3ChndCQ4FMd9nEXxdPMCXfctym5Ycq1TznSibDJiPk
fp7X8ElLahYGigJInK7wpzMHijUmKnBx/ILZIEZ2q5582t7J0PQOTGNXCL3vs5zx
2C1USQxIHw7JkxlNMX+OAq9DCF/jSgxDekoHfqrrC56wrh7ZCddMGBI3WzElPIr9
UaWdPq6h/TiReqFlO68KlRPN2+a/zp5XtbG2MMsKIq5Q3AeYBVVAButN00l+g3ZB
VL0HjrlXNHJHurN6R9CGiYMBje10Pd2lYLXqaLTgR7vQ9lJ2hBO3O28aEgdnHPeb
BHruY1sYYIMgxQJf3tBBD+u6bTrRrOWFAd0GpSZU3lkfOxMHAFkhT4v89hox/Ie0
tZgaytNsMrSgj8X6FVaEtVz4x3Yj2fkJgU+FBiZbaa/0bznf8Mxedeye7BOShS+z
roMNSfFEZwH/uU06WaDEsNCYpNzca9ahj5tj9GYaVlYLnthJEHIX2Vs7gu8bvkVX
nRkPxWozh4nPSST+pMgsBf4WpL0IZgWs4EOchHrU0q+/0Bb2kLufwFcIsmUq5GbL
4RmFHa/z/H+vPIPJnqQTE37Q+fjjK68H/zR3Ll4oAR/ILkPyJZQv2Zf4qFr9uHVT
EXSzZsDDTRgtkFtA7vfvBjWfsyrJFAuL3gzDND1gf0O92y+kplsRNidPKFv9pXBj
UTFn9KjLHabuSM63DpttX7XRWGvum9wxxMrafu+9ogN9Ny+fN1atMId3sSvdzLvX
rBEhpylHzMuPCRcMczdRVr3C8z9RP7yafhjT4qxTb6nzrQynuRjNR+hHDRJ2Bla1
JN2feVCNZNODVG1/ehg3el/86emKo0YW2iPpNcfNvjxBUpgGzo27ysbaFv2qT1hs
KGtcxaC6Vhc3BkrbTvvkS/zAmvJ988XpppBsty0+eYviupU0PXPkYhOUVyDR8f9m
voyREmvmLwTDh3eXP6871Wl5PqYx/v8S7hbKebyV0pvk9sqUk4KgJcRbqKHxBau+
OgxgeIpXlhlvLGbOeQnPfAzFg/LP7udsV8gnfSd34EljiOUDG1XoRoO0PptQRim0
7E0uqxtPsXqZovNL03NVVBQqrtXwI4WmgY/LKCzOzse8qQD4Io6lZiy50F6y2gyD
z2g2n4NjQn9H13zzyG3M7keVS/8ILJKhWrLmzKmGxZEIfWk+YIifoNDVTjWXXl5K
moDqXMnkr5bh9jNYAQI3yqsa40xpoIJOzVQU6FOJ6NiqX/aE4vYzEmTdmA/NJ3Db
R+9glWl8xmLd98q1cOwyu8ozQHXKSQu0cCR4IJg8DlTMD9VLp+P9XQdXOYeLA91r
NxDf02Bl7LqnrzkVujJaV4SrZMv26Us+60ZksBZB4rG/L1ypUMWJ6uCqxczi15X5
d/lvU5bUgHwUnOPaLLaGHnXxOa01cO9HzRdp9YjghW0KqgY7V71/Uh/Xx4ar0xyl
DSGD2VF2IbmIJON5AmjJHwARz0UKOBOQdpXU3KVTsQJvfxmlZUHcsOdWhkJnT0x8
LLt5rXB5g3XiWyap3lXeXqkRXHlo1vaqL2LT6oMTlqxfi7c/Rx5pkrgZcyA6c2/X
SabEKISeht6DsQ/0tuegYUXlZxZUH3/b/fuhyEhpo1uf6O/sB2o573v7QmZti8sa
SKRkFaag6MOOEMPoTyoXSEBqk8NeHJ2452+Yv+dIhR6QJR93q3GVUN0JQtGzVv/f
twH+VG4J/fAgFeHs9hnW+JaH9PDLywm0KxP1y9gfbnaXKtlqJsYg8m0nPIMnD7Mu
F1afcijCjW97GIb2lnaOXpZp6y39eZayuNGrU86C17o9l2BEvtxVTmq31qLMIFKK
OsuCaXI2cBe4p+Zjcecg+9uO0NmoZkLrjHWADu0/YjdiJ0SEdg6EmkLe61b0N1wS
Cm3QRrWTWz6YX/a4qfeqbsbcOGq3RZfd+1gMDM0GYaZ21mqqX4q0bkEZy+IatomU
RzMzUd+ZThobqevL1IqJ5FzMoORl13aqU8bYLlsDdknT4YMiptA2qeymRtFy0ms+
OFe0lk0sntnBu/ST4P91eIrX2FyT4c/1oVAjKL4TdTjBUj8Qt4jMgjd53sZd2XtN
qpNebXvlvrflx+3hYXl3RvmDdy0Pe/j9rMJMy8x3mdVN0l/+ERFYKG9lGndmZEDn
B27I3VPoIsDY4rRdZOxARyLOO5ZfSeeVpZL+yDd8VN7sQrZBwAQ/A5E4qOKH+a3g
Bi9p5ET1lAOtGr+7Sl6FHalcvRBwU8n0ke4hb+ArUIF8STSbbBtBKchjHR7qIIMx
jpIKIaEHu7Z0OBRTERUsszaLKevNBEu6tf5uGWm40M6EzoRfZnWrZa4mFxwAhHgn
55gJy22yDSer/Qz8Gxo057oDgRdp68s60azxOCTihTKqz4pVjSrl/K3J1ASfxgL/
kzwPGWYHau9LtO1E8tRTxg+G79+gKItHum89pfIJvf+OHmJbqfAOz9tL72DYendX
SO12QvqJAMlsOi33w43xZj2dIrHac4l3Bv6QT6eu17FvEtYPrwfluVebt9kdvUr4
V7UMVt49z3A6vSy9yuBVXrcYCqCFsvJzz7gxiP0M8H3rkZeYbjnGYhLatZLbm1A5
OcnIGz6aiDF5xK26r1WKUVqMgzIzj4cd3Vb95PM80dLDOrQy6rvD+IP6ivnIftmb
PZCKB8CKpSMXFi6aOEyI/A9prFTQaUmvPyvMFWhvxsMlQu6s/KviA6WFinVT8XJO
x5C6RW8jzJKnlUTf6mANqCKtQu4Frc9Y9o/QW1j2kXP9TGL2qURBHUVzwNagZVY4
OB5ocUWhGetJambpQe08Duo31SxFPAEDBuZYYIh2L941F4vf/hDfGbd6mR2LqO4U
BDyIDjKWpN290VfkfqViN1U4KycmkaKObrwApQOr2RHM0tbomkA5KrW9/P2zfy8k
XN6becOaRiYWegve1VJTZVd6QSCrTnH3NfvQaysd2VBgL9Et+GDSfjJhmqC9o3Nu
njHFufWqPakZPOAvIH5dbuKh2QPwgJIK5qfIC7cbyyl+/A7kCp/tYOCoFXxNkrSE
0k/L3DlqTRv9orwz0LFAPImcdghGDNBBmSHpum+DrBHeDkk4iJvBc+lTq5Y7Gk86
ONBfuZGlasQj3NWm82cwZUy/MIrq+SlGgyAeJagMh+4l+DoauZamp3TmLMcHjW2A
rVcpzFvZwUrDGdl6T19nqL6JAQVne/ranJkF1DCXfirsmI0O4J+Ben6QuOsWUc8G
tNdDT3oKvu46Wf1ymVzwcdcBwZXbsIug5D/+AGmXmANymi9280qcuh8uvgCjzI8s
BpwAR0jBIfY/M+oylWoLwnrxEHngadbGELfjSqwy3iZ64bU09RXIjgKrEsBhD2/B
MOclo+KypzZYYyWROoVVFKEDhLET9oxH+J7TvndouDA/HVIVvwt2klkgpOAbsLal
OTJYcQnl0rB2iK/XB0KupJGCn/bBf9QMm4hHDjbP3zukKX7AZnqZFUcpT9e/fgTQ
WGbRN5EDG7t1VC0tnvLpj/qFi8tCE39+khfa7REhj/psKzjpdZbQFZ5Zrbmjiffv
zqcdubb9dwnvoBfFjDWmQwKgAVGpZPfeiyHOmDo7dpkk0O+FfL7NANdJhz5xaB0B
3YKjFF4Yzr+WJivm37LivWM84g2NAg54G/e9WrGVi3G9CVDwG3Uhra2NggHRlVcO
XOzyZcQZFti00eCK421wy+K+9O7gq61T9le5UuNqgdmQpep9k/jP5svT0Ej8sV9g
6SCVzVZXXhE0VC4v4mE2oU+vhjo8mrmctMd/c9MG6C/eHkLNUbxxKxqTfJnybhSW
qaEwutZtlVh5D47qqqzNo/xAerL3buPlT4GiJvUwuZCoiCYlIOHz0nH+j3xPQ87u
6ZyGRV0Vz7hg4hvVWp69bgwUw7LqLTHozv6tD0YHb67bokxcWB+EO+mMnliKjqCz
B2Gy+XPgKmTyDz4/ZUTihM8fhS7opTvRw11BhJqBmmLXrUXvizSgsqhJipA7Xq5/
qOuk5NExECtx7mEoQwUs4YVPzWEXewLJJB9H1b+JUh1XGnVaiCCnlE06gKAEaZKF
GeQTS5mHM+XHc5EAd/3PUmoPEr1n30W9AvfC0ePuLuqVginPsskNIGVTRZt/S9Zh
lBPT2YtF8iaVmTpMtI1R44pP9gbsV3BUgub9ddBXy44peJ+IgDBSIUWTPx2Wdj1U
byQECqUPrFgPZZm/6iRayD0xbQx/xaijS83xQNjr0+t1zs9Hcco93euwpyfIckFV
ra1QfafxpU56MCe278EIXl8cmPNREBueIjQTNDKCpPP1MPZZDSl40xOIdrK1ENm0
IqFQlldaki3y0dnQl1MhaE753eSv6jO9TK7d3SLJIQagsMq5o7RMa8xkIYPiuTed
PafQVFSk+YAL5XmQdC2sfuuxStx/wazo7CLxXq8mMM2PwDuGcOJ2tWQ7PPz1PILY
hCNNw389LEDITpyC0QKrmr1mKVfq/p3pto7HLOoKA0iyEfQ+PejjrbEFcusXXh90
CsVPPLCv2tk2pQHCyV5T1QrnMVeaDaTOhqZirOy69Sn4AjiERh+AzCx10xmWlJWK
y3U/WmeJssaCTTgdha5I7E9u6k9YzXGWcIBkGiJpk5GSS381dieETMiY9uIf0AtS
3WtC/xfHJnP67ONbzcEB4jYY1YoKudneyo0DLEm1wRnBH4BbEjMAZWHzLW/oHD+C
2+hmqqQj7wbTICK5sMokRaXp7zC4HUU5Iq+KRCh56wHoizt2phCijpue1pBt2H57
FypsPzdWDSVCf+swkEkg8CRwyCNHSDEk6ci87BRP2SV39xhoE+DYK1mUGLEiJ1P1
O9RlENv8FA36J0+Vo56lpa/dzFK17h0U4aorzDmLyH9r2hcUKibdWjWQ3ZEG46al
1s5B0ZaLdMamn2Ys2L0HDCEBX2R0+gWIxoTmpEbvxbYb834SaIT/eOt8wwwfnyYo
3kjaUcYSZiQRtgRwrMd4NTzWgU0cRpWuJ7aTpFmRNRBlFhAsIzGNHUteQrpV5DWU
1B7EwthTRHsto8X9DMW6rLEbX1+TQicR5pgU0YzDcPAEbS/ORWxlgSpL8sqhh26N
EMGNx0lD347ycBRSlFsKQaYgQ3uYZJMTLoOFLuf+5bpCPaQlPA4P1EprvqPpNU/E
QhLwGmNjD79AyMKJYdLqhFgtXYM+XQP1Jr2LVWjLEGdxhEfrX7aQUEVCl5pVRlXu
VctwK7S/j72J31Dapykyo7sAJvuZJBvo5h8dRQrSVPvydbrrhLoZ4VXhF9n2HWVu
Crp5Z9/iv1jbVvcD8v6ZnbP9zM5fWqp1XRFc1ur9UyMqpTLBO1KFJLdWvR+2otei
vTVP73GiRgs1r+WwC2iIQ4vntBS20hUAtlxWR35QGIAFl4SQzcr+2CxitMgzJYO+
F8JW21UlzupkbEu2+4MwC98O3IjZNqXwApItH4iExXjA4qI+yDPQtx1YEcy+wS5k
eZw53619E68bn/r5YfT21mWuuzaU0qppnhNrbTuJ/CEXovq35UfbxqRYM4jHlS5E
i6lu3OW3PTL6hnMgg8298TY1qTJx+dNIdsTpq37APmj5bsdlTQKaT4ukEkt/zR4t
2GOdenvEhXigKfbslAD1LwcA+KRstc/V/6aNd8AumrNvr1EIF/zS8z1SM2xruYO+
GjWEdX0+MA/GtjhhxH51A6UWuEZFpu4r489QTb2HCFv/k0SNMH0eVb3B8QEHUGQs
FjTyykMqqhYT/WTNTEhEagiUTgTE9AH+TtWYDgAL9Wh5gO+frUX+gEA/DeUL7D5j
n0s+P9wu2GtqNyOlu7zySt0/xZXPWCDpacyNGY1MoWA/VX0gn9admavTt5ctwouL
tvGdVrW/iWJQRNwdrFDwh2Oh4bmkltEvw2OcWmw6Ny8ZGxyNMgrLYOTEi9Df+92+
xt/A1i1QXn8bIMG/lTEOnmL2atGEB49gue47lLaHX4RwFCHc8V89RkT0CttdK0r7
FI4KicK7D6HUhIZXbWi5Dkm30ZKyRuZx/6B9s35C78u5GFW2tHF8zJo3IwtnzUiz
VJYCCJzq92ZH43PWmJb97/Wqv22y2EYdOPWVmCiq2ye1q23DhgiSl/TdmIKI5eJh
5jHsiodojZRnKb2CTj6g9PQNxbSUMbE/CAHKI2CooXoDpg3HGLg8ie07k7Ij09bZ
T3t7VY5PngZzt65e4Ezumb/6r5PoW/aGOrdyeWEpjcA8q4ga/adVXkImiB4mTqj+
c9Nd6GCRXOeAVpGjlMzRheIA/JzxcFvsfV6dtieYnEItkkWFWzOfbNP8IH+q9F5h
1Khcm1w1U6khxVXpuwTPpgYElSxoYnmTNc9bGIQHhkdC1xJWcOXYHXjemChg11CD
sbGGjDP1NwlfTlsAq4GmLJD3WLZTexlw/EUQiRHU2pUaf2i0dSCT3i2tbEKURdZx
0nVRPbugxfuSmP/yFSudageCH3uT1OLm1RHm7ov9ktAsOsz+Ldf7WZJsNoLBl5dc
5ltIR2QqgAt2fyT6rf4K1fGoNJx+7ZY2dhg+3GybmOP0YAnQ3ZNDgOdU0c6ETlV8
SvSfXq/Okp+VSB7vTN4y0ZZv0qAPDEUnauGTGD9StqQhga3BZwa8ctOS3tiJ+1CN
Zt+XjM8D0n9i+aQPBGCj+LRolNMM3cCWHQDzE1yU67AKWPkPj3mvSQdpsXQUNnqZ
ncpVofPGjm7IhXPRimwxduExdGZOR/QhBRRwOPX/ncrx9FgsMCQca0pkgKRFJLJ6
jjO/2Of47bqKPqkzdGAnfoA0vp9IeZG42MYW+Kxn+q31ZPnrqQKnlI49RhLjO1my
zUk1Az98mC5nv+ivJBLPju11cwbDUmGJRSI5aEoxx/5xa9JmSAi77+CDlIYNPoJE
8wWKlKRhreN6Kt4V96bpPqsAFcfcQ1EhFpT4EGMBg6roQOamIlSAQqt2HQVOCVtH
qh9MEcNXHjOTTQXEcR/yanRdKyIuhYpOgnHC0z0jGuIZZj97U2n6lDMgfEGb71E0
+5usz36vtBs8+pxy26+1bX4IWwlv+Gcp8mc3/zKexZiPfiogZBcromUvAkqbbXQ2
epxqhnG29YgnVOv1UcujQ66r1N41tbWnHsz4q+yFowug0v5R8z3hhBTJctY29x3H
0/4i73Bueov0wDiZ5L8hJlIKsyIGygN1H575rU1zQ074FnRY8VPdLbg//EuEQC+V
1pqhkuEe+P/vosp6MQFJgXRADO2tOAnreegx/ZNj/sBvUtXAzMFRTT7Ue3CWthGS
KKDiY/9QAi0Eb+AkC32uIzg93CAuo2mU4j9WfWd+f+IMEvOBw+20YetH6kfW3GLQ
5cfmXuc1ycs2lv8O4bD55cZ3WEQUPVCTpVrpB0GkIA9rG+QA8O9q1+EL/5Ss0q/S
+UBc/tfjadl2aWOt5cWetDjWrbyQeyc1N0UaGxGq2t1iEdkMwicQiBxm3ERtJ2tA
IYo27Tk9aFWmRkshVkVfD4xHp8ZzTkGCpvIyHcTnrIKlLZ1Dj7zcS84s8Lsyrq/W
97DIQBBoHWSs7RHJ7kqEh+bAnTsw/KRaBNPmm3xlnCsehk3BYWSDHWY3WrODzETl
ZX1Ii1StY/zMKS2RshdN/K4vWLwr0qvBOjt66PaP2KLQFBfYT0gq9MhANsP1MfB2
XQbN7KZufW2JwXHBHSekWfR+A650qH8wdAmIyqIPBRO0L4BKgkUm3vzUPViJLgeh
g2RBwhOdwlw7BftVe3GBJJwHyxYYP7b7/HZLh240I2WsVbh1Xtj/GWWipXS6U3bc
SlPo7IDOEMeLyzZLE290wnUidy0nT5SmpVFgZjWfz6u8wehk5t91LEdmR8in4Ssy
2cnlOJx8+OxF4xHtRozh36xOXGFLIrkcb5+MLQ1DanSYQw41wyeQZS68/zzl0YYn
Ivm+8pSD7Y8Kg9dtV8ucapex3S0SDpZwFRKe+hTVAhQ7lUkg97zOwE7WYX6ucZ0Z
ItrfvDtD4zdDEu8NMkoZWo/DYISOjRvXEJClI5jy1TocfbvT1n6I/DzbGnUZPmhL
5rHuw/j9ZXbtdQJ2YTjZmejbg+W2UKt/j8yRAGedZblyovg2d0vVn/7u1BUezPBP
0qOUCuGGmFWGXPAcAI7GhacCVHMocHn8Yitfb50El0mps2lxKbNWvtwO9QyWLN59
squQWXDQ6FXd27nkMt4yFwYEvRXM7WJmtLjV02755LnMPrjsaliuv3jCsIEW5/3z
3pKVwQXvsuMXygHCW7E/c9m79KgPfAjNPpu7a8wbMAumjUMeBz437owZCYygcprl
R9othl3LHwYvyq4o7BrGOWsDbJvfgP3eouCtUWtYgrnnyEFu5Wqry5ULqx0qnTzF
ruhiAGTZ4fZT9+jPZasCjh962ZroxKx06T+USwo+hW5qbcttcgoy9pP57CufSbVJ
nH887Ai5oez9c8JgvmH9dcVzymh2rVWtOejAItiFUysljwLvh0HZNO7x7kn/T28c
C3BKRW2vbjHnpYy6Yasj5EF8z6gQWpAFzEhPuIMXAOvEa+KrsJwzg16rDjNAHXpF
+swBLbNTlBlwUzAXZDbqQCexUIhlThE+iB248NWexFRpwao0LORZmCtSB6vtlcBl
Ut+CxzIbDKdBPpF29jp6u6/CpDBx/6uaq8+xz6Ev2ol6SkdjkIxSScQyex37mrnP
06tl6mBUscJA867wazXhQxFmJhcSj1jctAUG4YiVLc2+rk7uLD0YJkO2D0gYw7G1
qWaKFLNbNjc0WcN7LOZ+CNr5qe2DCtX6KThfpIMHVH5pI9cv7YEKK5FluIv/SpYO
/ZACzYb4s+HKwSPrM6iDgXpWwAlqkMzwOL7g/etvecZhDp9Ods5JLDE+Vtx+FoLr
CZ/KKNzu9mKqNNZw12kzFRcti9X7YO79UP6e69NR+1CthdhnNEkSCv3pVZFIpys7
oCmJ6IC4kCWYV6NHuD6oJ+Hv0HRVeho6lwiuXUW8Uk5kWsxtGrPVkaBRQItG/zVu
e2WDBnd4xf9e3RUzHfUZb8NUcXDg4WtRVl8lCF3TaoxmC7oS1RjEyJgXuch5rEvp
cp6ENvketnE4AKdpy9zCk1Jpi9ej+eF9bFIFjCXVveINLnVCv+57yD7sCy+mFweP
cGxCH5To9VPt0hfKxvrgNCh7BAN83jTMMbchqufI9Wa2MwbE9NnSO23DhFMHyqvj
laNvgTev0rIMwQm35BLN8qyBexcWkAMDaHaFpduEtg1c2NQyeoHxtdDnHcAQKplQ
uqaG9LaBKoEwWix6hOeO/iye23sNPa4aCHRuEhhBzpadq+kd+phLXqv6mWpP38lB
r0YfuFg0oo9Dtjp6n/Han5XoS29KmRjuSaJ8HTC07/Na9Rgv2I3wDGyBhlcJwKaW
762Dp+77KpskwYsxh+xAAu7a6ZEU8NhQ0teZOrg7Peg+bdb9dqmmRMW0oz93+1VX
bMiiDfBOULNyU8sQNuyODkVbxzLyxHarHaVG3RRsSm+c0eaju96JebBWxGVJCFBu
rEQ6vk3Q/+H8+odpxDMSViyHMLspWFeOl+ZIYdGMFllH1bSCwkJHjHa/4FUPuqfl
52ao+pvFNp4WmH6EfNvAXS2iwErE24SFY+/xV2vVog2YWQ9WRYygTOhA1wpGCluq
vus8SBqn1l8cH03GLlxdTW0Nk4BcDoE5Y4c5NSWcA4ovpa9dea9a6+7t05DrHv6+
N5SljgKQzlj2X7sYywuNCGv07Q45YL94bXdLHuu7R23VyvF3tDwOVtlbAjQ6SgPz
20BqY2Yhq9jZdZqLmZWlIbKoaDCVJu7FWcY7WLL2jHDMlh6u/K7Jafp+icMfOFk9
YV1nnENl905gDOVOLRqFh9OJ1s9QikaMPAVFnB/OILCvpxC75nTpqZ66tZSrFe5l
tSGyjNZ9Wtv5xGIq5QDrKmKhW+y3EoGhFpN4SKXgtSlPtjUwC44xPWNO5IXR5pJn
vUj0Tz20YDS4n94rbeZwu2QFfhg2V/8xI5v6q3wlkgI7I7kcfR9vIECiCwBkbwMQ
FznqNs8fnxz6Qwer9vaD5HXw9Wt0Mrx7HDb7Cs/nIOOZblX20WeIV9KNtfFrnMko
iuAoDYeXKh2v7somokDlNw/lBDnIREzSWmcpIsoLSh0rJkxC8yAQIgLMo1LY7RUX
0VmHr3cwgAQm4R8yjEG27AAdORwTYwQ8r7ZqbXEwmIDAw9VQXGtxmGVOTUSz+RwF
AVwzH8pXO+8yjtHFwPSa7A/4rE6+uW1B/3exBQ0FbeULS3uMX4iWOsZ1+R0ZZfab
LeodKMtOq/s3oApGxI/OB0yYdtOB0n99k7HhuPV3s2S6lqK/YqBfQlntO/cHIyye
2En+9NaGiY/9t/BllPeRpBw1jHdXaF0AFne3Nr8KtoBmx377iILidu/iu3+iWR0O
Nl6JaKEi9OySfiyq5a8v/4nXOvMZPJInTKgDJqg46AnHEHznVRPNdM5poTUCvCJf
CkbCPar3MucD2qRvcCDWdv19otNz8AzlCPTZv/p/oaOaQ9iX1YIKqO8Z7SG5zmoP
Q0xmDHWbJXev/p/8NzmkDOqgQ59BZ9x7k/yGJWqNliP16owVLXCl3CdL9TtadxnN
XQgdbtnfpRNANKYqf0Xw8Efv/HCmULPp+1Zq0JNsaj6aYXYn4eRDkEqoIlVHD1ex
Ben45esXvhjcf+JDocw6OlrkwHbT0VbY7YME6qHljeIlJ2iVmLWoNaGjx+NCl528
GHYYzYrl090JEVHvyxI/m0CkLUw/SvCJhMLgsInX7k/S6iyntrXgXDy7qurFLK1n
jYuaIuXRVmoayHV98FUs+Oir6URUASiLmDKrSUNOnQ8hRtgrENBlNRPpd+lKEbUE
7PIfArRdJvobnVRigUPb/O1+CAmwC0ofqyFby0QAGmBoGcLBiNCoFR7sxN2mCAVW
heLuTPmR8zcvbGZPmtP/Hw8qxBsFPWoYMFpsMmKN2usE3kwmCa/sGnvWRBrxMKai
7T9iYhWknXTi1PHxhXsMbICPzjJkwEXMMxF8f+YsrFqfCITn/1lhVy5ZxMVeArLM
w/pJ6x6C1vz3qnJR138ZizvBjjXerfzbEd/yyEHqV5Q4IM1OUoP/tX23EDbG/87L
qnMF8Nd1L4NJu33NUAM7bTRE32wUZzQrt5Af8ancXK1YYmrMNQsN9HzBCxCswF3N
0R+CGhWxQCmhFU8immmnr8XALfAXYRfbZ4VbfhfMxepgM3XXc0twCyPnKO+nrtJ6
fRCnJJ9vV7pfdcllt8/5mTvHnaf82ekNJIqV9elmuLBNh+Ql9m8BiQxrwmFS1Wae
Ofh5u8GpXl78mCofPyV3LyYBOdKYM1fmzKiTvQefdUVlki4PHyEYzvMn0UcQVsum
badrwcQ9kP59suRft01BUJTT8F5ZW2hUq+HocHmEtv7daR/Vbe/Sx56kCBmQE+Yt
gmgWPnSo/lORIh5O2pUIZYB2rwIEtpSC/pMoly5oN8Fggo8FNQmHYH62jLBJWnNb
fucB4YbOep9ileh9aY6EnzdV0CmN+RJMT65uv8VEEdrZAAh7YTKjCOClbDzoFvf/
HA9xfCZZS1QtbRxL3UWsoUJ25dItZITb34NnUAMQktS8VaciusGOPGk5PNblJQE+
MKuIcMwpPaN1yiuEX5z0QysLsFgB78yziupg0W/cmyXchZXIJon+9R5Q43r625I6
LTbBsqhAZ8e1myiuEmJCgndlUJNCZP6zbziMi7exJUhL8UX80GJutf+ThxSJNzf7
9VxAlaDvaNj5V9YttfHFV9ophD55B+6ZkJRzYn7LeQgOih+KficAEs6hPWzNUkUe
7mqAsc5yUrJ3ps46Zkp9nk5Rf42GFDgrwpspGMcOLs54/02RrTzJiumevV5UCxS7
UUtWOLZscvGUOjMe0j0u9tFBOoa0JNc4lQS/StiaO4Y5ZyOq1cTi5bF1L8mAnOM1
lEADpg+k2Cc/Z29Z1z4wW8CcM2s5xDigdnjNae18GjeI08razzKM1g/YNkRmArBR
1JKQ0Plj2qaqaTnY8HB9Di2j7f/9R5yAw+54p1dCipF9nvIf0i+ctTYuFG89ztBF
+CL4A9EFT+/RbMariFebxwTljOWQglrCWFSRVxWrQgfcupaXWjjK9RBOzR1t+4KP
q1GAOOztinwIhrofuZ3s/9yhtccxpZacbFPp1ox4hvQhO0PBvzo4GT/nUQFqRdF+
CfOzJdE9kM2ZHSiTXDz2iyT37AWNv9xFdD+2SVqN14pw1vIFBYQ2ZubHQcGkFmEu
xKnCXK1DgsfOdFE83VdnLBMUabK6Egf3M6DHHGLrvABi1B5ZSw88X2YkD8qB2zz/
OgW0Rs10T7wutu5GqWYk4+PLRxnxOtJG4jDGq+Bs960TZtQWLOcBmjZ6U8q31KRl
l4Oe0bXfyeNizvq972l5NrgJkXNawbmw1ZJbF6nkyu/HANTyJa0CVm1c7YVjinoL
Ma2iVOsPnUDhZAk1JjGQYUipuD/tVa3Lulkr0rAv/eyCEBfxCR7+AGvhBY/XZZd1
mAmm+PnBNjzKyuzIklY8m0OiM7PWZmhlNcOesxDlsPiH7M7Uzih1HDfb8ER8bxNs
50PCT1bLOgvlx2ZmWZdstf9LSggw5GrNXhuL438rOLU3CzUfjlIu4eJF4bSisXcY
oYN4koFSntTHT9yQjJ4e1ZPtVMnerioCkEXgPv8iEX8p/8zl5PMdv3TveqqEXh61
RGzR5acbznlYG0MTsAT7OLsNKMTZNZmDubIGmuLOOmx89J+UDIdkDFn5c1g488dm
VFFGAux5UTlqXAMXTAparln+5nLKBoS7jVwcODymOEhThQr4wo6tUPmnOS664Dz5
VGtYG1lFp8NQYRXltlCXIAPy8TbKlnou5MYcEhxS+2/RXvBDviZB2346SRTLWYtQ
gUW34FhPsUtp2SkHTRh8BmK2VLdIylLQkF/y1ZMe9mp0AfPzbjJYZsIgAQyzQuXm
h9BCyuDffficrKQr9Y7vSkNuJWr20hb4Ouqmgucm3SaQTvzEmm7AyFkLXVm9JcZj
fXColODkAxEB6jUbiAMTTXVEyR8I5MxjYFPHywhIruOYUkXIyLICR1O7m2EIYklC
BigxeGl4M7wP5P8DeOyeNuIrFIOqvKlirCdfMhl7J845KDjKrOybhuZinqflLLzI
WvhzCYlmyp9p7cspai4YR3Knx1Xh6ZVzJlW9B8RLXxbdsNAzPn/9XqBB6BoMeYuV
xJadlrgxNBqoI8izvorQtkvrAiKReUgAk++p9yrDDIfGmCSJOHe19IBjdBX9ZaFO
6kWlKj0ZBi6sj74uACkTipkXWTWEy7enGT0+gbF6X6HNjIRVIMvDnOp7k/6ambZb
o30lh7e3mmLM0wWaoP0tO8xGADlde84ghQB96suv8BjZCcLPewZITpTdzkz4EpNA
QX8DJnbXeBZdpFLWBJkcJOK/cvfPwnVo3zxa0/q++G9uiZlZi2NW6uITiFMsUqee
jBXMQF6ngH2VqN4s2mNSLi/HamrqBemowWNadX9wnQPGkxZ28mtUPWLOG/FBv/Uh
245C2lp2cZuG32vuNQfZ8zTrM8Pd3M+ymhBKLGtW5IC1DIRxedLTvXuKHAGYctjZ
uKOc8FzKAnKGV4OA14JvBRc2AIHVI+4TkPnE9xk7zEIKebePhdG9UagQ5j2v5BFc
17YZQlhq7vWyC+cjNuja2LYmhFEqedLcQREcBxemsKBWtZnQUH72Fo31Qo71gj0B
AdvPc1Xqu/fiO4b87SVzduS52kkkanfkf3oF4ex78GG338W5OxBBgF+MyeYnWdse
bnYXC15Dw7FikGAn8EXeY/Kbwa2wESKr+DpmM+AcY/6rtbHSVBdzYvirtBTaB1Xo
cS0jwBbAYMj+I1G8bWLuxq3GSNhFDUacXSz2vMXWQU0wFaLDzAg/xQfyMGiXw/VW
lmuTZcTWBCekyphMyCqBCw/Koxze4kW3WC3i3tUUvcnQYbc2GMAt2ed8Z7kaGNhu
RWxGVc/J4rcBclXuovSWMHxVIj2ru+oP1XsWYWwOA2SNZypnf3IclvcPkJts/oVA
yzXwfiRogMNBNZ8Mkmv4yaGjHjwRf3DPZGVYzvWEMOrPLkWNfJzEvR4Cv2b4Gm8v
6MViyUdpftJ1VRL6OwJTKCs0WKDfABNpS5nkXjZ5krAIP7GzldDF0x8i6Gz69Az+
w3Bqcj35u88X6I8V+IpAkvveCu17t1PSLpqXwWGnF8/CoV4b4hFqZZcWupHkf0QI
EQNymFt0xCPEVo9VfIlBh2RFsaftZNHnkSfttfphkRS8+UQmh0rfIj7CFn3qEoUw
lKAlGb3CVJOLCONvaxciV8HqlF8ssT6hNaRp+nxpzmfoy63H89tNpV1QJEOZd1Nb
qLM+1Dt1bX3KtGvOrBuRajjKggLh88M0y8maXOif5J/wXJ1HzqEo3VdlpLLMZzjU
NJ6Gd/ARKFAnPFU3Alm1Lf+IDg3PzXpa/3LiCJjyInR/PznwZgk/ATQryylxKMBa
ZsElBEcDVC0IyZ0KM/gKQhGfbXkiqvilN19/FjdWAtuk3QM2SJKldpTXeW5TaQv+
KKJjLJ+HNnTc7/I5tw2UCB3KBPr+XOlzZUnJ3KPS2tIEY5KKDL0CiNgqAbwE9Xy3
n5firjYKcsW6zvNYA2P5O+VR14+N1DvrYBUUvZhNYEHp5QW2Q/vPFGiMHzCO1KaK
A1wSCAc7NrLNlIdlPMT5C9LZam2PK9w7NYdY+ug6NLGlM0BbEJUz3oldh4t0ggUq
ZKNaq98Nkl1EX7G9dMfmiIigO9ThzDhST2pHZG7mo1GT6Ky2c4/JmERzt2gIObNI
7hcU0ksu7kTPm2PXYDc007Pgk7c7GjfzPdAAHtF73qjADyxzJ8Ox45OlwRGyCdBN
YWa/lOlGEzPRuYh3T6gsbovgfF5mUGrK9tM+isw7j3khiyGIkezxVcRglqJ8f17Q
VrABcCC6FNkRdYxbSAcW9C1l+upY1BDcPSb6a5OF2iwEs7R6h6KBtXsByR3Gm0PV
ySlmHZK5jlg1BuwlpX+Witg3DDdUVUNegKvOZnINIw/1ib0iEQ0reXuwKlwMpXMc
sELUOU8i9Io+mNH1yI0paNwT9N6hoz7J/z/QJPIbqZpvBb/E5UIIXYLtWPFBU/JK
B8t2LEziNsc1Zreza/h8+ZtS7t+o255WXwZ0ASOpRx/g+TaiPL6CbiuRQFg+uaLr
19yCRrsz6DA7Mh4/t/7rHisJu7Ribbf13bW3ZMEcukU8JIs2dzOEKfaTVTWXnMtE
XUQr+gB2EyoYB7igZRBVz24ooT3OhOJPXEu0O7HJ8AHQPDM4/DeMUcmQKkL1Aa7d
IDEPU09+qhVrDXh3x0jl7ftPJwqt4c/hDzSF7TyFKG1tfHdGne4LL3g0ywJPx26s
6/oTmEtcu68ZtpdyFYhdrPo3TFaZmnkMvDsr0MvOSOhKGDavv2LIRV8LvGoAsj4f
r43n+0b4xvsGBofsSuEf9h/dXz1VGHwfsZ3Voov5ny8a3EYhD603czzSr30AapS9
8nBTrv2VBxD3qVMY4m1ItfS/UYc5OAoHjKZid4hF1f62XE8PdKU+/w63X6csEy49
tcU+vlrWftPAWvgyEj579/TLeRNJubxYnr8QY0Fujxy+ZbFcFVVnwCp/E3tuiqTf
cgIN71BRamf5qtez4wPHbmjlzWlSgIDgWjtPJuhLlrtKyRQJsoXPYOU2FqIFZq0j
yNdtIs7I0zD+f3rNHvxoBOYyIxLnRh9tsjM1b39VqTNlkCLv2h6153urtFmLWlZM
jAiEWGuLyIB5DJxPHd9U47LIu9+VC60dl2c+TEa5IElLo06KSkKJ8TgKVLJC/HZg
S1fWG24DD+njIYdn7MoC9VnhEglJSGfppQUtMso2+PgKjNUOR6MVh9Dt5X9b6ben
SM0Kqwz7Awuyzwy8SKiBwHpQw+DJRWA1XNQSDdBmhYwG1x+XgqlO0E7cYy1HAnXt
Euk9NxmMfe51gcgUWoMTyA4W8N9HyLoUJFDuLb4e2OmN/3bl+m7UYO6dN5kv+bcc
SeVrVfuJ+qdGoWPPaOGLcuG9xXMAb7zHC+jBnUhxu2Y/MhCRijjpWZzJFUWc/fGc
J8+0sQQFmtlTwPANljm0IvO0T4CP2fPgvTNH1ZMhPxm92aotCDRqIGX14qR0MO+x
vcxflHCiOODZhWxzhXcpej/fiBUhv+7703DR0fg936sBErEB62SED+PTQp8ir88J
SW2jv81+qhLrVSqO276GWa7kp5SwgKll59LfCs2InyjQWJU09T9LMwsz2bZEdXqF
LERKzHdm1HCKjLuHQ7u6Tx6VL5NRk28yvlJdotVMu0AV7uujUK2ZMLQJK7f7+bhm
nr3xJ+qj9Fx3DhPxyl6sCcnV7kIHP5gIDNErkLSszRLOYzUOc7a+zOoAoSw20NBf
zGR2p89m8EvoTapGskaYOWDcW/fjsfQnqXFFWa8WqtSKNTHanw3advoZa1b3eHtE
xlp3zEWel6cjX16Fm6OmCJ0mwaSPqf9MEPFwyyqupZe5BsXYaD6Kbt5DXYJYV090
oeGynsraYuVqXXXD8Qcte3rNQTL4JvfYRjRor9C+AfKWCAGZmi++9OZHCfXlnJpj
apmBmhNVr4acCP/SiHlrsqTQSwEElxadliaLkg8LoJpMB19Btxnkm4ch5rmm2NeS
BAi0u9uroUkxaCDvVxTjQj0TKuQvSy6meXmDMpdnKerPAuRLuQ0HqbQZT6Yf11b+
bttGDb3aHPMGfwFGsJwh383a8Fkmn8NEal78ncXsIfEYzbOdynhV9Di2dU5MgUwB
lY/OplUoGXbgd8RnzP6+SCoYYrNLVA3ODu4T2XBUm1XEU4FD5nqDHICYqh7Afh+p
bg8vYthY3lyMMTuLu5WT3URr5oKod+JEmEKiyNiAvjn89hbRWhcPqX31WYRAEwgM
BCY223EoOf/6oks9socktqBL9RZpWQv4yQ0P0RD8P9Vv11KxRwh/2XRjXBe83dJW
lNeVLBfYR/re1lB5+ejWIahVOby0M2tCojf+QKHJfWr6GLHLobquVVrXKVN32/si
K18mJUcucnDjYekynRuZMJKvPaV/EnOkUaXIv8nYARdBqMI8Ft9xexenEznCcybb
WMue06Cyw4r4l6arjT5OgsuF984P2czsBdQnQErYUZyX0EOiLocVpnbHCKDYr33J
eoyDWn+x25DicUKOPJyPlrzNtHPOGtaU4io3rWWBGTf3Yfai+ON0ZQdtt3K7AS0u
wFGJCQc2fMhr+eAHslzO3c2z5WgVWvntPlskPildOTt8gK5794wQx8lGefGWszSw
QMwNuulwGi70vzZA0DCWymWpR1O32FZR7xtPdzRgfpPGbAkUqT4WCpSRUjXk5x5E
gqVPZ+V8gdvwq3chngGZzArOkdCfXyaNw4RyIpyYBgNXuNxlBzOxW/JIIqBXbx9n
Ef4EKbN7d5pqXw56QyTp5kQlbN+sFEkebFQVz1JKZmJgo55vkwvwFoxERuXcUXpq
7wCigT8B6arhR20fVKK11YoEmyD7F6g4HIudj9FzxFRUVsG1JecD3PkXuHk4qteV
oh0NUlupSvlpmMg17CAJxoiH+0a6d/4StVOfzEbpfnlHMDgvtvyHSqfrlEOWqgRO
IbmTSwIf2lzq7Sv/sIiCco8E0bWjqYbhQLbjzE/Doxk1VlYVk0K2xxLZ7eT6eqx1
/2CrAjn3/GlTRyeVs1Fr/KBETni5rhIG6wHcK1He5j5A7aOLFVKX6x2CPtIrzXdj
vS3JcmFGfsq7wo3fDJ1hZzQq8YcHRga32VHvrJrMUIet5IN9OZhM0pnD20HzRIyl
WnrGrV7/2PPlN29fpLFeTzOWfCK9iSygATsgJPj4ICqWjmD/wySw16TXRblsEaeP
EDnKKCKysViu5X1zk/SknAIlAl9lKWf5VjtkyUUZJ50eegmdgIYWVhYrzQRJ7pNY
FbUm9R0GPOfvXFgzEpL1BZWlteEXQz+aTWK4pWRViufd78LhfUvaMw69lZSKiCKd
LcC2ptWBuBjsJky/SzrLKG211QESdva3YZn2NpHm/GRbQ5XD1OoWzNTNXOruC3NT
UJ+PY3mcwc4iGRS5AC4FFGrDKFrOwyx4E9QQMtwJlEaA5cjlvRRwVIqDMMzmyjw0
FZgpsKpeX/y6999y7ts1e6KgkKG5grEbaXBllNORH5VPRx/uaQ90RfKDzZSdbT7W
7RBB4sMI699d+9+E8Y5AiAa1xhtt6CTDS3SWPq4WmDCQGcwXHIB9Qw3CYO61MUbu
AsEAae/nTVQvyeO1ZM+JkgeMVaXbRgUxCgK189MK+CaYYA82p8iWphfe8rQgi+QL
VWCmANxBfxVmpGDvjTf8NXSqWiWh0cCYKXsbwAoykwvOmDwEi05cPhRsFPR0LB6J
CsaqP2CWGYk3wIdjVoLTxAfzuNEYrFIislNgOGKSn1hY1EJFV0D0/obYhOTCzGwK
G4OQ0rN3V5MxKybyi1mFz/RwolMKqQlu+GHLzpqPypM7qoGUTbRi9G+/sKM0QeQM
uUgQqMyteo9ChukFFFJq4slXL+4oTQDYf4Bg2hYxO7jF3beKkSZEtTTFaObe3Xbb
b50VlpXZEftTI9qW5pSQmEYdZ5DTOiLLYSH6Z2AzFpenKTb3M5tGXOiworZ2hmbo
fnbrtArdA81vpyP33v1t2KQK0vJ2JnDFbxWLI9v5l+KXXHqHrgdiNKylLHOHesw2
XGaI5VANcO7NKOuqJnxZJklHgI0Xcll8utVbDlSg6bPN+y5gBlK1Sv7lzmYBZGro
eqYKdbIXo6bAlp12vX0ug1yLHZ9fWBezC8talIKSjvhfH2xRVKOohlHubnEvrgkn
KOQnqGWS5WEW5ap08sqJMKnAcq3N3Uac21AVoRR+dxwwymqBf8VZoIc715+eUT8G
Xnoc51h61YlkTPzzpTTWkdGfZm3wxNqYUpsLzIHkWfQFizlDsED4/5U+VodPqTGC
7TW4jDUweewql/mW3mkQnZuZLUex2V/YUJhH8H4FgJJ4I7BBk+PBgnRXd2ZP8RD4
FdicnJLMBe43Fs4C05c+QujiT11IATSpAwAo8MFSAAoL3LfTk9W9HemEcJfKXk/H
GyQn8wR7SU7o62YYxrrnSBTYpAoaFzLh8/N8j9YsAt0T8jQMM4C4yg6drkBmG9W2
/uGQAHnfF80pa0VWCL8iRng4eoXt/hzO1D85/OuvP0nH0AA4ZylCDvZydlmajAHg
ByQ5x3UwJtlxSFW7nB+UgrtcW1Z2Mfv6UCRaFNJLywoXcscBzPEAKjo4bGVLCPwo
0hcQImaYXjmBUmORL3whqvIAyr9GJ13o946jiHFSkB7icRAAiJHcTLVSIOps0RaS
nTMDcTJvESE+4kQURB18uV9yGO+BcectwOtVDr8ku8uDLPZha8Q4p39p846LAKbS
+U3x00JQuMOchZq27h94Z828LZXqdmfWBpfMXzltRH2MuMHZXVoKXvKqzV0LT4Lz
QsCso3q/xvI6wxwEV4A8ooTtqZ36qhvC6cVX/X4Udh8gkS4fJt46cZ/HEw1DLrmA
PrJULug60AcJwwgQ+nTKMeLax0SaMOV4FZhZKFUj8c+KpzkbvbyrhJ7XBTrSc8iO
Mvkv5ziLfytIra8B+KtCwAWcRTjWe+3yBqmT8Bc1VydLsFiVi2xBXY87hryolyLI
DpKOJdXUCIJ2yrXsNy1CkHLZKAyBUJ2fZqWu5U0P67ZvsNi40fTV/buCW1kN7772
DLyQ+Qna+m14xKHmuKWVGfz0x1E5jovlYezakMjMwG5D4YZurk3Hgmf9JcOm+Z9U
LGluMCTRVbqhrdhaYYPo3jLHJJd0WuzyCGhsHcYcrG9ZLPSnM0wl7KtfzHEPTwXM
dNc7bUxL4WEOfmz7V6RKB/nBvN3vKepKa8IYkZ7udosgLeGFEmGW7IqHNRMcQGAg
ILduBqyfgw2Ig0aqGlVB94m1pJL1Tb7c8x3OwfuHAVDHqBkddFHO6AlW+TwEBUMB
Un1o4a4xtcM86BleSLpqfQI165TtjLdUoa5m50Pbj15yJUqu2WG4BpvmPUa3ck8Z
/G0bKEr7xR/txRK+cgRkC+gi53wcRmzzPbKDkRZnyJ1uxj21B573gCF6eDlxXt6l
C8rtgBrZyurLYTwx5CcLxdE8CtDYs649lPQaheY3FUuT4HogMFgrgPv0yERAP4fL
NXFXnBlI6sX9gI00uiajVeZTVziDUhPr8ytQ56EG2rdYLIptsbKlWhWu5Dan5VdD
RSsq69+KZVlkOOfl+vmGakdUNMTLleh0hJ30sNRs7bZUM7SWsOGsGPNEqJsuWCxw
nY6WHz5jQVC5Lpm5xM7UPCnd0JTC+FWC3C8F2RjzgNkvcI1Ll6xiua7qN4cy8/ci
TjSPQWBrDtn7SdvrOragqzSkvXeTmF5mbnthBDXpHU4Vf06dx+j4CrqFvcB5xIFZ
Pk4BPgDWWEoHkXSyPpGIX0rcQdFt9E4T63IxnSSSPtTkkKzHY3Wr4tem55qWj9fp
TWGu/5Wfa0qNYpMrCrdlDhPvQlxwYtI/59FRNTylXubazd9eue2gYBuCw13dtEo/
9hKcowHQpJDQhyg+uExn2LBRXCM22J8P8xPtGctoVcC4osDB5OlAYKlejDEyTrmf
jTCZeNTDalYn/3zNCrp+bwq2xvxgsVsaybFzidCSyPZ81PC2JKFLHH0BWTEqY/qC
mZbHphp/6R8xK53Z1g6iyztMVVdjSA9NAqSVCBRAnluNz6F5BsSECmUSldr7HUzE
WBgKFcyh2+GaH7AJDvjedt0odHf8q4ZI2mzaoXN9JKYfysGMBs1KcDMtjd4wCkS+
o8h1NBRObFeP3MDe+0akEzZ7u9JXUWTMbnMtcPMhnilVqV8XXJmIo7XynHGLn2gX
VOTcKVE38roRWpLd6UlMEhpSjCCgrzuZtOzIxh54MGG2E8+jNMVHMitrzX225Vvj
J+eSjiYc2u1RhoEfS5gqJqpEq+5C0IJP/cFsKSQQ2X8GtTQ+vuGa8hh6DELv6SuK
tBs3KumwmhWPif9FLrR2/b4L6FdGd/62Sj9UTootGhKBFCLf5lZdMJXB7bDqtfcG
R8fuAHp03279Wlwh8hUvprHmJHS2Vcu4moW8O5wJDozpMDhuOv/6wSpUAZQXf/cm
scEZ967BHk2/OkG0i4rxDEFP/uUtJYzo2KoBrWvRViy84rxT0I1289Swd6Q5k4FP
N5Zvoc1/bQlEsk+O7VEK5iJvDVntcG6VwkU7ynpPgsKtwgrQAkr8En9TpyC/xalA
vs1dCDLfeLKo+kwrKNO65ytjEy8IT8FutX48zwGil73xT5DxU1Aibbpf1ObtGjGn
N7Wfm7L9FCocYD1pkplzlnNgFh7FgaHGUKnPWI9ZcxbTH7EApLne7ycEFZ98Zbcd
fD6jhGZjiZzEOh+QU2QuZGPShz7RAFHjsG9Mgs2YFELWWiNCLXlMt2rcim6jfFAo
wW9qnrCnBvZRfLkux/CGyNluu2ZFmZ0Bmmw7++/kW2+ZyVoFyotQQrsV0uoGxiUh
qUzRZrumuKnHP7tyTvcaKFAbKObuXm3b5EjZfKopnd1xCgmUmbqQpiZDJ8EWTyx5
oAXTciFHXNKD0mqNVonyAvulEorz2EfQbxY7wY1GKMc+guFrB0M1eu9Osb2ZTCiM
nlQgR+1xmWsPMviM6YOpWwF8thiin3070HeSIKVGghEpjVkhFJp1tHwpDgdHXK6D
Ws7zrx5NBmbgAykZ6JHKSg9ISCZU4sXMJxCk/wvnUt6JWeV6Evqz9gdXP6dR8yJr
jG3wbs+T1Buh3Rtgl7gDXakaIzd4I/T3LYoAqwKY7/GtEYOZtsmaog6YTbArfAWo
533sFJsra5rDERcggUdd+duShLd/+Q8TJAQFKRcm76JtPBvKPkWvur/XFz3O9Uht
0D/QJVGkJ58I5YgmLuEL+cLiyj2a84NWzPRhZPA38XO2naTyprfrDBBgQUeBmD/H
k05WDECBsBbc4/wOOin8a4gzvJxlKV2AnE7rFRDtFrJwmBVxgWaV9cxri5mefsXX
jelFr5AYxhhzECR16rXOm2pbeMnpymQjLD1W3U+GIQ6DATPF9mo8PY+S/Bp5lUzX
Lvladaeue4JknsTGxsLPBHXUSIewHkQT8VjyOxo7WnC/NoZEGJl/23FFDMY+mGFV
W7ez/iMyhAFVr05MJKMsuJEF41rav2tLvaroz5/YrSoD96qHJutyGK1haQDdypn5
aYvLduaRYjxa1xYbDbIRh6jDTl8y+Ri49ZR5LiGkGqWp0Fpz6+Di5mniSPd7qL8b
N2lglft5u8vvBCmixfnTJNrtReEAI+4rU4M3dtzBrOpQDZbpFvTeL4I7bKUKI9v/
AHiEZR2lxI3cGIWtUw4b+Q6CVfQyq+vILANX+xKRKIw89ka/mysHTEjb7f7FMAH4
+80Wrq1Ul7cgr6usCV09QtOC3wuuJtIbjVTE/cljowtst2jbIKIbbuVlyGIwuLHS
W2yRwxSvPfaS8wMA5GFQDpSKAYm0AEadKlDZaxV8HIjerc4ors9nosDjUI5a9L00
PnNYc9iye41ykxLhKaAJ8KDb65XeOU7NFOzf9yYTtFC6duCSwOiZZYHwQPbFifEH
wuKjlnlfLmm2d0HQdP9kV6M3wmekxKPKI2ZsSze3VLW/UIyr5/A4hi1ei74dUBk4
945Se09x96qiggXO4wde/ull+ErqKY+lpa5nLb2OzfAOEMabrcYEcpFlKdC9dpuM
BiglKY+kLrZZQs1acqDzTszKuf0pNU1cvyBkyrpltrajDzCGFsHkuovZiLb45nyR
Y9s08fK4l1/cBFtw2yGvSntf8oEPWTSrcC1PGwzDEa9w+xmvnX5D1Ixml5emjqCl
O7j7F3oZnAeQRQG4NtuMWkhUH3bgOwBlps6LC07/PHy9M4eu8lAiCBSZlLsg29wz
4ICiByWADvcmqDenDi+JJ/3o3B33NB3AZLEHdYzV3rOxj/DIbhqJ2zN0IMk9DlaI
Lz7haekHCxj7+122hxJ6IVqE3a5JKPN5CDOgddSdkig9R9f+apk1G9PgpaWhNdXX
ZR37DirHr9hQKnH0zCn00MyE+va+hwpu+MVdiH9FN099sZCcUxflgTWrbv8nmblz
7ASgUN8A6h/TGPYGyDqkW5K02puU0J+iqJGFpMog+wL8FZu7fvKd1jUU73opm9a/
uiH2tbXZLeIMYbJylU6MBa4UAp50PM7UUJIx42iY/EI6t42Zx/fRk+GBN31brlgK
wk3ztgnb9iMgQtnzMe8ihEGx8dXXVpgUuQx+jre7wXlmfRqRUp16nERGLF3oRtss
iWmkkfF2TqTahridS4yHX1IC13DHgSHxPNEnjXL/lET6V6zgtdW7LC2J2LJflpFI
t0/8WN6gtJ/pYRfOIvRQv3NxzJdrQqmofvlGYv9Wf6mCHCKhmrvb2QeCCFFTvSPJ
ZxRIVL/Qn54PjyQezxp5KtPWS/l6IouzDuf9xP8/onXmLQOz/tA/+cGZFi5X3LrE
9HRo3xW8HbvfV8N0S3XgXze43hC/FXef+CSA1c8/zwoPdt9DqiWbfke9sS9WOsLV
610OptZUnm6X4zNHP4uKFJ6+xYmrddo6lWnhpMJOGF+gri53lK6xizBC3ZrK1wQS
285r5+m2PfyjX5kGraFoqHpViWqupDhu4uXY2/6z8XnTcTnWJVbSYUnNyoUMQdlA
KwwxJNTtEOVKXdsethD8uMKKh2n/qk9rwxIkgepu+aElJv1jRGiT/FgW5m3710qJ
cX0syNRLIMpev0XSam4EQoYEHbZnoSR9nMOi+C8P7dGF8t8u/77Hy7VWeQrHF0wM
SIvbZoOt+9EDN3x7TSdbTylmkzzp359f4zIgxVTYNvq69aXhevYwtHI+EULga+qD
OsfvPFqpTFkXuJjTnBRrUPMVhtFJbKIUI5ext8oJuvW07w/+7hKmQth64RE49J/W
bAhICJzItLD7qq/0+PC3g/ef+4yg2dnny7q+HboHQHYtURfOGFwl3/vpIZK3CI49
0nx6hQa5wjk3QsRIib9RFOOh+4HPEx8SZgNFZ15+nKeys9vVjwzEo623ejJ+VpIm
+XCuPPfVxsVhFqvztWAEqqxUODr7WOG0lPokVVbktcbUJv7czxIxeMPC5miey2GH
HvvxTFfYq1vJGsG/JFMDHFCIp376aIn/d12/nqrYVtjujwhmXibunsNSMPHjNfuz
qNb5JnbCNBtIV9N0YJdaz4Hx4PjGGmbeqYOIEiaWnerAcq8sjCe653intm0nlyom
VvxXpGo9BwU1wMjUOE2K5pDdGLj4FdnJ/RAgFejjFOPkgI4azhYeg7aQeJFxuTIq
DmD04FMdO0ECzAUpRIMf8Mb0bodjmZMhjbxagaKADAV3gSApvBTKdgNlQsPGDAq9
uNdjYGO8wp3tYQahY4zhOydWbh0lMhSZ6Hh4T/vf3UnuqgrfdkFF9o2E2R651nCL
JE1snRc7G5/QL8Hmn196rsOBaT5KWnO1Yoq4iIGMQzb3FA0tWhVfuPwjnk9aXuU5
rwswmh/IGgPJaqR5F3oReEopkzRTDU4wVwOGZcd0SO+0az1dIWG9U8jQv/D8Bf8Y
0ysZc4FcZHUFhTmAvCjjhPmtrAAnDMbOeXUIR+k5jExYRXp+P7nnTI97H3NAdXh0
EaA/Sxt6C87z4oBLZkSPAavXLL9Ijcq3gYLQq0aoU88M1LxCxE5CERapdHKoihJe
hbEbcIB2RSjsS/XwDTsRwTSRfn7jajYQp2WUEGKezX524giH98pMYx00NOKN5Emt
+oXUDamG1Z7Ti2YRH593VVeWd+Cmm4p3j9C460VxliWC0KcEHR7o5GQk+5NB6hh5
/Qsbn1lz0N0TMGW039BZHGjpLljrd0WRH5FBh3MPEZDNhL7FXFnFDtGoGtcZd+hs
tMouZkeKdWaMSmwngtwb1RnCwgbJjpsH7K0l0d0kyX11kXT31l2gG31znubTaekJ
tLZq1uy0+2z0qySkbKCMT66u2sx9aVWbKZhB3WbJz7MZtdOtDB3JJ8BSqV/WnoOM
PSpodO1G89vi6nKLiiE85JBDz70ZO/lbt9uqEOG7R0N7hfvQHHXwPUdzDsBeyGaM
+V9vofaAoPDbb/x32JzTmtNHSNRlHE0+KGOSwz/gs2SEfZcG+6HC4ZTClkQzW6y8
YY64DTGlw0Vss89j4n6zMIsIgSE4a1qMBA7qJFTl9cflW7We/i+ogAwLJfOf7RvG
rVETG3heSxCN9UEDdpeP69Zzc3tKq7PDOA5DrV8aFycnIIekpyBjLqoYsg6GAzyM
+5AZhZnb9UxPU09NACP1iwyGOCDT22Of0m0QrqkJfg/+EYYK0VqPqEJywBEkfzZ5
sXE3MBud/rn+xlfuKejt6tasEcpAailGfId936QcY7s7KQp2Xa9AeHFrw2JMR5bp
K5e/NHX0Zhlt68NFZskJKr9F6axx7RetW2lNIKS441DmXKBqNjoBczb0jNHl/QCs
A7G1cedB6INldqnZL8eLztsXEDeCyZGoFUv6IUR34rF5I5FbHV5o+rw5zhDsuFSI
tm67xFF+kMbVM+ye7Z6tMFFlNBEF33d5FrfRjPEO52egBDoWcNRILURY0s4OSjKT
G5guWB6cSCobmzstiv6OcDJmf/qXlCcvU9H6YWliT9aqL7Zj1heKdqOpgiJdiQMf
mps11nMob6fr+AnpwCBHjd+/J+V84FwszHsy+UQM20t5wTFiMz6zGz8Mdxi0Qcgz
BSFSDnb6u9rxDaeMpnIbwNo4SAVfUxcMB8KQ3Me2jlGxVgWS0LqT0PARz4tlR1i7
pqeQ70lA4WLRnV2+0I0BZZucMGZNG5+VuamAj4KjvLYkuOZHa+cXqfbp8Nvfq/V3
KjrxuwtecHXne+8WeCfiYSQmIUdWM0Am3Ko+F27D6u0lgELma45N8tnHYU8ZYgsM
vva6x527iVogw5IaKTrFmJW5EzdEy3r3bhTUmmDIQVVZmj1RC872o5PGhEcLAWdy
Ry6ySjhS02bVjmW0TjeD1gm0lXPcBg35yjXSetqsXZO8oGqxkEoa/CSRHvg4l8mj
LEadGunqkFh1c63nCQj+1fsHCWMgQZuld7D+OpQSdBhkXLwSI/izuorlnDA0R6Gp
9nV0xojddCqVw2BBJvvtv+n/mUtyzWgezM23PL8xw8upe3AQZQuqVGlX+QYSO7Pw
UFk6E3sG2jYZqWG4kpjb4XQvRAtT3DS82rbG6o0mHDaLnrNvHefFLzlCs7UwlHFW
UWpcD6EJVnpp1MDeJAhgPrUYHNnZD+dpxufIjETdkUK9az7Bqgd37yeGrhyFgQIV
EG3VAXcc3/pxJ/hCSkJgXEtbxLrrnPgxWsBQk2HwR1PHJjD6tIsiTMAI5nBsH2is
asOG+JAZuujPan2E9BxNyyIxx39zb6qorftJxUcxOhpu0+kBqdrO+BMTLrA30Kgs
Dex3i7cF0RE9oOBzaq7NIA5Y4XiQ8B77hDm01xxRwjvutzaEIhuX8ymlGwb0rUvr
S6iUPHZ9HRl3wn8bkeiRv4Krzch86z1xZyaHMLYOSEFf2Jah/LRvgexCgvPH9Q2l
2C9swYlD2qeXG/1DFnbsP1c0VcMdRHgR43Rh6HHMc7M+l+wwZg5bbPEdbS3Y9H/G
Zqj2coNmSZZHBqmCNpIN1VxITu63Yd9Cqw923c8KPdOOqGqEKTC98k60ensFzYsp
ljFvP1yPa55OBNCr4Q/enLYUvRt2o75z6dhM2+n08XibI+CQh9OFu3Xmuvxvz2tk
sLMVp8oCD4nbgfTZEvdxICziA4g2jz1taHyiRBJH0cpYK5LfGU6kiPsVOtHi/wCY
59WSV5eV5B5EAiWEpI4yPp0nOQstSIPWq2aUgnhLWGl1CC5rAqbCayWIxAIEseQI
0AgAjoY3VPGQoNjVXQyKl4mMtIIGMpjkoahOngGDgG8SnX53TSh9GXmnj3Yx1y8Q
GDXYh/KvX9TmUYmfBma0QQf731vlGjpWvC7G4k76KrTDwBYDaa4+DqFMF5Nu2UK9
6Czwl8OZht7N42Mplm87jH/7LSMacwUMUZNEdlUojsEhNP7/x5fcO0PBvDVISwyU
09gckfzmLBFpK++C/o+F+dgUHJMq98sNlMCSU/MlWW//y2zrh/e8ZpCCfoC4Ayiz
UfMjPJefXHg3LSEBVwqsjjhQ/9HSj5uLb3dXUWzSut8hBtAOXqV54BMKdH1ziSyf
0wc8a8k0cVmxYZD527lZmFaIqBQm0EWQFW816II9TDPbPdR50kkoAuMHK+sQEFNa
oONfps67aUlS4UZ3RAFZ8+novTRAuxI0hdMTNwLy0+6ON7WQaAlwrebiUXrGuAGF
8DHKM/PoVQIlahQs3KRwtiwHy7A6Yi/lpDoIS6W/hYhB0XqDD6YBc8Fi4xyLjZXl
5RRRj0QnAoQ9tSew49YkvVRs6KvrqOvU4JCO8rlmCnSX5qVGEdviOrr/hxdQBmtg
f+8WslQu9v4d8Qs1HuAy+8YjKZ7uZNQnANtGteXMcZCqViLFCQHkqPRo5Ks5NQEq
viGtZeZalwtje/mOQRZPPD0qLGYsSTkR2XBZ+6VfqDh8Cn46nIS4+m3WLzmocBkw
EYzjGBJlO5P1e3HwAOstOvV3RrX7+zs8Q70KeobKfMGso0Yvx3mym465FDAUgsHx
0IfabRT4fB1wqLRou8rgi/doXtwymDZ3J49w9Qc13vaOQajJRdtMPATRvVPjY/rf
LZUTYzscaGka1O9uGR3jfy8Z9RPFN3v7GlhAkEJa2bgpWCT+zvun2fuOjQRfRkJ9
7nrv1DOwe0kRz3pFzm9+yy5Qi6kmUFFII+HtjOALuq0j95L1AuvP6JpG28fVHRbs
9Oun1fVPOnhREKvVYPuFeHbrXG0BuydzcPx+XeqhpeuzfblxpE1MSMSKR14NttN3
cFYpV3g9OnAxAN5SDuBhnSZzlunWnu4Ek8HAQqiBOmJ/o9LAGfiaMyk0Lczyj+9z
pFah0OHeKhxziRX96SJi6TUopx9t8S5H2dNNJGo8R5/bIQWgj+gb6qSw5ZNRAdpo
oCnrqgnsNc+ZV6DTXneNg5wJEj/3w/AA+UEIMyueu4Cn6oJbSQ36asG7v6VeLa0M
fFtATPQXHP0Ykw0NOPVwAzm+M78mTY8uoJCLtnrydJR8vvTIu0kp9WELQKIk1kDC
3qdx5Ev/R0AoO2rNDaFh7P5giCYgnHY6MTXdgjxRmvK7MPJGibYqtcIkpgGt9Nrj
CyaixS69WKFp+reCheGyTHoAmsJIwtsoijx7IfoQGLlnr0F/os305HbFkYlgEiJy
1ZJKIfRAhU1R0bVUY8t+X6Doa8h9RLqSAan/qeVX5wfXvHYAeur7gYr827Zcf5Tb
ibHzmR5UGJQwW0vSqYvStIgi4t1ydNPaVYSLdTrn4T/P9qCz6QT98KOjyhT6+XNx
rs3nWQe/GDc5W0huhNwCnobPZgR7oFBQ3A+nx5ImqtTnFIOl+Q626aWrPlTfRclw
3/G7fvjWjPvZbPkRraoIk7z1cGZ8sPeVRBhOIwqiZIIPiduhuCf5GkuxGsEBarbW
100xlh6mIHLof2Tmbu2xTbwSLZAsUljwTey/Y5YYyweVZkfRXKFdw2vNnt5bOPZz
yIJTtT5MW7sY6dW2aUCa4KX5nLcsUVgFEiiKj8+8RxU0GwRVVkTMHsm0HtVkwIu9
nhI5zQg+VnIXdW9BkFlnKxPMcuAD8BjMHJI7fRkpM4KyEItWgR73wj3WibPlMomj
q1AGA1PQ4Gku80Vx/XcFbpjsQAhqZ/qVSH2GZo+wb5QBZz3ot8nq8roh3c7jchys
4aBL0qkYcFnEwrnLJH0MdiVzcJmn885qbv/NpKtDVHCiFrENZDqHyI8RRFWXDLRf
Rgv8FokHYFBTHnwAfirZmDfzp6EhLsia8zpe34PLX2Puso0zL4RNxESduHVL8wEH
jwVwzYsWBtdRZjOQmBzNLO1vu6fdkq8jhQyieiglERo19CPvloUErZLZt5FCLjig
UKRu1UYvFczCoy9virUN0yAXh8p8gFTLy6w9Xenw8lX4e67FtzfzNzNCwasBL1iq
pqJtxz2aorS3tar6k/hcx5K5IHeePaihV/s771Eku8HoFqB3NbNv6bsxWvIrTwIw
eP91bSIV12o+opUXQPDQxmh0zUjxK66ZRQA/YB5vu5txxtXgZfBpT7nUQEFKKGhx
XSfn5u1Gcn6tLpXE1gE4xozmeUA61CX8jgSDsmToAQKatS/BohjTJiFaC6Sfp+UB
DTG4hblulBEtfHTW5+aeWowHgyt5nAo1IHVAtZXXXnsniPHqOCeUGqf/KBkD/bAU
vsuAwxyzzuTbZNMuHwIdnSZcSC91GUHUZ/QnF2xmAjR4uEyJgmsa4gnJZPr7TBzW
v1eospDbCjroXR2FuiXUaWFeBriMUdjJ+DX9Mug8i3O3izwDK4WXgY8mLENvrrzA
M5Ufzx2gZY7v6tztlqKgOJEkeoqc7YBXBheFM5PrbfRJQWa5+Y61FMK41LqDPZCQ
DEJDQc6GdTOIeDq1W/3CT4/oSsSt/aZHSLKBV4FVEwhLhNmGYzWmOAfIm6a+8G3w
CTUCUAOEU5kp+CYJANUVQcu34zKNg+j1sXYS0lwSytPkZkOHoYSgKZzs8lVNxYPj
zkaigX86aB/fImjdjJqKi81TZUlSP5DZ5Jr6TlCAjrQKKieE+Nul0vW2DmGoqCRn
E2J3LWIQ6G1gtP/drwDmsJr6eQfVQw4lVLo0p2/47Y/euZ2ApXB8HfVxTv8QmMmh
Tx1LUZjFLuzseN4va8VmqiyVoEuQPOIlzSwiNrLJUtwOcF2oVVNwfMwdKCoLVMYh
yx+glNQJI12gJc/pT5tULNDIWYdq1aQG50GT6vUpGh34c0yhLOngiNCp7yihvOhg
wdWpAbCQZTo+/A4crJbzrS+GheSnUi12I/nbA8J+m/zp2i0AmsFj2/G+L0Y92Zht
mufyJMa+a+p4PfB4O383YgBWGevHFXsbQyD1EM9v9Wr7QxTg7CgJi83lMOZXcXho
yEb54LBrwHyEn9j7rGVhSvQKpR400Rf34oJtN8KXqdu7bkqmRzFjQFaqY1YW03fz
rTZWVkpLpHdU/+hVi44pqYOWSBrd2mrtebtoGfRz2Kno060FVT/L0iONxX6mAEnp
6iLkXRhDNYo6LOp6y6W+NqRUgrnq9K7x9OjiukmN67wkGpRT0/X89WxJINwj8HCV
ky0JiQgUm3kIAFawzTazWis7Wfm4DFdJB0QJO+onyobZXuFDJyxJ/NbqExtB9PTC
uM56pqEIbhztunMqvOQlH53JjZKjvqqucBnOHumA21C9/VQKecTegaZ3ng39GxnF
0MQgJxEiucNSNiHm9c/zdBtK99p1wXbCfAMZYq+/sRNxSXBq6/zoLJOTjbp2dxsh
h6iQtGDVHY30bR4GAKfqa0uN35oGEAPbk4EihsU+iL7JiIqetYzgE9rTW+LCla1X
POXX4eFbwwIERwQeqE3NdK4QRmMJ72b6OAc01FC9fBzYDzTPqcAVLAuInr4948co
v/UBkwHm+gZpikaI9J6kljtDdfEvjhml5muIXjBqolPv0lNnJJkvtDZAwimicf1X
azPRBqIfz1/uQeqnOyByuyg21tM+ycb+r1x3a+bmzqAivbUPpa+KN3xzqul92iPE
+1RYwxyFgyOxMIXwq7nel0S+fsfY16XBCUBVMYHxSpYk85Tm/12h0kt+q4UJ8fAh
I2aSo/RzSLX7iflmyH+lFqP6thgCVP815dw7HlnD+3BMMv37ugCGYfJdb59jaLTr
pGbhhgl3TKrupdWlOzX2Ey+LPqvQe+pISH18D4FQUJh5jfJVOmH1zJbFdjYuEA1T
UTjy6UTXudqKx7bXn9rcWNHTiiFLGHeexKvzF2qS7j9YYVsTyBVRJhbTIdxqy8ac
IxhCG9MtxgdZV0jOD2+NP3NnOeEl7R0eaRrw2EJcoGz9YT8glBVhUlciZ5pJlHGP
73oPmm+IkEo0pfOq1O+uwTTBjgva1uWGym+o8cO26yHSFLPwEm1wxqmoHNWyQEn8
Ti+X9KXnk3EMCDln1oJ/eeY0BTz3u5v6yuUM2IyK/3mPI995uirbSYTyUV5+mN1N
rTg442fddJSLERBISo2DEBgu+z8rnqLsgee/LrHjZU1RDjYRGG00vBBIjn7O4g8W
tAvvGrlKRekasZntNKIeS6kp0jH08Xaz3bcXdgch69LLPtnahR6zueIgL+WqKkEp
fLFRTuOWzoqsH8um1SCHF/jQxkBdvXgfv46gC74Qp8l2qimiStl5/kkhdNvjjX1V
Hwn6/FTm7y0WPnF7qmzQBFzO/DDHlzNRDoFASXn+56M/54DZdfIWeHL5JsLfYUI0
ZfWeOhgc/VeDvql6xvJOIHUl9mC4SrmKAFLluiE2jZAHR+4hEllsAi7lAgopQ8rC
peaIx7aQTZZyW3R/A6FyQH02CxDQRDCH1mfD74WTQTSronRMw0O95KgZSi7eNggV
rFxMBY8yN3DcT7jWhv+2WJhs4clmBA/kdLf8HeSRw9pNrvu33Uk6MOAnPmOchGY6
98Y7a6ixGcrQ7+hwUN5Iv5P5CQRjaglWjfY/bAQMNziVWHSJp7q/DW86HJ0xdE7Y
z1a7u1Nbg7TgMgPGWx2fPjfefr2vFgVbkuyPTU2m9e6pKu5+l2z3bl9f0OgOa6kS
BcuIix5B+8VqSUD1mvITngpX2zQKx2PwYXLGdySQGz27ntETmLxFlQFgRN4NLoAl
pzGUIdiKVGCgvImI8yFUxHJen4vCSWFbgoHvBNWUmbmT6RvsD4JOWaXhtOZEFt6p
nHTZM9flnZS3BMwKYEZR1Rg03044E9qFqW1qmpJnNsk7PqNZmR80RhYcdhg13YzU
IBBws1DoPaRGC/uSZnNBrsU1CxvYi36b7uqC6qjvLWDwE2l7MQOPdKOnzow69AX6
1UNcIHq+HmirJWVFzPjXBQOwfrgXpaN8R9Q0g2WSp2nE0XMKFZwq+hsVFc0pHKBi
ayTfKLK/puzauEMOiJglDOc4yaHZWRnQF9UjE5n7EMTEJ6E8Qvl0wurlsyzRGjGO
ZrBwKekvErGeXLL65oMd5AwE3Ph+/qkF4QK9wYF+cOVTXTPO89BnytFQfBWd55u/
j1/XsfI+Si/Hueyxoih9lv/ijyDX9OFnS0jiYkoWOgo3Uw042fZddhMXTUC3Ypn9
TReT2C22aPHx7k9TIsWpwLzhpQ5ba8PYsWFAn0opxYeKSbfax1iASX42f1xHastB
B2yQY6naGPe/RGmCfgvzUWI2F4nvQA8gVpTBYgBe9Z/DcJ9fXmmX/SjtNm208VuC
l67+lwo+hTTE3cAgkvHARx5lB/cgyAX3bKDab+g/rjkDIZnlg1xK2dOJZa1OyxME
7p+wwJRUZEEU9S69OAfH2+eyyZrejt68mv5WvVMXs7EqHQW+S3TiPLaKqevWmmSH
mYWr8YCzYEKAPHzmRZBgIQBfGMaUNMe+Pm4PL9k4AjlZHDwJUo44S9d0VAAIy8TE
1Th/OrYFjxQmvMaHnWk+5X7555qRvtVlC0jpNXulaHyZLXpkbHx0P9bw0Aq7KjDH
HZq65PfbA2hko/74XH7VvY9urNGCwJcYk/f+zHPkqHKkKxXqWzfRqd6RA737VAyP
MBsIZIP/2kMTvM/wvjLoDd7QYMynfL0OeoDSc3bHJRcnTHaSwIBc5sIwQiml0BQM
AjcNNZhZGdrxfxvgyVopydX4x/qoqW4tgriRL+m1cb73dw8fmDyWkwAUFHdHyld2
q+bLKdGylxkdk4JWmQtsjmw/g+RTl1phsWs4ooKTJfHfo+X6lHQwkJp9SFEJd4vZ
94eus3GoRiQwH5ZXwd6Tunj494MtCdGPO9QT+FiXUuE0F5LGjWgXFPPn3MKNCXn/
zn2N1u2S7pOelKMUpsmVQhnp2TbfZ79Av/E0Hu7IrTvVQvGab3znldIpUVTPUzdb
yt6eCL2eVV2zYzcK0gp1lFfkrwz3UjcetkAHVD73hHza7sudvPD1ks9jc3ppzjkj
uYIO2ZsvvS7akQRc4q1Nw+wwRHQ2iZfhIuwVTqDsp4XA6IklY/HB8VP32+3GDfi6
lwoasLSmKfZFaxJbz5yxyn6HXgfizPRAe+1j/P5bHBu2w2e4a55VdP5h1tXficUH
8mR+tHyT6r7Ej9qy1DsXftG/oSOrGqjEYoRY4BkYAHs7XJau/poBVHsGhNDbBllg
ryf3ilQ+fkJnCe+ethi2TFQYrMyd9sqxNIs6Nc7LLMXnK3VAiyT1J/Zt8E7urEl0
5t2AmrV9DO3MQW7qQUPTulPeM4SrzcNRwHJ+FA0DueSlRor6X0OmblqTMZqkbGyx
cH52SABxETrdORmwkt/jjZRSu14cEc/VByWIK0oHrI8ujHEh8pvkdkuvI5BrUuyt
VFMSoet7VLrZzw0F6OgGBmrckhFSOCIYBtgwdK+3/2ll17Lo2V3RzMYx5LpN8oSR
YrWIfMMa10a+C2s1NqmR2DyN4WkJPN0eEPzF9KAaHdTxdNS7AmW9FjqnwEtEqUPK
Y7MoIn7dSyCioWwBKDSeW/YtLVrnX20nF08UWQEVlTgutvu7QMVFORvw0owVje18
n9kw5amzQrzJkwFX8BACJalTQ1lTrzh9K/4vv+tYYmhYmZZ2OwYRsEqtNsyXqY7/
hO8zrstKzRdVRD3Am4B68FK3kV9Lv6PF0UHfrkuqWfEU/GBI70lXj4miMkUcqAL9
+3pHHsk6g05eC2QBW3QXd6FSIP+22Kz4+mbclAalPIBpKhgAPSg5nx9YeZpV0Jot
oxySQPUBTEkLe2FQKJyLSQEnB7gHVjCSyIMKm/MVD7RBNh2vC1TR3AWJ3ddrWSSc
8ufxyE2hgpUQLA6iQLTQvYHC6fgkTIH5/cbAo1GMo5+ovtleJV/9d5r5df/Hu/7Z
P5OsdTCSeF0KBGnlTzMX0CP4oAkVYMnYCDugAIvzaYu8UyDF5EWUYLZvLSwpcNzo
POblU7qTSjR0quU0uHZoT48dGwkFkZmCzZwTRGH8dk5o3gEKhfbB0hp4qkNKUzeu
bihWt9VPiCWTPBGe7wBCnXblUMEuYPJwqzg4srBdLVzJowlxC/wFHdKW8QyV4fwh
M4e+keafIZkCgYkX5aQjx8vPqMUIiZK1ARyuNbiXlGBdRA+zkGAjWuFP/5rtNLlZ
19u0F7VEmSHqlCYtYWDEabdPHroylo7qR+ZwRFC/MRN12ZGqgx/Kvy6xGmNEA86L
jxXIPdztMY+Qg33cDzZderyhMm1QSztlAlW4f0C0tAMe2gIdPHQpj08YCtP+ftBe
kjxHvVZcf2SFxNWnLbqI/nW8G+RG2H6jehN/ebXx/drZxlWfNsCLiw2RLQElJCTB
V4jXJ+8uGUTUB63y19dRVCmAj55mcSQamgZbp46OMRtLkSqN2sRhInt6UBpuwKS6
P0j/m52DuIGzdwr0sK2uZ3KisH9YiaUfKQO3VqvOFB1/dV2mX7sSjVcZTzPPUmui
T6SGkrgbObhdBVscgfsgXBUl9BWQVdILVT3gKkAI9wSMR/ZjM/ifrG1cWPiIgCTw
vz3fNa4iIoH3wQwhADIlToMqbYj/p2gstwn3FsNkz951kSR2NX3trfeWvfn+HZy1
aR1n0DN7mPbpy/+whSNbhcR982LZ9Rj98w2+34K/z6G2vR6g/nFv4FERxtNbM9JN
WpDiC/EFtgbwayFq+mH0kO9/4Wg7TEltgL7YrRFUthQDE80jYqyElEuA0+JF3qp3
sdPHAvVB5DO991lxlEVfafZl4wQE6jmvtBA68IANu7Sz/VnkVGojaXYLzpOEqg4M
slGJbtrP6gJ3GURxxTwWq61dzSdfqC+HLv/06fve2HS2kfAJNBg9AXXsfrCERLlk
XaQTlyUA5jkdmvTbqUAfQcYQbUpU1sblewU3+hI5kl0Xab/fz8NygR7i5xrhKMEA
2krRMFXqZ+cbVJwH1KZghAkLBwfiHfz14euhGqDNFU6bcaKWimnbOSl5xYoGVh9u
ZSVK1Je9URmk3RAURFgkaCRTKuDqu52BcdoQLyTXkUuqeBF9n9NhpljvAVFzUO7o
JgsJC1Fl4pEwgSj9g0/N/6DGDeKwa4iT8SX+tVrCUqnnEnINjWsuPe1Zl8262aRI
h6Jo6fVWHqSoOzidFuKIuhndrgUsKlAvk8mPJ8qSgexNGVVjMhA1KaMRQOHRv4y2
+tzpIhunySy6NljSBRfJ5r9NBKDhiK4bVouIcXe1XnygkHUH05YyZHZIXv6+237k
AM/gtU+IWa0p8jseDzKPv/d2a8ZJAZJ/tPi+ohDdaes5myFZEFkSkfk+NjZJZgXn
i33FtUXpye2w6GNBxKpqiuHHlqPkl12eAV8pXA5DbGOfbYwuRRV/Rhl0O5Sft6bP
irlI2XtTW3RpUGkDH0uwUaYtI0rbVx26bsrOpflUtyq+sc8qRMeBSPcS7pB2wbRx
F+a5wxJ56L88gQzmXJ0qQmsZ43tjOw60I9wkoYXxkCvz7jOLpfvWYu7seCLdKG60
WvGeXfkK/zSCN2EmKqL1Mk+V9Z5J5gwlOGUGgl/TshRK5Crx+ott5y/Lnf32Dksw
huUzyixtCXwawJt7x1WDkBiESVIy1m6BR3oExJ1lVJ2Wmgud60uFEQphfo13FkKi
1mMsFhvTX8FLJPlqG3DEsx6mJ2qS6/R0Dd/tcz8cRGBwPc+FkCLFkASvFujjteUU
mokMOSIFl+TvvQs9eGGAH80Hn4REmmObic5rJmPg/1caybVAw/flCJJsyhsnQIxh
7010BKcx1LD/DsGdDIdjC3NQPl8EYWx3xVEwFHwqOLCC8Gt5/tgRqEUcdIgdFTTh
2h7pq0Q+RUX59s0bSXEgSYCdJVW9SQoxhiSO2h2fQA3alI1LMPpKLNqySkR6TiRr
m7WvOsf0VkK06zQiozAHNExZsNL8z9DbWCRCkuKPoAfIDXxGsJ2LHgWmtnhZ31f9
zG5Dc9UzVo5C1xIQ+1pHPEWr+whxHMcGiuAjc56E86sMAohLbpCM9duYpdFlx5QX
i/CaMO6PROxmn6HLX8veVzOttulhANuWov2dTF30A3igB51/IiCxoOf3ecX9rvwA
r+eQpSkw8rb0FYMRhTCwOgPefj5AvS1sw8RkL0hw5PXuJB62N083DxvEDf+6iora
sfkLUkHQU993LnWs3SOT6+s1g/FlUQM8KoMTh1N4jilDZ0T/J5XQJiIMzw92wqqQ
C/pIpA1Ef5zn513bkyWLfiB5OPN/PN7bU1kzAjvaXUZPsrC7fYlXJbmhXeNrAbpi
OA1qz1Jj9hGxzHpaKsqvzRsAU510kjoPM+p4xDE+ZbSQxEqyWeM/GzaRKxXybFc1
sgVioXONv7vBPaxi/v9ayu+X9eJQgQ0Ti3PCWZNw6txVi2Kq0/O+4nlR1wuui9Pc
gucCwsZRGtlzIVpahcMOrxL/OEQ1vs1gTAnt8pw/PCTEI1CSP2diysaVl5lXV/dN
/r3+eClhRWX6D4u5WUrANkrVI+6DsAqS0ZRofj2IPmdxpnPNGokLt50/CD7bVln/
/nxs1OvP2I7Hd3/U8Xpg09hYZIt/u11A7d/OLc7SqhRCus7bMPLaMTlykqiEmp5U
C5brVVSrP8WvoB/wLHYp6u72Nhk2t6Sf9CSeBdtcd6agZVMwNVaO8dzev7nxM3ZF
Tn2MSbYnJWP7YvcIhJ5N6/QhloukXOAvITICb2BydZnFN5Tyk5rJcaw9Qb6N3XQ2
mQAmqdqR0/Mv1yjxiTFTNnm+I5J1+JtCQUYXsFc0dQ4iaqzLb0/AZSidBfJq4YSw
H21Ytplmxbbr6bFQoVonVtNDEAqb96mvKdeVJnyEhhOLUEvWA0Up50zVtZct2Z49
/wN3++42INCPrJxxMIo0zw+35BQCxDG46i+TjBMvr5MVmzMyPqwpLxZt6L6M4yJu
SBogJvOrYO5JlnSofpPJ52GC1CzKjit6Z+pN37EVPnxbsaGyfBMD3Hy7djuCqfsn
WlNCNeB9LrzOf8V2XquL2zl2BbbSa86putlQRUPAW/uwkbTCST/1F7OtTKjEbdM3
dKbNVh8YCxQR7ThFGJA0Dq1yimvzLcdKqsMaYUS8jBDK3Msv4pphlOT36ZL34LN2
Asl8VWsG5C1L5NdUbI5HfcgFVTkKVBF2n8SgVse9yO2d7xs/dZZFOSi2nyMIr36J
fRJky4gchhI48bO+MlZONC1a7ocymnOtInPVGTEl0WIAs0UXmJWJtdaweamHmk6V
FH5NckF9c6YUAQ1LkRaWfOQm26Y+aHNXfUG/s1odJ11ehoC6i3oKL7HqgzL4++NJ
IstvmmEu8mYsluKFqt7qB0IC9g7PZrWAhWQ9HB5FIj/Qra2tMwc49ClwqxogqPkJ
psACTcI8jCM6UupMRAe9J0zonUZIKY0FEYhg4//+TztnEsqiXeMHRWUWHjIWNpNi
7ZJSKEd9AhHp4hAS61WACX6YP7QC34Zp6+Kxf52DN6c3olRcG/UQttRxZ2BxIyl8
EUXLMQ5MY+yRUGJ8CID29rYGlJP2yfJPzdG79yQ+Kc9qvMY+GNou4vPNFxWcnvPF
7nQyE/+WzBF3FCfGfraHpM9kKZ4951R8LTYhQhpGBHgTqyCzK8VULPFMtWj+E43e
4+2eL+UNwXsl484rK2XHWJ+8OadFZHzX1OeNqea+E/mK08coXAoze5Tu93aMoZYg
TwoQpUE1imbIr79y2Blh525NPp2EuQ6q3gEPSsrY4j6cELC1FluEDkEbj4FuIfdo
KG/FzqyDtmyBHfj0jKA6ttwcawE4DEjdoQ8D2nX8ySDd4iSPz6I6x32U0c76+SB5
F+CHwt183CZhBpsg58cX2q9PN8IMIPGZXdFWNWbnwIN7s4VFsiwcryJ7ArAHJbyE
Q22cpx7nmxNRrOCY9c/QUubXjw4wDKSfN2NNm1qDB/BNQpbBuG5KFN4PiT/Hii2E
/uWqc0bJ9ubpIyRJ+5R4oiXNeL2uujpSEGNl9atsuFmPrGS/2wpZpSBJI2K5p0cu
5+b4laMltOSV25AVc8EkTIuuM8KKTfovqMuWEXALeb+IM+TRFD61s0Az+fWXFr26
U9cvDJcXYUHwr62Zs5LM5vNva3Z9HbW9inD1usY31i5uC7K91hz8ZutPqpUwvJic
vBi7TEoBl1SagzJhnBF9K/6EobUPTpCoMtQ83EyJknVGwUy1yC5K1oUooKSFiXot
/nFXcufU+KgRzn9GCXEqVLc3TfBYvLxnGjb1lzz1J/p9JmEugLEMiDgt8yR2z5vF
+Vvnh2mtbIQkPBN/5h4IUPx9OpQ9W/xo6O9CEYjekVaYts+soqPeUOUjjqkVv4yz
Vxp10b5kUt5D+f73nqCgDLj/4+8OHhHj2DtHqu7ZZFDK5derFaQmVm0b3k5jRQNr
a2egRG/HBcfBU4j5x5exVBQuu6GTg1IE7XFoxIhoGfDSWNIJBgn8pJBa5dzlu9X5
/eVKHvobW4ikr9dzcINQakbznPKX0gUSj1mg3mhkX1k7g/uo9hESh1LmnWrq2nIj
OrlJ3jWlHJkcziO76oO2PecgqZuGoqpQulq7fsR7IKaerVA4TBj2uBGW9IpiTKFI
6wcG/+Iv6/bR67NMGo6r+/brLnSgsmxGQ2zRIi7OYhmGApCAEmuNIu4kHS6z0ohQ
1yTk+BFYU1W7UAI1He/yaLXndI8qwzSAJPHbAZMnAJ0lGEytplip/Sq+Exh3YC/5
wSxnl3Gzj2TKBBIbHKXOuOxZ+XxPFFzoSCzwJWTm+5K/j2JN+HE6N5LrvyRKQciz
AWUd6L2OqGihxg7OdGJqKAH4pLh6nK9VCosPTNic8/lqS8nBdvteHWEdN/afV3NN
M2sb+ua8XuiXimp3CRsKoobnfBXA3r9AVNCuHlMePjW24Ui76hVqLRmWpo3lUpEz
Hc06xletKLD9CKOFfGCvvJnP+uuARShsPxtgfSiOGVz4/EOjOfMmpMRtADI9ehBk
zl0urhUn0xdhxAwtwezSzOvRglAKP1afpdF+rEOMj4rEbSTwUg5Hth8C6oF5qta2
JHpM1nqQmAf8NuNOQCnms/QMIwifAZFYN9m0cCIzrRRpEXDEYpOYZKe0EtAhrS7N
ovFMMsdZX5tMuxjWsbRMOIHHgbEKDPBMMaBlKx+41xrNsyUVD8rXbqQxfS976EQN
0uOlxzHjVDSLQXHPpgWH1UsiCN/GeIGYK9UZdsnI6xFGFIbr62NPu+F1MiNGZG1v
P+ef0T3Lr83JwmS9q0q21rXLvx7EsoMdH/UibKfQ/wT3/msd8c+oCH0NHP/4IPeI
zon3z0CLzxJ1rx8VtwuyLMlzhw80oZhiGh6kPNO7ie1fONeH0JDCWmwERDSSYERm
O+g/7VjkA4qOLOJff+OswNr49n+6jDj1yj1dt2H4ABlPUIjDxNz7gl30M4g/upyC
okd3so+0HwNQibJ2Tbk6D2HtAUVsIMVf8Cr3XjJdJOMKhlN/TcCjhW+Pz7GUwXBA
AiAZyczh2SFnMBUzFXOQIunGthQORDYbMej7wL8uz7sMyec+ch/1XhFZGki0G2Np
GP/q/ZwYImEpoiCK2vESzgrLewtiMbJ/ChZMFflZ1d0+NRnKIBg5nur59QqOrkbg
FXcQuedBpxIoZVAaaX1z8NKKbFZ6ysyoeJYJqZMUHudf0tWZ14IuC0QTK4Z9FnV0
2UzU1VcuG1fPAIqtcklZlizYFHlpMSCHYs0G3DMtkbdY3Ud5TVX6kbnpPQxrGOFb
7y5hcAWSptJTVUD5W3JBcmcRqWf6VeyKRva1dVKr7+8WowpNZcBGyHnYd4nLuxkQ
clF4ZaBdizzyTMsDoGAPxzwCOAaPEXylvGPiPw3mEHc6mgvpOPMJNEaPMwHqEja/
xsDNcALrvoKKaODsQZR1y1QvUHadkFM437IujthIW/R6R3uJYCZw+X1ZAkEA5pix
olxiskeChB8aKOma5msvW/rS2cRJeza+afjpxttVA08ghUfO7q7gDB4I+xv3TWJF
EEmiuSBwfEGTa8FeR02e7Zj9S5wA99spe9Hq03XqfkVaW6F+ETb77p3RBp8mA/aq
GmLGKnNe549QluN2UzrU97rULgx4PZoC0yMTKi+mKGFakw/Ls61Ac16E1Ap43eFJ
d/3y10h6pJODHmw+Febt4EpVnAyo+yj5YPGz9f5JS7ltsavwctsVKBqkF2G8Anqo
M99UpI5/M0mZJAbWMXMEcJvgO3PsUp8mZ6a3/9adSNgqv79AHgdS+37msJxliIxx
cKW7i0Ax4zwhUuwOJSEN51Hu2FhmBALMWaX5iURzwgL+Q4Ef51/i1lCpyrjgyVli
WBSqhM7C0cpgDjM/TEgmbN49B0ap+oGXrrNZ7kbi+laCa9fRMccGpidPcbQoHqXH
hyj0GtYc866hOmpx5nYm378ruNJOTFt5TV3LJfliFmFwC19zBg/24amOb4kztnoo
SulBY757PGepHpid+RUtOnCBMeJJtKfHkVkJxigLX4NVP6P38HaurUS0+khM+J9b
1H3D4KzYoXC9+oKJhpzGUyMsRORQ4tRcWAkSHhJA5iT5eafIIdNuK775/ccN4ofG
K5luvLLUfKWRfL4gnp3laMDj8yx2g4EzMaELuJEPFU2V/6M7ESNAehtPdheCAopu
oppSfBVX5sBlCp+CqLSz0+T6En5m+eDyB6n1ypKnnxd+GgSAwfnn/AaltTDwJHDK
RSBz1wtQWrYW/wfYR9rSTyQZBAZ09g6FwhWdD2Ecf0ag1+4RzfvyTQK1yyeMCHZp
09GH+d+WqcGO6j6RayP5PfOreatw/hH+H84vOahjf9WUNNdGyK6dohoxJBSDtYfT
eAiDaSvA/gqOzAZc6bdgpp8S2qI7f5LW6KwrSj4ML5ZE1N2Ik1DFL8FSJNibWTYB
ujnFk90uynikK7uPPqvdti87H4nWfmBH35iqh8ZoYaPrmcr+YHbCjPQChufR7Wcw
lfEhYLPRo3/+d1V2XksN/lHWLbCxSrOZebw38ydAH0LNaUTFXh2qH4uZz3zmUrJz
7+8fT/9HJE26/g7vDP4OlvSxC5JKJKUyzkrF3nDHlqdyV2pQREKE27je7Wdfl4Yq
6I7F+X7NDswL52M5CYQ6JUogxt4UMMwg+ZnepQQOp8AZ0rosfvryF9doRU+cHIvq
A8jGQ+6tkTkIJ2Fr8GpahXdezkZP8EUg4y+/dCpw/JEUXiCox6PVfyVFom04jrh6
h3dC/dfdevNkLzeG1NRjGO0w5bJGBNNuHr8ENIAy54OcsVkvdZKQ0ZmyMePCRSbo
t652XqjJyn3J5f1YeaaGvWm9dK0bgsgNqeE1BUCyXUZF4qUSEOQN7/T5JYejhTJR
cAbYTqEbQi+ICjPdmJpOh8Jl6aUJARNuLmeOWaGaNZ5PCgKxQKNaU4DFJRfeUyQS
rPsXcgLHCfyufr81ygC1Oqi9azNiiXuWedl2ytsSN804rXv2BN4TZ2zANtXsFQJi
URuuiV+LdHLCQwaGN5Gkqf9udr14+2za+Mw0ngtaAGyQMxSenP9jE94dWxKF/KPq
YwTDvzu7lfnzNDYngMKycLiulm7/dLQRgyr1KZeBXoGc/Xh7ks6v4YpRyqQWncmU
haL0hmEzS1NzXDItd1KKMs1xRiQbDxQVwLczDrK5Ufb0sTNieNjx9on4chknQEQf
VcRBzV927jhwSJqqzehzFUcMydvZcxgOl0Sc5CNWE26gSQeAwoXyLeUR/GEwDVOg
faMTZjjyA4x9hbN7kgZMI3QAcyfQRXzswUmqVgBbOstbbZkihTHJd3kD3PLs+7X2
7MqwZqz8EnFtonUucV3sTu6PzBvYyYzDSnu/P5R0DrhFi31b9yDxiYXBQjIC+XDW
LM7D8TZix+bTvGnX5DKNoWE8zlwbCwQX04yAaA+2NouL7RW9SAg+G2mO6kQNH3l1
shPazgAhhGmzFYaDKvP9Lkw8BTiig6cRqjpjMSIueigO4BWxhz3QChq2vTgBTmrL
JM2nndEVKvamYI92Jc6hBwPwoH7YkxIQttfNP/vO6KU5LZ/TKm5fo6l2qBKZTQTE
ZhKKzUsWo4HiF4w0p/Fd96mqNZEbFfrPwHE5ceGGQTiOPncsn507F9UXKRdZtKBx
4gvGxqs/kKdvs2JWtL14V08hre4EfNFC0s0sd1yHzLma0OmsCN2QHmKwvk7hjk0F
UT4K787jLOowPKBAUe8UmWZnOBHMuCSrzPzUvAM6yULmRNchNN1QKNt6fLJVFl9O
OBC0VO3/TjVGNx/HAqKOJ8WWIxMwoBkgoc9xDNYhyOQoiX36VVZPwEw786ioq0k5
fS+fUlloAiqD/4hOFLkHrstJER4vkpGDByznhu5XKJ7FyalvLxnKDYOB+6+xZ33k
Lz0fNZIbXcI2ltHI/DaIfBEhCkWrOTe8KOqrSPY6qHdQzUevaV8lNRA5UQsgW1TC
UbfmaGFKfKq4rqYZSPLivpRNGH4x+BOaWTtGMhZlDP2fiBaDBwzqhtyuYuOwvaRl
vBiJLJ7wT4VLnjB2JvEO0Z43iM5qmoe5uuY0FE5PVDgyqvH6z943qpzFtT9npnnK
MZpLzXK9faYR6eRQaXmt1ckdgKmsj9REXRGApiBZfV3YARYNr0FjhGRIjjCbA655
X0rNXOsPMRkpNM77tsKfdStzsped4CCvD3XhvAioRFA/+DE4U9Tj0bhWoCTsDG0C
pKnB8s4bKt0TQmIB0jlPzyM/wmxJtc/mvJW67+X+2Ve3LTcvDg+mFznmyuxrORh3
faKK98xVUOBzqkJ1tlNK9m/WopDIuax4QeOzj7pM57QfBordOSay2rBNEuzJLThT
X5LfBbHJrPzk3/lc8fd9bfijkMQxGY/tEY9v+9oBB88pxndrJKrnedj66ZYAbcgE
YYB2SeWrAsUssKLAD6RIeyH+QuWFWdx1Suvi2EUxCFOtpMtWEczDW+81pAQnBlwN
tLjCCYUjLO3DEDSCz4/2MnKF5cmH5VKQV5LTs5A6i1z7j5WDBZ51lPVFgdbGyr2L
mRo4Cajm/mXyHnJaS9PDSu/Uk3ssFLJ5q8uTil9Bcj7poqyez+nzuCmrATHpSRMl
7QS2GwKTz9x96k3ITgBsap0vNGHJgiaBRm1tMQKCNzGV/eBGqTJg5fFEcJkb9Kpe
QIoV3c8ofEAkDk1oAen0RgicTE+YN0wwXYDiqCzTXa0rEvxfM2+DSTpjLXWKpDYp
GVx1YIsBpcq0yEQKiuYfAItky5tWgFBZ0b0ZY7ZCS6cjzGpLSj4Db8/ojoCLX1xJ
YRxv9bRxkHCM8tsQ5E0aAhTKc6BbIbblDfVnKuaja4mhD52rkvPTtOasQHJHqD5c
fI++rw2QxBbb8wTVMyGJHRraSC7Zru7I4IAnPcuv7w7fLBzEOFPUL/IJ4E2QUEn5
7fcMAfQ2E/RkG3UvXfqDQ7J7EGHKRuzuPl4Ms4p/ik1H06TRzAL1xXRLOvo8Xhxd
b9+7SlABqVbcxgGQJ14LuA+rGa9LuM3kS3GPjOPUC4BzlzPCHIvXy8SHWJVEf947
0ej15Yzl/JqcidOiITfwxz2c+3g4cC7LCKl5mvOpbNDMcbk0bDHbZEN/IFeM9dfA
wqMaJMN+6uSgafIV9ZVoD4srblrvnNzTVxJGwOlwO/ewRzM4IJFaG5YaHKXgf4kM
t/AqaWRzJ8cRE3ylN901qLAfgAm6AZMW5rOAg+PmBluGAGMffAxxz8TGRhwJztnL
cIO+9nZMboo1lj/aTy1XwHwuFLsosIq6snbCdcIjMh3Ad4FYGGi1Bsa/rZCtu7k2
qn4zqrNHhd+khu3pKIFzwNni0iFIIAq7FzUHFwjvONwY7HxwUZhVnnzNk6YWRORk
sclBysVWudvBab12Q6HssURb4J3dPg9neEV60OhI/GWekMRLm4fmiMB2z852kgJN
oP/lt78pAKvo7KNi2B4yUD6BZWtaYDuGRncfmceK8A3/9+vKLrIK+Sr9u8EK7GSy
XygNQM2ftQK9VBjFKSnSUP6xOfUBMzSijjXlFZoNTwyTciSh7DWmDvPwmYDnFbbi
DTt2of5hfmYlBMtRe8EC5bR8Iy7O7cZ+sYAux8YbHe78mBpAf/kyl/SgfPRY5VWm
TXsCaH+yFRgkHq8iHDwbDLzGCgTXrdi2X6m9q/TiiU6CSZj05B88YNnaFp5JrhGa
3eKimFGYD1exthol1AWLhu8CLnKTjJKJIWJTx8AvFrI5xgwmNvNWwXIKwOlE4xir
HHzCH++o2YkOnxG56+U5jMRKsarPdf7cg/JPBQpW1PvQb8PuaZsvjeVF5ZEnAhRx
MSIWK0rHNlQD/uQv0+1ZHCDyxrF/8chTTQLllhtKZRu94UY160ahIIqIk3x1dcwl
0RIQ7tcfNhp1aFpAtvGNeXehjVleYTVR4XFL4BZeVkgyJxhn0i4p09mpbedy4qDI
wb+0VP9sKoalAE8wH/CFWEzyAXIGQhkRu7cgx/6+jxWpp8ZkwLuNbnXv6vXt34Qt
FfBQkHHiRi0u/6p5lULcZNsEulJZVkJ/0HLhKFDXKCA+sZBdZjrrD26RYwShtmHW
uUjjw6daGk9+HZoJYJwLMuaefD/nMgF1zA6eE54yUKHubmflrjNFWtaTaFDs8nhX
esCATj9VHuNzyB+xC+uGqlqa90aqBp2jeqWv7VaKtD54HfxHMUXuSsucIpPv+95q
SHZdPpYoRTvJLZgg7Ubysr1MOhJthpzcWG5qkE3gIxYGgOzx2dmdK11iWqLydo+l
YPVf4l1TAVF3qgyRszMCenUiYysdvGMVVMs6epSQ5FdBfjRCX6KWRGU63WWo7sIU
efwvkbz+K4tV7nh+hs1oSSkcbIgBqGd+URICvZWMsZTMOdKon1sN8RjuNT0eAtQU
2bL4RRceyuP1nkF5K+uSdqbeuG6pb036w+/7ReO/Fm/VQwdp2DAPgScBLAAXqoQ+
0OKVVuCOY9iKrOXj7bF+BSIAXczjB87SJoDCXwqdSgjioUst8VNpL7dyjXB5BWjg
n7GLs2sue0i5b2wD0VtIGtQ2QLz6DPBIy0bnagEBl1kTWFDOXApdYTGmICA4oT1W
wf5vt6zqlpARYOEMhL3gyCZQcQZv0jhuQzoOS6LCKS8Y5NsssTrsqzWU6m+fEgeL
eT95pRmCwWy+MKEQ8FgmdIRZsBWegzMC2Q7Z7I1xmoVsnjJ2llIDZFw9N842Ax0c
xG/GCkibz5gs2OYDZm1XkTxZDmuKnzNydDl0rv2MtnVfdSVQ++onACHUmctai2Wp
Gx9DPGAUjqRXFPxfUdFf81qA0cUPJWO+ZMEXlHriRJR54vKzQ51e5nYAYCT/uCiC
zHZWYy1GQIoTIX8y8do5MLNTQgx02dmAwlsOebRaxduBtgvvpSRqxOnkcTjbg1uL
y8m8UIyn75uaR0qMnaS++cypZgfancAcPFzs/kF9cP2I01PDnK+Avjej/UWeEN+g
B5m31s2COYP2PkcoJaSO03jFyjimiRbGb9YOWYOhRzziNZmKUYMbJtGZV62iOWHE
8zpd0yfgHszzJsQ2nGRQO8MxSa4Rzx3qQo6P2qivLxEHWtoC4izqJDokRtpTCE55
lus7LrCKIChK+W/ceFqXIsaOf15oWq4tqrmqmGZbk92Zs9rAge12rOGWvNOJBeag
MdcQQXmsacH570/sNXxVyGacMUEQC9Ak59H/x8dmUJnPRsRsxtVNHzhx2qWL9P6X
M0FzYW6raCwTc2SFisqRtIKaejcZPPbE+iGrc/ZUcek6BpfVQsYmzvFfbB6WwKcX
dCtP0pQDBuclpRE6sZmG6d3jgcYwUXqswg/PpIalsLHiQDDbdBhusBDpCK9XPU1R
3K6J66Hq9A1fDHDZr+NJonNWniBe11VDw1v8PSAhi1z3sbg6miPLL2rEuLLKqFyA
dpQXuHIZ/6Qg14Gr2gotEOZp5wD1bpvhPAYJePcPyKKfkJKKSEnf+nE9oD8LGzW+
er5ipcJFf1HSsvQZxzI5k7G648wSKHxNBQNBq0hJZPwxt1QrrmWTxlFjNOo+EUMF
UzFv5pFGH/CJcYzilkHw5DcOCdYiprKmByKhPc5nhQD3n6u98NzZG9ffyifbhOIC
FlfcqwhMav7VdLkZ7IBJ2rnN4j2Prh/Weh9sXLCL6g9JiiG172aCcOVCG6kVlKw4
d022/1DRK2HhJjfLPhOuy/RA3t3Vk6GcGcAzMN6udxvice8P4YTeSbxwYuKaS/gu
vqwtNniJLX0PZWW5h1jR6q2x3DkRnUjdestPC1nDx8HHOHW7JPViF/R5QPry0gXy
pboSnHAVyRums7JTwR7gQ4vExyhE54OeqQZ5YUPQm/3NApQN21x01bDnVlvuCnvk
gZYuFalZsxWzbYiqmYaHFhe2Bm8Vx9YePL2GXNn7I+keScMIQfhVMVl+e2Ys2H+H
aJjB8L4VM8eAi1/VriYtRrH1PAibDAdKroOMdBlvvIi0hbHH8z2Rg0jZdZaNunqO
6fEeq7kv7XvZUmgl8TGKz2EiNAmOYzVL2AeXteJVV7gxo/OR0YZSIcrF6MgpZ57M
M+cWtNp6TK1tA2+q49WaBI39pTVvkv2pE9bJ+FbpMK/LimYZCtfIztsFyhJgNRn0
eVRxnpbQI77+zkIvhprfAMqX3ECPBDN/5ihaEmwWovsUWrhK7bOM7oEQopnGag2A
1dwsouEyd0FSigwLvpVPExlNiDJYY03TOd6aGaP/xzoTCLsHMMmrR33bbynAVY2/
dNtjbSyKE9pS5ZOPOJKTzuwNqZIYR+0mIpfBcgQO/KnOsEQOGH9nts8aBWyaIXpp
dhaTa3FwtZN+oI9XebAuJmqOp6oSQxESRmuEsk8Mh2/2oz8zL1PPEl0qW6EUGrpJ
BKK7m2Pcjvm6ZiCQsZ+6JR74Ajda0r52au4NzqAqQFETD25DLLEL1XGAtYCCKHsJ
WdYERGr6/fiNW44GTFP9zjoPREr51bD9yoM8l1itdA4JNF+WresZthxqFL5tnSZg
CouIPORzjH9nciAjsdhASCCW4lG8JaKABEdaN+zcMQqLs3ux1SM2cemtFnMYPkPb
PUHeg2VRvBvVO0tr8SUdJ3KMvqSildC1YL6gQ/ve43zGYAIjov3QhjZT2V5mYoxZ
aJENNkfBHpihvteFPJVDvyudeNCxORYdQuPBHTpnA68jAjREzvs+/z9t4BEl0i5O
iu8az19mGOlh0p72oUYd/yqUmWbcEcYOUbP9iFoCmL/p9DzGfeuEcoxFCyryhykd
2co8pFC8LKEPNu8HJxqjrl0PYKDuZqbta9fWh2zmNhe6EXZ6L8ZsVjDa9MyDZYeh
BuK9dz4lvF4eiCKHc/XMULv3bPG2Y7AWOu3KcbDK4dbAZM5P73ATC9fX2xMJ3haA
pb85DzTw3ZfN3GFt+FOlotimg7nEI9tekMN9UBT4/UdBtLAdYRiFED1cy5cKQJgT
3A3JpOh3wi1R6aS4Dqzkj9Y7JDFa/0R9idTFNjqqV8eHxLopqIbxJou3GIhhm14o
C03hBzYXBILDcRCtZcFQgKnQ6Quxk0Q6LARCbEVVXNivy8KGY2wDQY/3Kid9rhlm
mh5YDZrDZuDzUiqKKFm6IzMryHiLKHq8o/37ghUJjfHus6QvIfUs9i1MyQKTESsA
uCaXJlO1zlbV+4UsIq+WcJBD9ZUpRF7mqXw1Yjw465dXJWZy4CesKKWmw5J1iAeE
tLbCs6+nZoCnI5q+l/F9jKYNmkTnjzCpDJR5tdmhzIcCC2Y5xqXaGRW7hRBn3+Q0
DEIPq3qveyC5LTyPZVDuvDXPvoAsU+pf8qgsz+Fu9utTX/BJgHp20wfks4+qwUc0
UmWwipJeEiMz+WQ2rdvOlyqKA8tobFmvlqAS+uwgCh6n7UHgR+2sOYartda+wZvx
xYQLYVkJCMoQyV1RPXMnhaH3Amkzn2H44KU9l03+oTv7QooSKz+abU4uXkQ19cqq
ujH01Aj/TrzMeIM2DgffvWQBxYS83GNMhrUUevqmGI3fEumXm4cKO8lSqGPB8cNu
igoTYPKYgwAKIrvX3brwym0MxJrBwG1HacderE/lEeylQWyf02SWmncukmUTxugD
MImOEXBA65K813Asdu7iGdSM0P/TjId/MONmezHqL32gVDVVUPB8v70ZfrPQ92d7
SzyPNLOZhxFthvEEBFuuww6ZtLs/Nz8WozcPEbHOnHoQYwdUI4XPni8btEvmCS6a
PCkGwJ9JLjYoTsYtuWX1UcFAeoxBeDOBjCQNuXACNM6NCiPXtqnAv1M+7KR02iah
QIAh5Wf9wW0A0EM3SS11j13ukrCxu0dTXJWkTlAwDBaOuofE/o2JjBTAHpElzmSt
LJSec1wSVs29uAEiyy3TOWEFM5qD0c1bsLm88yBmrO8EKaxWqDlDTNMAvq8q/KIz
lMuZRSfZXuC9dM3CmWhpn8x8smdZEDQc/IOlhpst1vqdkmZ+d3bgORHVU+qfe/rm
645ZskvMJacVW2xt9Nn8SHogFvZSj22NBi/MR9LFMrsWIsgeDKvuz3GkyqY5tmnt
44aOas8y1YjtKHXsJ9QxTU+p7p14dOFozCDjQ8V2fcz/lYu0zXfwLbAFbYrG9Hcb
Qs12zT6X+pCXMuN9GIVSAIhwr+bsON/vYYG5safC/h6Uz+khzHgJvHwQKcBvvwBN
pY7kaRurhM4eTqm+7xc7gyjI/ROMBniR4eBWH6vpn/oB5Gky7KrJ+Xc9XHfg2gp/
G6+6pcJViFjULB/PBt5E+BDgJAYa/2R0mUUhRtzsUuzfJYTK8VV1cvGg0tQ3K4Sk
RSoHOVKx/MhPC5wdrffamKeIGrPdl5zIyGR5cfb0qvKXoK+wCFZEkM4JY3BdgW3W
CWwCvEcAtYc954Q6v73wUIQnn9M+P86YTrFusSXhggioKAfvctSKe6Zs6o0re9Kg
fFfJFAiSNisKEFQh4qk5cbZdiXnYIWcRXc+LVcoFE1nQILiUJ8D5E8WUekkJA6Wk
5rLlsDad21bUVuCXRPkCKuM+EaulNW3SOsrJ5qgV4V2w5qeWw8h1PjuO/My77QHq
iKqqO62GFDNjUoxVDDG/TCRdSCfq5E/GReAWnYIL4nwQbm/QVqxruFU7rkP4w3Il
ntWPtru2yWLI+RsHNdXwcGtXE8/1Fvdi5RLcEJOYMgO5ZHDyNYWtI7oY9VUxgP2D
aDJZXnITI4lNlAYR5HUtQ6OIz7eAOCZU4aJwTFq86dPRxUuNVeO1e2RP3Ee3Y8TF
j8Y8icVFjcn0CUUXaO3z5ATcrajIQhLdU5LTdu57A2wFFTYsrzrdmWa7N7RwdCwt
2bUOJErOalH/SRRGRs5OGSgAgnseElwGJU1RX3i3PYG0V7fQXCVgiBAhS0hqo9Pn
eUYLBV6DAgfi+6NsjCswiFhMwqWJG/cvbmA+3lwI7mFX7+D3EY19DpaaWMEIDve1
ekHLQWs1mfVR0CcrTAV945nveCFO7A9p1qUzRBZfOzeuaOcCMJXqM3cOxcKhVXyQ
rzWeh20tU0Go0asDt5yiigBc9UMJ4fgnaqZNrhJJwm2n+70vUwxtjJb0aNv2klPe
u7gRxNxF9pAJZ4itAj4LggzOBcbs8QaI4TKK3VyMmtnYUV3GJscgALB+F5JyBJ8/
kWYH40jBKCedFOVcPKClQy3gDm11YBDgSeaPfKdNu1jNzOkci72Pd+LSTpH47+Bh
rAm1W1DKKcIkyQ5WnxolRNhLT9psGI9QARI7K8eKOsTIAk6nbBwC5DcV+wve+wCC
OI/KuOp/Y/9CRFidNfF0bUWtC4NNiv6VCPc8y3uaAXa3hXH0rypGEvwsJQ/DmAxH
YnuLTIXmJCEU6wlluX5wp/GCv2LjJ9Pk/lwj7x1QCWe1xKLrfwXm0/xYabysFyyn
gy245bf/SThDDZMmu5aLf+H+7OkkrkmbyaMmAZibMc63JVf79k5NzrW1dRKfXCvC
/vCd/S7AiW8h09bvY80nUFuy8o8yCrV0C8fm9wYqfxeJdnVe8MY7u4pmA6NJvr1B
9smQUPRyBHTzsLlFiFHl5n4hVVHd9DlwcaKMoZfVQEDaxgeeQYQui+MulBWXumys
QbYLCRWUQFmJ0fJ86p2jqjvVM1LVk3DnTTz8eJzt8BrJgm+JuFJgMZf9BLurtj7a
qlhjLmxFGgPwMF7paKo4KIBnYNODEQS0MxWQcPF033sGddJAP38uHIK+Qn5DhXC9
0xbT+uSCd3JLqbHXKCFuDGTh+pBxSVgKEQ5Mz6ykUXZj8R7wFT1E5Wz1hYa+CdtX
qeIB5mLjTyPlvlZtIEItOQHAGJ+hbsgL3p/cWjVttrx0FlKi/s0dxbbS+6LQCIxr
TAWMCJ9gOMi8mkpJwSFJE2Oo30IwcD8tMTx78S2GUuxLLhBTLSASsUJVppobC7wE
qmWvYeIkdj+G9Sox4driXgY6bH75BtcPDhcWhb7wBbG27EmQeHJ6n3CUi4v/iq+d
OywFIoO8Ykn25qeBDkZxKQOWxXq7EvT4qLSbeK00SoC6EfN9/cPPdZpQJbh2KWSa
ZjQGvu8mrvhpwfaZyjWw0+gh+6WEqSeqoGIeiD/fN/3LG7JIBDI+nr9DId3kZwSj
3CzkhaoW6+4nT/FO3+s5iz32IiplpMPp5y75nESHdbtIr4FOg1gWeGwMXB5oGdM+
SleopLv+HEJPVOlqJ3k/DlAOszNHN2r4XWwj7s++ssu128K9ObUnHB6+ofEci4bJ
sJoiaxUwfK4nt0gUhdhE7IQGwMnsv7I+3ZBHm5/C3QS/YKUefZsH6Fcius/6wWIp
cJrnGbZyc4e5W52JHTwJMgFh4NHldzbAOlX1/MayHCLbCT0mtKX/SNXmVE9LvTFE
r4mMiXwZOFCG3qRkZAyr+I6L3lPa4mbV00tnds3eU3V/ujiUd3MwmkqqsrcYDFDC
OsP4GxIYiAe4zTXnldgrrYPCqs98lVZr/aDUl60hpYKOpF03dzKsVOV1UZqQZgcp
rCXWSFToOPOAeJ/C9QFQYutvn/xjyg4MiCQ5m9p07hVmCpzDQOTJ6GJ74pUmrVRn
fldtSMx+rxo4aoTHeXn+Kk6auIs86QvFRrcrxrxmGzyGyb/dFuM9IjNKp7PTVobX
YwgZTOwLsnAfLt3iIpP84ADz2BALJE27M8jm5JQbc31/Xkl8sBEK3rSTnbu9BIxW
bHcpPdgCFQHiHAE0Cv6Z3/nf8X1QUb5ZTES/BY2LirLAwMKxiFC3uAZw7WlsbeYm
8Sk6IXQUzF+YI8nwAo/kUzuhIyRyZnPstxgXZ9JxdigpHmUoMlivb/m+xAskq9BM
I9XQNgR+d9PoP00RpXO4V/yaU8LiJTmOWuBmvhwfmhV3UM+IrwIxe1lT3hb/mZGg
r9lGXrCUKU1hbgwYKR2YhAUa4sby/5vFaoj///Ride7FHRYEfeYR3cRHy+Pd+lH+
hvDhvoqGWqlmKFDYdgUbub39aA0+N9HL59ufCt8CL3PKihOwsJXQMLv359HNe5bQ
BSvJTU/DGXkENcFhq6k2NsoCYSrhxxZuXhPb4JDx369fBQVnTsHXy18sQZvtGdQw
LqNWJjIYqzkxXUja1tnRGcboG0i9feAv1KbQSPCBzHfEb/mT3RHP4MuNKnegrk6P
Y+w/Tu/hl2hvtXGx9XVPOHiSjIX5wUlfYK+Di+n2wX68sqhAP7PEOMR3/89SkN29
1QQbGDepcU613zT/RIENyheIhBrGOqeP+qaj5mNaxKVK+BU1MGSbyO+SN8m2fORR
cPTMhQRxRtKWDmxId+8IFAEvyeuxcWQ3/HooJllABX8MBilS0Jo/zbKYC/9ov+p+
WQmGd9eSUvpKIyvSMlYXzs8+1LWNG2ydQ91DxpoSsw1nhngw96xrmEexCiXGE/Wk
B9hk/ipDMJ8WDAnEWTeRiF0tli5tjLOTdN3bJV4lobGpO//f1QpowFQ0j7mK5PBb
LUy2sdwBfSseyHGENzj/I6Z1yX7LAD/siMACuolDX/DpXXc5YEA9wMSIBygLM57b
c/WulA2RgIaCzOCle7ZZCmiO98puwrebrYMmdj/PmSMnpfYR4v6Gww7hrmSBo2mo
CYBUX45C6wQJutIMcHOTog6UgGu2oB79iWbgDkupVuREx64XHhtgKVLs2w2qD+fF
hTaWFLzIiMQvkM5WZ7RftxobtUDkzup+pttrOs8+/3m13dqmLLG7XKk6e8UVqfoZ
5SwWTPQ6QS9xKC0a5pogdJfnzMemJkW4uWvzG+XTR7cOiIcXLwKYKfHxAdDhr8gS
O+YYW/ChEfdi3rEI7mWP2P+FyCECNKoN3PJ0wOgOTgSJ4cyjqAmx+vSnLfbUgqU0
SGIKCenlqRsdx4X4jKhx3k7zF+bEUBJ/JpqZsLQXS5owSv9JDXHGcftBLN+Smh73
1r+D1Sm8m+2Z0Zfm2o5fe2BCPBYf26CsnZJn7eu0nhF4WfI6vgxzsRUSk7Bz7+6k
17LxxtlzvqGjURyPW/BTbnLi9P571NxjQnCHL9ZW3thB1PE8XNAT2hciL5n6ewtJ
l9tLQOeqSXrAl6p+s8hXMHAXZWMgxFCrFb4lY4o4bF62IfN9OhgT4zWXtlbeCVEC
aV2u9yqRWRQPQLgxxTciPZcz1qllwKlBA9CsQ8ihVOFxqeX+cprk2vrptU2UEOGj
ljuNB8Bhm5U2he6UUNwkwtrViwXZtbR+/nDcpL/tPkXLkmd75z8SbaPQ1JuYFdAA
vdN6vdzlPVR4iHNK9TEZT+QOs03fTHg+H7YIuv1sfMs0YJtqNG56q2lvqkDkuzGd
XMsjXpzu73V4w6ntB6t2qtx5FLMmAX/DmvQDYDoBTGMxyiZu9XVsIsPOkhsbhrFD
SCLKMZN0zFzJQv2QRQKoqW3//gGuZ0tGtFoUMyjWTumnGCz7sZrGsNx4VJ25Buwz
pT/2m7NzAQX0uEH9yUT3P/2CgezmZ0ZGXeE879aKavbXNT3Jg0J0vVGrAZh6suvV
3CkM9to0OOMoef2bs/llroGWE41JLC5jhqpLyv0UC+tJcb/JllpP+GzqKCKG4Cdj
/v0DdvauvBTMiLYM/bgA4X9c0gY2KlPP6gTeDU2UVWLgQbo70XkCQd2dmi2baB0j
XCpFJUMDhRGEqZdJi016/GZs/VViWkCtcaFkAARbypqt/zFL4QgNigTq+gl8kj2R
z3dvb3C5sOKdGFyLLtfJ3IJ0ScmlOcOJaLAh3l80OYvIRQfPEfcrZfIwNNGkJPiy
rzBFuglbCPfHwfDoGJHMukSIYGSswoHb3Y0TvntDnFhSR0hL0o9LtzG3JEOm8RT2
Zj8OYD6k8MIJSZHBaS39Xp1WP+cQnF4XCUxdLCcCUpT59UflzczJrxggoFTxWlBp
SOK+oIWeT7aslARlYjz1iCTXzhn+4g7Gzm+9uV6PyChzI5kwjX27U/uQJcY8Qkfr
gCrXCmfBg8QVwSPQfDidUYUX+izUOQsXGj4c3xeYY+prEp/nmLs1aoP4zgsMJC1R
2PANLaIDDlXt5ZjQp/jqhZwGrXH59MK1PJpxXhSkzB0oe9c7/gbsd10kZN/OEec8
Y4crRTSillXsQMulzcBQMk1pmUHNJywaje3n/0GqEi4dP2DHwSfIsdPzLC3NswxQ
oPiH+Yd72eleiJr81U165V9FqybBadIFqozkiwMzYJpJjQZ/ciJs3LCyFQ+8GYom
hh4U4Pn7WBvZLL/1RE/vv0/1i7gtKqkPgU4HjuWSJwySbXZG6lPT0PWM4IzbSnRn
G5YzrL0ojHOKSZuPFxxQqYr323HaYtmUXxMntGXjOzR7FdixFZYch0VEoKDICI8a
NqfhgPj9lV4A2VgOmiSOW3A/skAm81KqHFCYP2dovosEi/MlzXv8uKUid+Bb1VLk
ziO1IowgHWppTC27Vbec/+pj/xxTWajAtiOZRmzXxM5UgjV/apPq6gkVcE8zAN28
cPPSEpS6JCcGIVEBeijdgOluvjSIefiK8ddz/f1oqyfDh5HLfhpZCkuUWdzjT8XI
TAQAblpTtfEQ0F7QOUxwmR+Qk09q6eCl3V+i8azPEP/vNHjaWsJkcL0EXJm1ArMI
+rtRLPF6iKcdf21Vx5FkQEKd/QM8N3JBsIhYJhiQDdAaSooo7schv0UlZ2xdiC3P
Ppue52Uda02gtk/C5ixLehwKtWkCG0FWOBehxpbyh6DIcyxU5xKibTctHL0xB/CO
3dj0B67bB68CzKP7JkbiiQnMC4KwrIAP/uUqnBRDIhKyTH+++eoKnEpNc/vFsuYA
bjH+VxWFiZNn3ptwqyamInSg8FMjP5isXjvsGc00xtQf7k43sgbZn1vnahkpFS4P
fuDhMJgd5yxyuRAMT7WkK/2EnXQG9Qvz2yTgjg3E6NdqHrVzgvJ5XH7I5Q5Los0A
XduPz5CaYl0EmzbCArud/R1WGHno9j7JsHpePMfIK7ZxbuuyyQL66Mw7XdhKccB+
SBrxB9Hdu432Z/hKavXPC67BORP19RT14JcrHZ6ShZaVE45rBnOLKAc1ci/BVJRF
dnDv/JgkfWHr/mcGdFlEcnGbrm4uwX7Poa3c2qGyye80M0jehuKkVhraQUTVjIQy
jwPx0MrTXB0cJu4v7oob6cstHIjWkTSqfHnPKHwjT/nHAlVN/xDG79+ZNLed43zl
MDczLHSz+3UVWehMbMlSgUdqMT3y83NWDzGnhKA1BkOvYumXVF1aTL/LdvDYr8hl
0m2A+fftBrEMQTfM/73IOmAsq4qRWPZ2fEw2tjWYg0oFQ0I1F3XPe4t9Yd3zvdWa
Ps18VxlgrhL2mwuLFc+HQYrm6YFYnY3ekC6wyUSxVloEHylvg+drlfiKisYhuhth
MI0EEbnggFtq/dB19faDAZvXbsyXxq6EMMOTc7gT7Avh39750vDYzrrT5YiLLQIX
Z9ga5CtZWU6HQtl+u/dsvf87mEMUTA5kStn/vFwrmQLIE6mlRMs2kzXSfV3JZ0/w
ODIYrq1mmblVC1s6DZ/OMnOnA73xnhAQKDwZdvUfGGi2r3XcpN/KH2fBidiT85ch
wdGksezNrsRrCtBbK6krI5KH6sUDYevJ+MnBfAUjMXcCzlnHLRZUwToVTf4eMJHY
RlWmgIZKafSFY3u+oSCxFOlr9jE3DyDxL3sLx7ijLsr8+onBihkGA938csw/AQd/
n5zFQUc1sScAlf2BOvD1C5i0p+Cn4W0kzFC9j7qjPPSNe+1t+xaN5gMH9ZjFHtyt
iAv+8jVdwC8UqjL3AIHmdtqDmLXYXEPV++8TijSFgLQOpthpWnGp+GjWcKpRx/OF
bl7LpYqujP+YM+HAJCjAX0szaecf8dbJymoWOf4MbxnxSYKqA0OR0XQOBt4Ttxry
R6SzYuZ/r6tRhMFzMEWmPF7WIaFiYLoGVthDACHAK8Y0etkqVMD6aItwzkdXudam
JaPt+Ekl6mrwNX7KLOox995LkQbTnTzJPdziXS8LN/EP7tZAmO+oiXr+3uGI1P4H
xvp0cZt5YCf5oJb4gXI3gYniRmuyuGNgVe0n6GTd5+XkRkbKi1X3HwV/VacVStrZ
YxlHk6LZHfN2axs5gVBRFjuhivQ84Kzhh3aMbcOOEpcRAGN5bcD05Kv+CPPtQnqI
Lazp9gsScm5LVTdtGSxaZqaRhZMrsiATkaHWXL1mJlJChRtbzv9xZsS+UpU+TaTO
jNU9c904XRO5pEuYwH7JFmQvUILCnBdMrmRaHdFMV1ATcS+P8dzG1Y1Qw64NJm1l
jC4yrs52sM52QgxIYoLX4PwBzoLtvEZXWsw7jf8JJEO2zpVJczJnBUclI+GUIBuJ
M/AGJT0EontJ/eZWQlaz4w6DUqi4qZ1t57rSJFskia5VwrO3/8AoYdcMPbX9KH+7
qDn2obhMlYRcV5/sswBBzn1wd5h45BjppgxF9lGy61XFq3tPktaEKnAzBx0TbEF5
+58ZFq/Ged16jjAD5UUvz0aGZvE6X+p6A2toqU5qjaXKIZhL7wQyZ0lWnGE3bzqp
XmWT17Egg9yWSn9vL60IW7WTlvnpj7nDjmwhVfxz6f0ha6jRMw8Qw8IXE5wtiEPW
lMHmYfB1hN4k0QzYg7USTGEmUMktNTPw2aptX/2QKLon49L8gauLDteJm3tRkIKe
1naksEHMQptELQrxk+gR8zsOggxGGTEUW+cB3MCabQ0hKsPjskBaeAKMfOKGzrPz
9xBZaElluzK5kC0kefPtgZU3C/5cpZASFniabK1UAmryZpqMSLAU9SYDqIdFdPcv
LtHjsJgWb2vzUx0jyKBTq5MGqv+SJEEI7Fbbo81ibHPlHyaso2zzZZReurLz42lI
1aCP7m74sSJ1N2INsJc/ygNp6qc4Bz/m8SPmhhDcj9nSv03WIGfPhcxArgDL84i9
tzgPkHPn1dRygvwmGstatlBno8TxfTHlKPYFHBGlF3lazF6Ugcw66CHgntV3Q9s2
Atkt1IugARkLys6eKT3bSZjfYR6pRcVunYinvKveikft7mpjoEERkUtWeztiibHc
1eRWomn85msNIfIGfvYmNC3MrWsgGbK1Fjrg0t8BvoyVoVV80hqdSZsCs9tHNbkt
ybH4X6720edNcYDRc78sjPGxF2IF+YJzY5Xcjjv/XzgaEP0U+StPgi7D4o8EALSw
TSy/YBa/k08/q4t0QU07LoDUVCxnBIpnW6mNWgtefLdZc3TYkprjQ+gEnPJgVN7f
lpAMEdSyUrn2sid3ZSysO3b69cjdFTv9f2HsjftsGh4LTT+l5vQyq7moSBXhutkh
dsWNv5RIpkYCxiy3MzsVOCyKk1L2tNZpV2crL5Ps45ZKTAvahbGTg803fmZIiQ12
0Gy/NGIDZsQiqAWeYc+gUXGSYq2KyvfoERzKe9cice/y4M+JAqDLQB3Pvbq0If3v
wRsjJuNv6vYB1tX/gIg27RjBoQT01MTyPtDaDccwKEOZqH+Uwy+oQxVgwO3SGSyg
EwzH2fJKNfP65wVUN3p3vXRGCAsQa+JUBnarkJEQRVb08rT5uzTm+Wgh82hsV8BR
h9qqZloqXNo0lFO7hyRlZks6Nh+IVBHEahLpFUy0aaT+8r8aanFIluBFClGaxI5u
x/d0O14/UcDAZI35GQWxV6MaQ9Kc/ma/DJofZ/RpGtznBbk8LVG4A7zLhpWy4teE
ftrnuRc8GeTK71KPwHrrkNY09vsXR+15QE2u/a9dl1PDlrNQvGgKoQg+zfLaB9xg
uzxXR60IgxRNH+UT2yOB+PO6szpHacP728GzsuZyg+8USVaKyXJ+dlxcKcicOZVc
rWgMsJ4868lvNjQ7UD5i2EZz/Z5M5iPTy8Iw97THrrUvAAjGfAfihJEXpLLwApo4
y8gg23w3xXYZaarJnNHe9zdCVRlxQlMTYgp001RXl6vvtgNSgBS8aaTnjQBfFw1C
2qMWBofKKGQ8KiNzoUO2zd3xTczR81WXrRuHd2SBxUkL9PdYmYWrcjJwtco+S+Ef
PGtQfYj3wuatIRgYkEhC9YkmmlmArykb4OWSlMb7MTvg8o2FNcjlZUficiQap36l
ah/dDmP31EW1z1Ms6CsOXMDD3/LNjORZdbw359onQmw8/Gjhu/M6lW7BMAeNjgal
NuMZw/LvuaNxNCBkKmG5F4bsiCDR3RKVWGCFT+cNVFp0JUklWwGmWF512MBWHgR2
DS4JzsC8sRZ8Tn/C6Luk6ms3hzmGnv9R1ytPygAcrwsnWB3DQVr9ezMEJpx0rCit
mle7PwKaiV0EJKhNYeEFgHwQyj5wZCW/yKL+5RRAk9XwiMd5qe5Gn+gIjI4z9e9A
/3ptlyDRLc+8EFpX47FdcTaPbyKKf5ruzumqoc79jgniHtGiWOvOV3irMYqiJMv7
ltE72qx//1O3FnOdSTbK47JqZLA0aT4g6PdumhraA0Bp+0dSB54BYO7z88EUILu7
YY/Jy9m5ZmbAN+ZfWKw3lDTyNHtPIfIeLj7dg+UQYhR/5CN+dNc5E5J1CkOmrCln
mfKbWR5IDCNNCDZJe1GH+lG3sVwtAJoOeyqOFxxcZ0ji19dHypMwQhJ/qbVZo55O
fghwdprQ0KwUvda97jBTASXLhTmRoyPrPoF4t1N2xcrX5KPktTpeSkATl1fBGsMM
K9uAZO1AztW4IpBxXqgpX26ISPX9/XIYzCNixgxeVh5ybFqVQsLnRRwfW+wgwE9p
7S68FHe573PE+wYTQPx+4zkzUWjxHvjax4aJOIKw1ZPQQOm/7qWeB438d145bTRs
P5nEdb1zI2CmQWjqqcJTWc5elaQ+1m/kK4yGpYqCKIn9t4eOysIf64xFQaDqwrKg
6euKn1xPlnTgfa5UxKR+eoBf8i8nszVQzFvJdAEmBAlQ5/iN35YwOS44gM+M1qJz
C96OANx22oJPaICQ93sPC3HMVwtqbpk4LBpFjYF2eDJpFS0sCfPlxGpd93vtwJOd
c0AFPge0jpK5GfKRWsovbWsyPDBaaRFd4kk1kAMWPRoy843++dgdmbv2xC5UEnuz
Tm6lPfOqHWYoK4ERJGySxrmwC+PtHISlPpT2puRdp2L3n6YflYbEo8I90QX0pt9I
+ef+S/Y96T2dDyjf2EmNr7QY27yfIxOlJLNCBeUqXfoW6KGsctV4D21HJV3fZ5hJ
qTahRKI9nOv12ni1R5agCQs5gghpeFTB8UxRxiVBq4xGzVTcsse65D4eYpzqEXtm
DwjkdFboWOpr4oZvT3N7DeQBFyGRL0gjmjNQjpIxUyj3+8nf7YYXlXlwiQmQYIkh
x7Tg1qcRcjghDFj777MVpcllNvQtk0La7bfKv9iTyE11OdbbI+w3XidUw9ni0dTZ
0RSkDpi9f2Wo4HDV0SMgEfzsT8zV24JzVG/KiLKfr19QjBLwDbK00K1HouCRgg9J
53SJJ97qzlmZCMOedH0iHfNayWTb4zpgcl4t5ph3I2m4lxNa6T9/0L1N3WNUsGwm
pKtYSKtwW+PooDA1VQQ0BHjzU7kGgR23Vo/mvLKHZ4RysCPWM66eptHeUZTxEWEl
o/SeniN8sPo1BL4/XYG6HnUw11Y0PQnzsAfq61X7kFL0hL3XVWel/PBs0p5jKMzL
0r10WKpQfvOqRKw766H4jYkTtoEx/nfaaxwwIwu56sguPPDQiMCvl4AH5FCsZ4o4
gYzhUUMNU7ECJ3T/wQSU0/QQzGX6Y+cquXZTfwR3o5EZhd4a8atz4G6jbZKFcU+D
C7rQw4u5ME6nTIuD21z2fWPWCau7hIAYF/grPvycc2XvKCEwNM1v3h5VAjfx2MW6
rYm4E/9Ge/CY0l+od7TaDLWBjyj/wKNpyqHF5YM0rlk6fIKrhZXkfOAJUCfGmBtO
7I91SnHcLxe1nyGYssHShrbBforXgeMepfTg6/PtMtVXrLVOYsZEPEgehwEBxkuZ
x/34c4Dzfq5rxiE37+M/MsM1XdARusmpruk7baYZkfVf8z5Aq4XhWuKL6wcvrNuq
HUDXZ45Q8KWBsHjw0wKc6iDMcAbDWcUPKxdMD5ZZGMgWXabP2gNmM0BVqizv/zpQ
VZcrNzkTAQajzPYW3GbRV8eFOKs7rv+9KQnWd3cdfdCHC5kjK+BXTyYV6NcNlxTX
4yl/WYkCZUCFtHPh5ZGDIdooZ524LVLcWi8JxKzbq4WLpCZn5Y4lwL5Qg9K3tR94
8kyT3fxJnctwq6OCn+Hrt6BuqLaK2q+eBBGEmlF7dhTLsrCVJM8SRpgqci7iZ/ni
5S7d+korRGjjEojGyDHF8vJSAL8zt1PD7rXU7a4vq6lhuereRxghfv+Bd2U0xhEA
eXvNaD0ZtDGJbpQbaSVdscT5tvSXgI+ejmIeVYNlPbr1z67dgswEtL/+48p3TRN8
w3KmDPzWJ2ZS0mZL1I9fPk/+eK+ta+HLiFa0aMv3hl9SVT1gUSECk0+/HzxRhNzw
/ZwG6BzDyOZZ3yAARkASRDNgH8Kxmu+ktXfBX7DfRcztmZa1sBhT7UUd5U1rxqQG
GtTF5b0jBSH2L/NvPtSvuIl2VKe926a+2uFPvSM6etvjp52eS8pizrHGt3kdau/8
Vb6OM5XP9vh2m0tMZ0ghS9A+0mmxI/DXum7T28oD1ho4dbdHfD/i7BCx4dhqziJ8
Nf33ONsZnwACWwgZMEolMFG/VixqxPotaVWpg4zjCm0DNWsa2eSZZSvmtFKWAr57
/o8lI7PRH0IaEOCi6a/X93haaHsjbY991xThwnKubAnm4PBdrpL1adb0BsBYC66Q
J2yodVWCQvV7MOyjZJ1mBiLPwccMZOLKAL1u7k2fptGKjmQm4XxRnejnrMXhfPeL
zfxjSUqAqUknjhjJCKEu3auQyeUMuHeG8pL30pdpDozleTiep66YmEusCV25lY3K
COfrjaDMnflMU+IXVycxV0zzECPSbg5EabwwtnMIBUE883mkICmSvUkpcvCDWOtS
PhTk4MwS/eQl64xEniLzYhYbSJybNJzLmY1tR3SxAhRb/Tx7jDFcbhtUiu1zeABR
bTYjszro+qlNoUoN7woahnvoFyKPHX7o1Zo/RLZHETn/gFswUkIHIG8bz8ieNmNc
Ys2oQ3q9jTDvcKqQRpAsoCtEHxbUO4UTW1LrRk4xHQve6PoTSga+vwMty+Q8nDrw
2l7KKjfi4a8kjmGxozriNEuNlNyMIMWi3jEhq4if0Ky3LjbrqtcwglLKuo3eyrR9
esVIv4bYrM5kut4A42cielcVyQt4/bdjRjPN4RWwI3m8vbnWG6H3w/TY/0WUrX3q
JBUl7tgbJGoo23SSWA4GOgjHCu+diNocHljI0pzE59/uH8E7PsmOACJAkLam3PWe
EjIQ6RgRQjLNSUmkGviySb5cJzd1Gj6w+jwqQjsuE0WbFxDHzlDcolImJTQJcNZu
8GO27nAuCOJU+A1cZDO0VnkszlLVSn+yGm53bYmA27lV5WjENEF7E01vRrkr2Xn/
jg80U3s/y2yjnFd6wA7q6Dzp9GJkKv0L6LVE1VMqNo0k0p6Ed88R++13eiSxqxbC
xtMQW6mFwVjBTCAJM38Va3zE9o3Jaxa3Xainv1GJSnrdufHuJgUip50y3gk5G2pP
vuk/t8gQhokEkjbVH7cW94Yf6mmXBaWWJ/yLAW8yBiGnIAmjkdQ+2TDSRBaMUtOk
lw/5o0B51nJ2Li52kMZJYjbKHfe0i79vipLMtxeDGhbH2ubQXu+gYsgxWsKAcjt/
/o2dTO2zq+IINPCfbepNhKfRvy5sMlgK1uM9s9KkFQ6fQ5mu9tcpHz4BM1rItwtF
UvH8Tak5Amsn0U3yGMCjITCN66O9NJk/N3PxKsj/LSzrj06ccP/6AYJvgtEtgmEx
0T6FhKGeUUh76tfKo2y73hMMqpIchFmsYrfbP4exMjbpyNvWq+diBdUX917uyI4l
IUZn4P18cJtERP7VRR+KUa27N+j+mCayiThY4euPazI98uDjf9PDWmE87er3pjKO
41yRel+ol0GLYUpQSDzm41CytUcyMmrQa9YcFG0o6icakpMLjs05dOpO50xuQbdw
Kl+TJ7OHnPPwJi5eGC9CkpUsKmdbk9zhXhRHIGVPesg/UXnBJBM7t4/vuKNEQAEl
pRQb1i4De3LTPfYjDLOPprNItWOmV6fMTw5PrPjZS+AkU1o4obj9rUdcGK4v6R8R
8o0/bCkGLWMXFeZ5kiM5uTsw36Z4uiHhap6sTv3TOPkWCL3sCBvQgaAYRIpGoV1q
cnb6cT+/I7AWmZbAwvF6vRAH266BBCc+YCTGfD0TVK8BnBSw2yc3OFNeklD5E7t+
UJdhd0rkrmL/qRqhdXvE2l03/yMHCUyA+9K11GqFOxrt3k3G/oNZ3/e/ZjFQfit0
E0BZ12VH4MyeMjxxsLOunUhAVymyaaLb+Hlt867nQVgtliPLQ+WKDkn6vaUc1kMs
9LCII3Du6hrPmVBZaqrR0uN22aoMcsi36YH1FceY0ZvEHxylfsoA8MdOgkYPm8/J
D0HBqw6f7Snsz2MGRebgD1t/H1FgTX6Un7QGV1x2LjD2OD7+EVuG3jOKivsq0nay
5EK5Q17s9xuR2VPiQq51QeeyaSaObtzaxt5ZTvebfBII09tOLhOIQxIa8jBv0UzJ
fH8LddsWoSVXzw4XFI3HOUxbX65czai6KeqHybj5pIO5EBpMkjYQcBjgRSs7NKP8
NuIb8ImwD+efsHoWqvmQQ6O25SE9+7LXY4VY30GuDW3aX2BlGHSfoDtQc+q3onA1
b1tGye/LuCAZgNXAP+ixYWQ+8Hf42nvTKe8i3oVr1nr/WslkIljnri4faQ1pGrIB
jGWpBzcjek8o0XSDZwZeSYyQFluREdgl2aPacNfoW2+nwYZN/iZ+bnIM9PuxNn2H
hwpEktgcfLI2eXCVdGHLYBU2rN2ADdeRkYIPftAkI5WUzQpPw9HJAq5JfiUphsC5
PPJsNPGtRIsaEbyEjMr/SrzGZCHwwV8QAZU6Ps9IaL4yDTsKyP3IjN6SHpkv1zwY
0xUs0hjT4xY5rl7B+1bXbzMaGW3+FuxUlvKXDs0FnItIDFGKyeUHRwe7M8rBNXVQ
H7WslYy8AVn63b23ALz62h8ZD1GsZR4/8Iw4pnbfStjPOxS+rt7/V+E8r8mUo6zf
OHKzKEdEg5Ifns7pyAK6tvw75macxWwdeLKUqzOm32DsrHmE2ZWLiWR7Jm/VT4u0
m7aSVGaG0hyTbD2iNEZF4Zbe5U0McHxrZL+b9WMmoDBLO0JrZ5mmOrjTMBfEm+d4
mFsODw9EfcblcL/WBjJIRueXv236RBRJDB8Ti8IHQw2DqDhL00o2DyCeBFCZcWxq
WLF2GIPajqlQvHbrL8rPY5zOZKRFmL2p2DhaM55WelcRPHOTMiZrbdqdLRVKEf7d
/bSDUusRWDKTdkgiaCuj/ArLvLWw22TnuigT1/WlvP8UyWdwh6HlVJJ19q/ONSq6
Ixyp04APz/LKMaDIOGfHOow3Xwm4WgPuMCBzIF5HSacziMuMqp82Hm/3ri0AbTsE
z7/xbV2pFslXC39lNT9KYJONrigZPyvqpH2HYOrHP+ECKg88T4mpskxOLNXHbFEK
XvPGtSYQMIsWhDEZV/o59trSVchuHZ1EhQYp6NgJTaSrjpO3S6ze47w9vtcKhiJR
iq2T6F+rNrqAm3MSaAsmlzOM3eakfMnVBjScEAWGAPZuACZyZU3MYVWVyGJz7jPq
IJDehwzWdi0FSnN1fOpUy5HqdjOU9V6qpvW9/Ipk5g9uVSAkWY7IDulLMSVFZAlx
sID6+a7exRe5YBdf5HWD9N7+aZ4DmyC3llG1Mw6XbXPQ0CyJRWWQGR90ScTbzQTl
+g3r2VnKMSaC4vm0jSQX9ONCYwBAhHY27FvllhkE0sRSe4JzjLcWTMiL2t9CYHC8
19IeRt7p42fOcas9PeuZkAZrfLHlmDWzJUleWeFOwnELMgSXuk82yLTDqBDnnCj1
V6/3R4sD4OIgWhoy1poKkSScICXJvzvN0xbB2Svv0CqBMNKLykERXrxbBCLtEV0S
+nlD6jh+OiGNKnIzILhSMCIwAZbM/NSUoWqtgoS+FchcLaexQ63p6nEul7XYHp5Q
FYrPKE0rXpDTXe59mLiMzVujVf2cH4gmLWO09F6V5BUif/nXSCxUi+CehXzZ97jG
t5mlbyN6nK6dPicS7Zqa9yQu/mXJ9Wm55DDVKDG5f+kS3fzymESw2vnVm/DqL5c9
NzNd73SHmpG+xLV2Few1DzL8E41dXPT62hnoiIHRToTFnoc3f4qMD+R6LLe3nhHD
HzrMSq/5Fkvx4iFQ741OY9IMjmmBaVfhaCzA2fjQw3KKZQfXSXgh1KtJXuVPnn7Y
K9LG1B/Jk5cIkVLmmUklEEs7W/UQIhLU2K9wWEHCSfrOEuZdqQqwLsEX+DXo04dQ
cbwpsEfLocxOyIJ4S2Zp4Lr884QQpQW5h9Ud5Ge4nY6lzxDOTEDTI1Knn08jIRLb
oWbx9wk6JxCMXZh0p345eHpUMeVHVnQ/Ujq2ty2qAG0A7S1iu97WDhUIXCLfz437
u2QjBWblaijkcnirlI8REJism6BOTJsTjfeGtMaE3FtcmDC4s5LwHGEbwNhAflks
o1o34yWbAqHS7kILVfRZbUcLwFHjhtHRdUqtzlMBkajG36SRPQhCIOttXIF0KJek
F/3TzvR35iCgkNh64NF1LQ9HZ+GM9llK0m9bjRguJlL1sjRHQB1N6PSvExIGByma
sa888zpOF10azvf0fyHXEL15j74ZiOVvQQhj7Ddmqlgel17B16hKFVzVx5plLspa
s7JxFHwhCfBUcoOTw6UMoNZ8uGAaqPwj+8Yn2R2KpfvabFo5j/eSrADWvIG+QubJ
Qf4VJzQ22hXqpTufFC6/AI6jHcEho2rEbJkXy5vnjG30ebNdIx9MqNVwNqRQUckq
MFytvWuu8D4rqqxCx5gxlAK8f0GX8JidsEDS66tw3zszOIYARS03D+RMJw7pW+V9
UVQrbRHPiVBXip7E5dJpxypfwCCi18xX56o1HUh8jeP0fWHIr4/bY8YVlvwjGN6R
oQwXdhdh0MHLC2651JcL2dS81xBFf4mK3kHuHmnInjSn/Khyxxt3ZeJlb/H+gOqL
gXxdw9pQbx16XYQF5JcbJ0kHHm2Ul3XMiMutERmW6EhrM73vbOP5Oyj9W5mc3lbF
UuN2OIcwzYyK49iNmZwJSAJvg0GX1tKBu8TIwWC1zqXs1Su0pWa9Ruc4qytvHGD2
UJC7e6k6w3LzkfLMty44Fp3QypmD9UW8vD30H/K5nu8EURPT+P7JFA9c/QFjclyo
BS+QdD7+BeEF0QAqezI+xFUgBKeVjI3VS21tQVueNGebd+RtENwNfHpPr7/MzTSL
dAtIKjeYeS/Le2ceFsWM39cG1iM+opRL+MQi9F5ZiV0361VqhDSDCgYy6xX3kH+N
DYTJ1opRg7pYCJjF9OUrMNVhu8dMFqTQmtA/5k3Wu63yExIjzVXVGFxmUciA4dHb
cKwKBDAtfVrzxz2u4kNP5ipvGvVvJmUg3+VEda2vbgQlUYfZk71sb74YBEFFPUTh
cWnQsScpBIAnR9hcdN7V6LJwCEx6+7Wp29iiT3eWdEB6LYJur1EyQiWBTtyMng07
XLL/OMmvyWhGQwKk3YDQ48tCj0hUHjX0UJtOrBB17RthVO2/jCDNz7EwK0BJeNpq
42zNhvVXt49p0ZUz1RLcbHxZ7vAvxAO7xQXycz+uZu1+a2DPgCRVCekIuMjav8xh
iglJ3FNxoYfj3rMJW//r13mAn95idJfAjXqROnX0s2YGFB+Rn2BaPChGsT1gxQtr
uxFvzcWtwLmVu0ICcsQ13MStnffW0oWKYMpTGb92Xoeiesxv2daeIZyTJLfsCc6E
hqM8JZgUBXXKk//I0dyYBZJ/xfZctO6AcO6QHZiEmV63PHqsOmTFA5G5V6UzNaI8
XnVBv+KWZApqeTq3qnEE8EDe9YFf/jvOoNKJm5PrWVAhC8NzR1TyZfGhUajJorUI
J5untovmWoZ1gk8FdhMuviah1g4bLr0gVVMVW+lW8AtrRLUAWmdTUwvY+Xy/VBHN
WqfHEvSk2pRguAVt/OpUE41gXwb7SSt/mn+UbQxvCx40MU5iyYfZKgenMYpjKhkR
BOWe26i1vAia+o2Njq+AVupOqQxZyox6kJMj4HAAt6BDqU/c22yDMGtbDSrkaVFo
diTpHhvqqqDKw2UybVCtTqzzwQtojjuiuSNFQoW2LRULA9yGT2ZWHmcAXKzmM561
AGne7n/F5EMwl3zO87rKfOCwTFKs7aVIwRyk7SDY4vZqT944Q2kM1GpMVKhbvfEP
NL38u75ms/3g60d8Ve+27o8Cn1poqEfMgcWMrijEQnNWSm+G9Mt3fi7qYAvFWmas
/zXj9BPOstE9N6gYITYFXC9QMEsu9shdoqiuQsTA9NBj/RSr17nhtva9oKUvvmFV
fvtFmmXZBlbhMaBmcuwe6Pebcth2VAQyL+tWvGo7Ee6o6aKLxZXLmVI+OX1xsLKb
Tgwrp5Ba1YiesojleQ6OBo4859xyfCtBXdSLSu+siB2flv4BelZY5aFSNYJm2KKD
4jQvQMMeByCkWH/+t2k70WGWKK5o9TsvmiE71Th7oT5UNVY83HxdKEY5P2zhCw2n
NizjMO+d8MWzif4YS7Ob2ut5OK2Uurpze6h7QH5jeAIeQlxZrWi6TM2qL6YiYoQW
3xtZi/IlX4wrhwuAlG8X6S9TvV5GNUTYSfroEXReETcUofzmlXLUl6Aus2b0W8Fy
Uux6zVsFVx9YlJbIdj+Ih70RUf8vJhXsZKD9Ka42PWAn/divbyNXXbukdqgxA+kk
6GT51cU38F5I+2ZYqlFxZ3Zr1ivtNqHEKprN5g2LGeHOe3ur7j3OMsJmebR+qRRK
MyRh5MneP0jhvM+c+RU/ywRU1tpXviWaaSQSN8iSh/xR3grWMH6nRXnmom5K6BLz
QXd31opCXVENvc1LOphpbR8QwZ4VxxrkAG7WrzdAFm5KGLlvV5s2lbRm2UZnUifZ
rJH/CLnw/HrgeSQw4JQCH+vCByGkzb+tjx/Q8J0uw+2I3SkoP/jITCWDzl7i/UMW
2XKUllywuA0EXESxe64e8wbi1vx1nyPGPI6dM3jGD1j1aChcaYZexITATyiA9+MI
MjTvK62IvZz5iPlkpLMp7NtygkVyMXce/9yQAANmrVTnCDqybh35yoygaOHXXadS
HWwdY2rqvB+yAosciGi+h1RiQqp+WNL9ywbb2a+O3uL37CTccuU5h5YS2lZoTU3K
rG97B60VNyKbu4iK/P7YUW2VgVfYKm+4kzd8vIz79anaa8tKaqY+4+EtvpM/hL4g
kRgILIqkvMWVGOuUPEDGCAtBFeRBrSRC/4FeoNZCYrvvB2l0vaKHxZdZcJDEC3vL
nTJphgqTYOhsgwbjKJKasF5GXYmnoL8MVv4jnCYqhUG/MTe8Oi8Z+iOPrXmd3tVN
X9t0ajRN1vR8ny0iARxzFVkcsVPuSvkWLcaIgL4ki24KZQarodxtfAhAW6x4Ys2H
X+r53mW33S7dX9cQ+9AnHSY9XL+pe2H5O0NeH4TKPVfJv4IA0AGK5POX5KbFjyG1
otLQrGvN7TrVWJfwR3M7cZneAY39SrxXkjHEGq9GtrLmTmjgsZtkJHZBgGagFoFD
7sZIGnQT9hOjA2QDlWqNyNOVBGbA5blksoNGk1dU60sYR6VI6SdOH6K7Haqx5R97
x5eO7oWZ/804+VFSV/M/+HQJrftjDrBt8fMxn2P+wbVdrQaADkGMHYrQ76WYX3x/
QkJby9HGgTlk6GfZ1bznlgIQq0jEYDzID25G56cj59HlktIkb1gb0GRW4GKp/Y8E
GBrQeabHc6FSc5VckyAT67wv/wOUqgkzXiG2loYiRcWRxM+m1e+dvEZQ/Llvp1O9
qXXsHO+h+QRwg6UwvcJwR/k7uQesrRqU4tlzpLUZ0rE/CMvLNGG3BHvTHxbHKN/v
F9T4PvlIszOnnyb7Q6zit+NeO2qxpuF+CXrySYwHDtEKMIurrDfNCU7NzrO0Uwir
JiDAHgo9ROndzASudhSZiRQ7Scq8QbhmlbOC6HHmCa08qmxNeCg8p+Fbb+MayUGg
hmYCTcBJfABxzp2TmlPtfchf5rul+5z0aT9B3+sku9vqGNlcQp4EKMK35mls+Utv
OpCdKC+kjyT1PieF7lktsZ1jsCCojscM+U5yFeNAq3GShNjgvB7/wgXBSPujaJbC
UnYBZe7RhyMBcLe/fMNKan/ZJvPl5DUxHdvq2nYa8bJxGrEl/FpO5DTU/kZiVaWs
FbzD7TJDmw8geLBqBJuD/ZUJAAzR6R88M7H9a2i0GV/iNmICUx3GCkDNE55wq1xV
XLItoTwjs/5oMd+bD9R6mDvjkIqoUuLNRMSGiiNfgoPCMFw2UyU67BK7M3RjVe4g
O17yvq8vlBaZWp5I7gfc4q2v6w2ThCALxUp3+Nw43cxGEfPBgtgyScj5ARXShwbf
ApvYAXgMi5FenS0ezpyGSCyS4rsoPA7MEteFHk2TpKIx318DVXktd6sr4JE9mYWF
EgXA5YLQgWTsXTEFH4UI6QH1YINiHX/e35KRV47VDNpmBgF4pDGkL+grEFqfPNtI
gSPk0MFhHT+P395ETbW5DlSp9tou18ukvkynrEJCPnxCD/Jjb9KeoPXgEcUOzKsr
nUiphk71itYVmFt9RDMTAFTFPxl3TXDZfgGoMKUio3cdCCgx0aaI1H5/VUpp0R21
0ID1qye03olv0VooVI7+oUHxI/cbSeJV8rXZ44USWH6bXl4Qa3k3y+CXhMcTlST6
68HFEU+dA4eEjh+hHY4R+Tb+m8WOcXJH6CmR/xYj3ZvMxYOhaJ3mBuc22x8kh81S
PzPkHVq+zRo8btSR3Okmj0AVabe9h4ffqqSs93b/tjSgHQ86Q8C1UBOeyAXZHN7q
SF8/tJvnTKVmSGy8F59PlwU3Hx3H8OAJvawQfJXB1OqLHzGnEO7F9sFw3l+lhfZF
kki0XuB5+F7DTFgOwh/HkbOLx30s5JipHYt8at0l2VjxoRbCp7RqXJ3AeJiNwPy/
UtoysNB6Guc/sJI2/q5ibKR7buSINQHgmZ87GKIDwheCT/0h840LTBglYI2RSRkA
6Ts27cLVYDqZTc6xgfqnjeFsyxkZ+tmdBRqLGV/mxlhBLMBo/EkcZNXWLhMHFeGF
MPYuBy8LYtuqdKRT8b8pHAYzTtgDpXO/5iD08r0hWfQwE5V5gO8ATjMQmHd1FdNi
xsM6MnuR2tlAVBeLQ4MGdfhrcGoccFLp+4FVFHbwuFWEivNd9P67Iqnj5NO1AGcY
zeqiXGur3FnlMiS39HQVGCEaylGUp4hkLqHYTxaQE9XfBKsV40l1SNdfjR7yi2zz
PDj657ZC0L9qAiNq8Cbtb+QfV+NTxa5R331kf/QpQkE+CHkZW/aXZS9w7VQWv2ow
Y7Wjfo/SmJ0JHXsEUCPPQtjialsaXffKA2qP6dJhmTThFAVE0GcKx8dobU4vBPtm
03B4/niPFVZAjWB5WvqPOEAVS1iDzR7RfjFMBxvq99N0UgO0tg8X2ltX2Kz/3LfV
SDi48TXREfbCij2rLhiD8RJK/3VdQq5NZJ1LFrpmxT3bmJNen/wxpdT08mURh9c0
DAk5wGp4SVeWi2AWexStqERhH4PwN+3E8X0pVwm8x0EUaXRd2yrKGdnYLISWk2oF
37WlfP7YIELaCkHQsLAifQKDSYlH2gvZf05K6iulgTgl2G7vYkWIRvBI3AIjo0cQ
uRU5BwDxbiKIC6RWbwzDaw0rFXkwQawHEOI+IKkVOVr3kBythhGU0/z27bIjRAXv
BIvAlbTelL6XTYP9IWtUJ/a4JQfnbD/tweJ4KBby0GLa6U0mgwtZ1Ghlt7SsR9u9
79QRUNBaeXqx3bY9B+MwoHQflEkGxYGOwNDC+N2Gh8GC3tmwT33WoXPuBiP3aLZp
iQqBrzD4oCrmdzJJ3rTTqOoeKkVAr134PU7fdSikvLXtcqTWDMiS6XltitqOdczo
mKcLqp97B+QXLlUY+c3cZukX5EaT4r+pKi3LY51BkSyl1FK2HjnLTe3MFVuMtGlc
Q1LsZMWz9qm6YCjs+k+WFyCzTbpksxtrmXkkwMgJZvXtY9otSO/dzdAlS4mjXV3s
Atzq1BrFB+wXxa/TtrPEPCxUfSyC4dWnLnLPUQw5fWaDeIqNYwClrBNtewifWKLe
pZLtdzBoFdh3YhN2svrKrEcj/6haZpeF6R7qQyTHMWaf/hq9rX0woLES0ys2+4+2
lFWc0BLDDUr61ftVDdzln7xhpJvgWWNAVfPnebppjLdKay64+YTud1yc1BF6RLhD
Vs/xBzoUZ83/OfwVBKX+kMBfeBKSJgN3BBsijoPxZ8eBk8506epyxayEjKviUdVw
lfmbASLkj1kBYvCaggkkM2ocJdc6WdklQuk6b7K/JezW+R5zccgHPsF7YNMLBhdc
/n0F2fNjSHSl0h+hI4dzyRAsjsRAuLccbhofJGc4J7bpIlv2C590+L5L/fL5hmlW
N0pzRuZfPbHAuLMzjaYo5sOqGg1OEuLvwL5/omCM4edPcgaBwXhXj3+9aA9Be7uX
AOGm/GqnY2y9Cyzc4fMA2WBciTqzjwwBRM64N1nGhmyapMr8we2UqtZRwFftojKQ
u6G7vqE4omyiGpNnAbxSfNYTNAUUUMW2YicllWYi6AcGWMCTian55iBYSXs1FKV5
hWamMc48zf/OP7NEpVcgOUlDYnCOde1B5KIUUIq2BbYg2JLI2pgBg/QjYr7Q+bYp
nI4VziUfa6u5NwrHwiBHIIOJs1fegpwtzmWiTaTe5F6unmOVkkPJtyUnUtDpym7B
HlPgRXEqKxsTni1Y4qCCOWLLKzwqMh/Yc/WIsqGYt3QOKPbD9ybx9nxLvIwjhv1a
IWzebsLtCVBZy2TvyOVtybuR/sS4dI6KgcpemaEqZsD/QR1ZweNpXM6kyRLW4n5u
FY/ou4cf8PnxVVeAzZ86oUca3rEaUh2dRmLHkRLbAhoHAEB3eumeIthbdvheeCnG
eWmvkOb+gvigM2EzH1u9W+yoTVEqNxv42qWDn2xwKs8KhvYmFsL1pPlBE1jmAcqo
JIwVxUZe09YewERPSNIgrroDmkOg9l6Uz8BDVZie5Q8X4PCbZqPIR+eakJ953Rnd
CfswdWrebCCo3SaH/G/ivKevXb4LQxjwjGOypQlMDH6+9SppOlemMTQj+90mj6mj
tmJpz7eI3IssyppX5JdD/jTSnscVjDSydHsN/EuAdOsZAfzew8ibG6BjqphzpvEH
QTbQeAJBHglvLYH5VuP1d4D8nk8OHpwzoEA1znMiFRaMzIcL6J8s6U6Tp9DY1ej0
fJbZpw3KW3Bzmbf3qkXwGSPajX6ymO4GL8ODKYlV/w6tpSNN7yL9m73SLIn+XvG1
ienjKc8kBdY08aaLVTEgust7nv7qKh8l9QENUWFEC4291fvpHuTLcEYlpD8GeuEE
D5eQqHY5v/Uiyi9fv3HitYZAymBXKzrr+1//am1daCqAJ3aiIm+o1tiSdkePUl+c
fFECjGifcl+pTODRnqDTH3h+wW4QS/tg5FqqI/k1GWRYKwImU3MO7IWeIl3ZtLO9
d7PaCIgRERl+PlyTjAGO+5IVa9niV6NaN4v0ud8gXHilIHYjNSNm4PBOjz5IZkJp
MHrQeg8GNda5u2e4PwqGED1A6jJNiIbpDeLVWBT+E9g8N4HFF6jxjIzb5Yz2/ySW
vPkm4xtvvtQEBSJBHwC4OlHMU1dShtvSTkvP/cN/UC7Se/D4cUu1+PFG9lkU0Qwr
g1uw/odSJabtA3JKDiTUU/r49UzFcsHWH13hTYocWTZ/VTC9x+Oy9vzMdS2qP4J1
BFUKvZ6hSebRH7baXaaJqgyqR/dwvXLBbY2LdG6EYywP1Dd1O/kjZnuUdygAzpcU
jsdQ8HeQjK4toakCiF4qtqAMGphmQZhRsDF9Mx24Nk/aeE6Q5aBvV0nEDPExq1Y9
T/k7awq6DjBE9C9G7px/ZzvJzIq9yNPH8wKq/A6N+5fffqfq1iePHjiWd+vesUm+
ec6UqQ5FstoaYKBFASVElfylxZ8tPUspa1zFN53maDagErEA4H61xhCZIZjPnaGU
EGhSu3qXkGDxV5dwl+l5gYCGPKDbATpBDXsuJcToYGeafxdHe+WV6rYwtpW42XVI
vfoBzXPKCQCe5dt2RTJakAGUl36DAm0QcrIV/UahNKbCmKnXbsy748qRpuETucBw
Qp+18upgurgPV0Ftm/xsUo5GbHfH88JsAAklZEjs5Vseoac427lPjCR/0GWrGqeb
9ZxIKYaipNnaPfuY+2urTs45keWgEKIrveQKsg1pTwISDmUQgiP2V14f7jcc5RbE
y5ZgMuMfwkpvRg06HQ19lWs+p0YIfPNS3hiYTfVw26Q2rQQhFON6DNz5fwfTWLvR
YXIS/Gs2sEaRQBERetihiSa+L+kYMeElPAMXV1JOiOyMNwJCOiXWyuZk4DmtATwr
0NB7CL6YiZbErPhvjkTlxccDXcb5W4h6eM5KN+/MfriO/B+95xJRMThMriW8nnyD
jRycln/sinnXwBC7UhFT7IPzQjLXgoUkzqUKgI0sx8dA8MRCBgVbH9Z/EIXevqFF
z4h9cs7/1eFyquX585jAXe/f+trz6rOSdA8cuyr3Much3T54R6ZAD3PWbb5yWifn
bD4ywy/KpA56wB4A1Gy/v09CH0aKi3jnemca/ZMkO6Fw+HyIgspVwc+NPJ8HpXSU
EiS8rZpn714wRgil1IRn2jyLCvVfd7bR2huWh+l1BTmw4HFM3HqvVvmtOXgL051X
gH7ZiEEtXet+rt7gbv8Z9LSIi1e4jG2WtL2OceN+MD/Cdz/QeBh9Blz9OHUlJCFN
VWicHa0SAVhgyg5gBFzgIv168IMqn5cXcMsHusYurGbdt4P61b+WvkcV/+2sANIH
WzePUAcEemqr24QqYeYjt35qNJof9SUkg9SGh+TajJUNpgQrGVWeSL7HYRwt8tim
fmqUE/pyd+1NnIwaCRgE+LyrRDL/XQO7fz/KaDllwpqtwzsIudZJRT3U+R+DeNg2
RmrtZIOmEMuEoN8btyzEsXz1lqlVG10xF/gbNrYHzwIggarssRfa8EN8nt7m4k6G
0OKXxHJFy6G69mf6Wf8qg5Mnle88eZEbRIGJixQ5MCGnRshGuRO482RR5O+TkMSs
iheU3JWginelxb8eJLtpB67sob33AHNkt/9F4Jy/606YT3Z1s+2sxQUyCRpsKMZV
EhOPuAjQXza7TvKl1JFrwaf6uf0qJGuv+6AbVTm4PwpoOks81W49NeBtDBK2ci+A
mupr5kbr+2o6qeXksw+aWyzbnoMyEc0916L8lYFvcBXWwke/MmPSUaBeXZQZhKY9
w70qwbPDJmK+pTG1+ADUS+Di/nQHAqCxLsbPxw4OGNgrUU8cfVQ6XBqKBUN8IOFk
Exr1zOiHWmezo5gs1VTGqh0fl6pFk1YedXO8kulm/QJWbiCMkHBW1D8RaYVXd9R+
9JcOza8C74HOikKUeeidg09afHugL1UeozLy6Zn2BeyDNp9LswkxgqSLRfyZShm+
2yc8E79Ouw+BaqdV8ViTX0u6wHfD1DGeBJwLeKUx7qsDBNVl15r3aHbrpF9rZiV7
Q79NS5CUlk+Ye+fHMBmjVgkqNXxGOToKAscU+52HTt9drzobAyZenK+ZhYLqRpfG
7XuD8NGoHFwyUttAuW4Ur+XRmcqdS3QJ442Lpx8MV6rJmtlLOkAom5mQHy1oRnmb
zINNERteC/dId0V2jSG2w44DjkT2PDPvu44F0oMbj6LQqZMNDYrEpDxdqIBG5jvx
XTTYnOHNXfBjZfkmtxyifW8fC0ZSBIVcghpFWZeIXo8dbz43dRXZNCWXrFsu4MMH
TiiXc1E37AD9iJB5Ac1H3u8lRRZ5CcDfcuGk817kS2M9pi9oIBwiuYDP6cd97KIi
PwNv1r5lfZoPcBgcmp5n3o0noJXulO0mhAH0M6kV1ORAh7ADe4liA7FRBqn0DZbq
QhQ9YiFIP9nMG2SXy5+0IN3nPDQ3uu67HUo4cWrgpFeEBD768si7XakUvo+X6Kct
vdWa7JdM9dx2XWJMiKzmzovi3V0nfO0tKfF17ye/ypFp/mvZ6/LGMraskXy41tgg
2b1pUdiQWSQpN9c8pjkXQtw2ONVvi+zf0hiWGbOaJmv/gTMsiQlhP6DLGlF7DihW
/hzCbe3jszLA6e8+U4nByC+d0cw1V2foqlwfCuEwlyqLF8xlk4i9a46qIvG1Qs+q
hposTg5ArSZRslWyxJwVbNEIeHi+aI3+Mo8rGqpFCRiWnMKfB9Lvi2lLg1nxbjgO
IOIJp33Os5CA7ksy7SYIY0m7Y1pCohS8QRu7+sqwP+ctUlNsvsDYPjQOUrt9F0X+
kdsZLdeHzqcI/N+44Su6h/VpbUY+V5lEs2aDiPJdm1ePTjznu0OyG0vbGKcF4ddk
7aC9QVdFlU5cdcK7kHQuu7S3IeYmZscBDeLQKmLx8iXyPwSSVytiPyrellh2xxHW
ynSx4+Hu5F3EERfdN4aTzM5gXFVB/PnhfBHXXgXHk6E/OKZMDMN/M+1N54PKOQkw
V3D7IkqXWLX3/rZqlq+zWZi5LQ+JdcnbbGUug2cKCHQ4UEVXbA0E4xp8EH91E9fs
dWV5WAnVnZCfEL3alocB4AvPxLwr/M1IK05OgTIZUoIfbw5rBFbC8UN6VEktAtq5
89Jbj1RSKpEQuKuaoenTblZk2zlSZuBpinOWK+LGVxf94t4J/L9rubkEG3G5DemV
FCe8XWwA03SrUluyk56yGXAUGfwjMBcwfsSF1DhgP7oq/bcUJhBe3Ggtif3DniMt
DvKFFddcF66FpJ1/mLQ5yGgX1ZmQPypgtbjirtKdaN6B+ALwnK4kdJdZWE3O7exs
QDaTNZcZhivxtUKMnMSGuqC92z+phh1oQqxZgeZG4F1ptLa+nk/agE/czWF/pNA2
mU3STIFnBg3c0UPNkwNSYNiG9vFf0rR2qvs4aHRA8n7INKMEUCz1nJSDXzkmVY0g
JUnbmocpPT0aGxI2hZuGCptlx7Ix4oapzpr+KPwWDAHP8rT2W4Vu4PfLWdILYQNW
eRmqr9VqGrH5IXk0SjEzBAUi56pfbCX+wRsgPpO5dArwuFRYvjk+SR9l1QAyy4QV
HrT0AYen27GfIXC5z54Nx+PqnasHQtXowdayp4sX3YGM/6p/x9Zgg6BPAjuCyies
PzH9f0cA59hyNJtDS8v4rPwKIE/QjgYMghKAmvPY5UhEWgtaarqT5O0Vn7GknWIu
UIuKLk8KdihktnM7Zi4tnTwUIYpTKGhnR5oqDR6Ija8SWRn2iTUbSJETOtBa8W9x
hDMHbRX/mIA/ZRXKAnE/fvHF2wI60o868roOYdq67ahEmveBqTbNI+xeuiPE/LHS
fq8chqJrC5cbaX0S2hlbgD6MQG8YTB0a1axWeYG4ONepy2x9aTs2EaWx9fjpyePt
3ekawKfL/JZtfoN/aFtVMNpPucYTtkI8qlj9njFuGnYhEtVGxkuw/P5MbsITXT3R
uzexxbkBMzQK/+MXHZx4WByR873sKhDjkAzDIavrf/igrf5AsZyMqqx0p8AfR8cp
kJHme9Wuwg9L9Rfzjr3xBVcVQopm+izkcs6B1sw4HpjrvQmHay7WdC/5H9S0sLSd
KCebmJZn1lsiqoFVCZIe6axvBXAYW3bHrqbuJzpOoFTOCtFsmLwAfZC30TgdGkq3
ZBPD8hSIbPoREu2Md0jo6j7SumEzSOWdw1r1LjwFgigkFGZl02dAYwhPG7Em+HyJ
OTtMh65LjGSawNu/022gwTTIPFFFgrMzyyLBMF57qKf7C7wZkdojLz7Hyw1OrAVH
FROdrgtynhxOhj/JmrfIJXpgPDIYeqlsnhFKwgjqFt2tILUUgG6lcx6+9pT3gFha
oH29+gDS0l+E12krHSkFHfYhdJSdTg+zqXzSbXzCsyKw/4NHpqnQgtLmUM/13d3d
/2wvPQWmMLwDzhRHRUgr/yb16O8zaF9IyjzRR1JNx4YvvRIDvvuZe0zl6jdg+eDW
oRNGpwKT3CHxEi85J1tUjaUSXt14DRXP2P91595/jVpkJ6+bequrGJip9eLJiL3p
jU6WvX0hhYPRCE40pT1zP7/935HRonwR4UGCqwD1gxU4vAU/I9tu7f8qEmNvyUxW
44OI9/e9AezZVwcvCA9KxPC+XhZLvo7suh5z1FjaAWbQdT3FuRdBgq5gi1th5C1h
X/5Cux0hanSido2Peu8u5tAD6sXLzudJtR9YnkS0QdASB7HzjZnN8zLllHziX4b3
D+nv94EYhe1yUMCnyAw98fWTnHae56H4DyzCedEMla75sJx01cytJmYp+1Z/inzK
qsAkEJp2tVcVFRkujlqIowiFwR29/+LbpluLHYUnAxZZH06pyeprC/19VSErkg/t
bUxoHnEVpsntQtKvTjvxh5jKNNhlg7SZjMx0Kfpr7m2ErUVYT+IUacpYmMrlDvvh
rvOTrzt6UdvV2wNpocWknm+H99+X0jmBaREJgpe1dqqtGTw1YLSrFatVaD8pbYUx
Kbx7I+z5WCnCvuRv6Y/of027h6RiLVDgoQN0hUdN5F/T4wJxbCEIJFlU79kGyxVU
vHsDClDpuLno2y4U0hsKkgI8Qp3rKp1Mv6JPdUh/gO0abaZhPf6cqU+II5n5Iv+5
WgsgvGD+FhrjdVv57LMVHvAndXUidR6f+qyhEafVCxqjjKuTB0OW5nhrQ22w0tzy
qAysoM8J1By9IYjRUz+lI5rLzIIrKf1qagwC7Uu1WiP0Vd3AYs18oeyz+9UBhUFF
8VbHNn9Ag+0dr9bFrWMTCAqgxtkbGhcVE8J2uDh4DrXmVowbOitHj3KzOlFqD5d2
34zbI2U//WK6iGm3QXMlC8B6GAaqqlz5YYHXO0tH5b4WbcU8bBoFRdDF9tb/cs2B
U5CKiYK6UXL9o0piWHEikdhmhyhLhow0fL6tXET9TaV8t/1Z8DqIOPYFMXTfWO10
eB+E4CD9zlW8I2mSovEvEq8dueJmVw6Y6euzjeePmHGnOBq+tfkIV42rNVc9YLGj
qgFbZKeLkV92pXYiYoBfiIldglASLv8p5dnI0iz7GhaeBjReqCAZqeUWQl6nJYWk
hrgU1pcl1XuhM7k0jXFNzly7Rf9Er7bTvisFd7OnRIa3z3DjK/Fjo3nb7N3BE/4B
tu5udJaGmvce0JLsV3EcDwYHo7ElDXLNF5xmeqCzAdVkEF+3ybArbUYudIyQ3Hal
1LoZeMLwKWNTAYxm+5RIyH/eTekKXlulFnZR7Cg1Bbsh8P/dzGTiGTtYy36/tvPF
WgPdz/cAPiAU+6K59i6qyc2xWOImtXd6nmOLmwsgf9KbM0+Qla1U1VVmICp/ExOk
hkgSKsF1ywZV/yRfQPtYqaVpEhJdR/reOIYKYTrDAdX769HP8orOcfSdo1UXrtXS
lqpw8guEhokFnTl2q2VN7owqw2kM6rmXkv/kKpGt9V7ynsR2VP8NRNxuvuDUTSJa
J9DYR7qX6nn6gOKFM/ptsglVpESu0ITGDJYeoAViRfFayIO1up3t+Yk42c4WYEhe
CBpmiFraYMZ+o6AUH5Q98M+1nNTwhbiE62F5La0gSobA9rigLWZiIJP9dSoYdmmY
fFG4S3Kka4UDkTLF+byV2c1fa8Mx116bQhqupeI/ZD5MHOZQFWRRu+jH2yOqN8MC
OmAc70T5EFUzB3GVKoZDIGsc6sBbGXFtpFbiHdo7+9kCo9EIQ+3/ZJoV8mNwhGd7
u7AfaHl+pbYQPZaiUnXQZmxFgjyGH4AU7AiwOS2CaMV0DJ/TOZIYm3mP3qqBBj2i
6ITPf/T/rv9eCs7C1KTK+lhLH95ScEW8PpgIyoeRAjk/TbtfA/376F6BiTv4NJpv
+Jb3+92zT8PsnW2kFweHWqz2AkY5BIX0BQj8cHopH+1ktXuniL9KaKTTUCCI6n8A
MmHRvSbqwGQR7jjHn0x4rfVGaBtg8m44K9txqE9/qBFwABhKOzvOZuzgVnCegWYY
zqudZpoWmSwpP36EZf8a1ado6IR7AXMByEiU3WX42tFLfEwglPhozcEe0KFCwQn+
xq3wXdWw/wNfLt6oK5ycHvI3m2b0qKQ0qyO5+VcPy+EYVcnGykyhwZvyp/DXFk/q
JMgqgfvc3uOdSekuh2PT5bIzTxPFKqC2Qw/zsh//nGvrKDHxNgmDDLa87bIrw6tp
fZUW0yxtwvDVeJQJ/zlTnmfS8iaTd0ntZz7UoIlTGedWRttsxPOGMBXg2HHxrkFO
WxkG7uusJLmaFnmB1OqF8yZsQMEAgTfAQpXjEdJhntzpqfJOI+vcbbGIaygjWDiM
JzCXpx7MDMP/BAt932P1k0WTP8Pc2QyAKWCSoms1zzhrXpV4cXgdpBd1FrT5SF7U
s5AxGSdphe14nxr7eg71TdQuQKaeKimXjjig6ekTLHTxkW5eoMED/mAx+SbM3np1
9hcIYMDGKl6XhqU4pWPmUdPBfx+owqF2dWJYtTh2JtqiJ7wv1tF+y395z/NjkpSR
/ckCeeYI19M1DRCl9VuvDR0vai+sUfS4kU2vhBOJr8CNowiXJ+Uq6Ighukij5tB0
jaTORFX0nZDLf1ongYaNdOkW9tacX+r1/RdLpcPhzk74iIYVKa3njvH65nHozaKW
NTdA6Tt1Y3b+9XWh+uK5afOnwBBjNALqccJNbJqS/YVOYmDidheye5h3dLbO4MEr
AFh/P9vmDXVTOlKmXWYKZA8/lFwOZRKVXdeJElKQ6MYM7VHYgEP+dfZHr9XXlQcf
H51jXLtuqTNfxPBJHphzfbtbYM7TRdUIz2nVHJ8h79FeTUZ9uqtCceVMcFT0uxES
LXiunRpN8BEcx7LaYiJF11wu3D/nwbeXWG0lPVYae3mP9aIhQGc8rAKaTOqB2/ll
p/9WYhvK0lJ9Kf7PVdOVyD4tu5RufrbW8GYtyIdL4tF4Bs2QKa+mBj9hVio9MWAv
p5BW4WxE55GV4EpXVvCRRSOixwtM6+Z1EfOwthrjPwEKKhorDSww6cZuQ1lhfOwF
u2/2XRqh0FmY3I54W7O5OdxSlUMic1/33uc6cBZ+X6FsZfqlq1+QhU9jxOJBQkPb
PKdCTBN63ymE4eKE7X1jLUEeqNohOFD6oloq58ACPXcHbvs+HPyaT7KIXGgyAGeI
od4HxpFKH3/y8IY7ACwg5n36s59JzwlUx02Wsk2efsjQ+9HExyj2D9ZAXAdWQXxN
j9LDbswstoLsLSO9ZRArRDTxdCL/ahwfGCX8rwNcfmq6Ui9cYjtaBFtg6FtbjGdF
1x0igmP6+iH5DHj0dwr4mPBxBBlPYDzkp2dlp+MANgKxidMra9bYreEkM95+1v2D
b73FoW50xuikOwmcK/qYFbPUIWbr4asrKMxHQo5BpoGKgfzowfjJxsTOUWY6vKc3
yBzysONxpioNPtDQjt5kCiTFwNLDWmUvjSm1zdDSse3l4z8AhitsDpxob5CRcxKk
0X8EgTMDo75zVti/9K36VTzfs32G5jljVo0b/C+f2M25KowqhfDZATA357fGlYCq
jHp/lvL76BKK4+sfGWZvudNRQ++0jocUFol1S0xVThZu18CHUjdoca1Kd4kKpP52
5MhmBwKodzl6yGEtZT8AHy2cseox0b85EIovueMADXKKe00jJ/yagrN3NsA0huvf
zIe9ebGLFl4fvsvFrzUOS+zbsEDPp8/woGgbf2ST07FXzQNRlzACx4gWPSu4tWI3
dLrhSMxatOYJXdpP2vPyPPyv8nKhn01y9HfjqjCBvqe206ZNkzUJcEdXG23ncDk6
6smkhXM2/WcX/dph9Emyxoq46xAXpVnPvIbNc6rNjyS8HGHo5Hfezr5S2rRwaHYi
AMWthRhrqCwbY6MNSxNOrBAopb0rAoC4lnAwh0JK/4UFnXASq+JmuUNWjH38Yegs
yF+/ArJf3QEZI6MYIB3WH/GPmGP3EICpQxqjS3y1HtkQdP4p50bBhasgiCsCJCBb
wLFHLbTgHN5p5e25fcOJKABN3+2EZnQVGtBah4z/ykl+3CPk4ZJwp9OHoT64i/of
HwzMQWq9Bi0pYl4+h9j8IsA+40966tC0N8k1nPJdfedUxwOpdInG4H6SxdpAiC+h
0NQAkkH8MibM/QkPRLUPONoLgQuhOe2+Yrclszd+xlQmlPgIpdKTLkeRpeperJgv
k/ALWLi8xwda0mp8bi2A8WVDMGBPQJdhTMQZ5tvIE64MuGBCbkFYCohNTN+O6LVe
UeGZLZkFUJJZ5oggi7Q/mAbvfMX2Pcfm4TeDv4dPM0mhaKN2xpScZlycJHbeP2bU
4vV5OzOYGZoAcQqBowLu6tyGrb1e75x+RsnsWlXhSu/kjgOCsyc+mKJBzeqRLBXQ
xe6GB8xPP6h3wrRtFc9B/JEg8CXXaVmK7TREzFkSG32zjSAiQcE+lBJj73w48OZU
oRH1XCckBr4y3FRAUqUQWllI319xJl/84rnbwgLNshNdUpUGgbF5vpaYpSGnXT6t
qApvZ302DOO8oaP1xR1xftHEJ4Pl9g33lFGBkQxnFgmQJVnkxCJdZ1I6PgEAwo95
sgvHKJvieAugXwEFqqJoh48lT72yb+pVaF1X6xNyVdup0layz77AqVnhLPCvYFD8
3AnOdxLF5y9RGYmQxG/gHr+S+3yNGzJAjSp2zidk+YodOWdatJ6CSCglpA/YPA8/
pm/8Ezw6GdfOKepguqgs03SKpeh71yhSeOVU3KfWjbXlYYUBqfEaWi+usVDs5WDK
J7OSMT13hkAB6Xg55rAaSVGj++RPZA66cACxQDXylvxo71GOVdmsHKYPnRWhaBoC
78bEi7vkmocN4uK2kIizgMqaDgLkw5430ElYLL37BzHKYZvWmMpNiFbPoM2shgdd
ZBNujoYd7G8+ToqThNTDLdjw4ziB1ljj3AO4irvoVNKFRCWD8dGq7XR6JHpu4AXM
B0Abk1SMBhkj/3UxYD+1X2UDKm0lsyw/BxdxoMMwo6bTJVMTGqx1dp8no5S0zMCm
vpgNBLVykqYUvu2xK3sUalKZgEbihtG4KWHnwGJqxBqKlcbE8xTTLpfnSj5U0vjg
DiBXktG4qK4hD8AZxc+yRGIUmsnkIjziYRcfiAeY6A/O3dw0S4GU6zTusA8w5M82
6U3yeJ7G2+fbOsvUjEiGseiq3JKK8dhOef+q5SopY7eNU5ku8uA1VS55Potzc/5b
D6PddgWA6DVGtMt3+/nqW6a5u98UIvp7enYaE8tmlFJT4lBF4hWKKAoCCtZXEZfF
91202ItRx6J4BDn0X+vxFUagx7TAL5ODXnDZ8yjehV8BIipkhDgP9v7X3Ewptrh9
pfygVE9LUBsjDGt3pAAZG/BNOWf8GX3Hi/PfotPbkS9Xt3/zVhI5MbuH7GHfcmHs
uT/veNmdKWzhrNFBIihla2S2L4p7U54Q50dmkRuJJZXb5EgzFyHqFi7Yy+oYo+GE
54xv2VdvSN5aPwzyGOzcrWnW3zYMIjaXR6Sd7QAK682lKQm9SrX80tNCQjuf+Ism
sBQZxAZiaNu132phJ8fvTEe6dYX8ksqUIILMpm5GIlAGLJkBjcnlF2vInxWPy6s/
L37o0EgOwYDVefLCCOeGTA17AB6pC3ZfZuxFW+X+qFYGdUEpgvs2LtDy6sGZkN/c
sG+hw5jcwk5lxskEEkbTQhahmba+u6lSneb9Eqraos+A0WNPfXrLPhZzixg3LukB
o9TemfWgS8mpDMc6HYnEJns0Qm9m+pzwRxUNWyAtq/jA7OpZ2yWk4P4s/JkExycJ
wunT+F7EKtFkgsL+mX7Jr8tYVn+DQczQ83R+jThHeqv/CfCIyDy2iQlyc734aRtz
H1dHdJFoJ9vuYLPFF4PLvSvIKL3fdtHdEQwezdchJrVZGdLH1JlHCp5U002cy4YT
NC4f3JaOs4nXW/0Zk3fHDW55dgNTbgF/U/aYo61T7V/pVQBfSQ67IDPdsQNSNO6s
STGO0KBF5SGpkk4lMEQLoYJREZ8ry3Quypm1aXUeNGaa2IDpA6rhscQEKXU1eRbk
8a2iM7pZXRPUcAuinHQynwiKJVTakW0ZAlCDxZH9RMS5T0H/QxPLIMQ2wkwt+PVD
H9+PxkjUpI2rVFSlz2gMOsk4UStZUOxac3GY2IAnXgC2Vsx97cgPlB344KEjhHN3
vkSwMsNMK1bInwzsVVzRblYD870GzNfrYJ95EAZRbDLjs1tXxZtOuaK/7szmIbwP
BeJZHrIt8MwyCDInDsZyjkB2sAokwdPDD+LJtVcxFikVzUsEr+Hmpzy0QzoH5TB0
lfLXLc8xnlzF7de8m+PrNI6rTgF7WJHmDVxG9dnukypErCjvcnKiIjmEqd6e2E2x
jdNfSuVdhEA6g5tdBLIIg6CPE43NW/PtuXKjRKvkCJ3pXt7LiIB7KMUvmqzYxw14
9ybLKfWVEITEaQ77w3G9eeA/EB65Bxube/rX1qkiHgeiFtH1L6nJXwfxpNPiGvVQ
J7fFSkGTEEydOO68+w8TfI72BC9jkaS45RQrAJHhpLVuWrJIlz9rm6sCQ/dmuHrN
xTNd512zyqrBJfFWBxRYqJ967MAvLfRk1OZZgCn7X/Pu2mmrhFw6E68BqtLA6TM1
PHn4yqlmhANj33mBYyLdqhKU/X7a8ioA3gdgRioovBP7TGr0VUc2tCtwc+6IBotC
s4Z8XkqU2NsboxtFCqy9LwCPgbkMpbWpcIV5LgFFqTKoZ2wPN+JTGzYEIVJ0BKu9
jktJAX0zUnfNPE/0TzwGmZcSdqvHRqBMN5BuXBEC4Kno9epSVZkZ9fG/zAYn6Br6
fKCLk7snjElc1W1FbxmBTcMIv/KzqP+jNkcAZ69ndVbN0H33HyT4lVsOSMFskq8/
ExaWwCdFLSF6xZkfwvBWNL4uhNWh2ykNd240zAI0LtjfOzlxlmn1AAk+W9bIrFuZ
rm8abFLbnTANxabKX2wXLKq2qytU1qC4efDjrdOjsJjY2ElSH0iDSOlZim3CmAaT
iv7Yzge+Vxn8lyQsLIr3DnHLWFOpnxtPxfMRemxWmARLetXrO+fofmRvJiKmWFbl
t93/S0tarcmtgzEjnZrmasLKo01ROk9ojDAWgKzuUQyvDNTb9IMsvbTiPhm9TGbU
Ejr634wipZNu9ipeHPua/j6LjhJESqIhHdbOeRXYOP3MqqEhIXsHC4g3OsIHdxiF
xkQwZi8Wrl1N6NOMrEqzJUhuB6k6I6S6geaWJd4y8B1C6MAfynLkRZA2eTo4JUh9
HoRMYfg7BAyDIUTXWWdfRtCtS9dfLAn8QpAi5Xk2vZRVIT3PeASWB8XLcPwRQe0/
ggh0ZQeDZfcpdtWylqnK0CAEa4dvJByq6j+IlmOdkxSoSsoQ4JEiqMaqbPcq96VH
hnsRod2Lqnzu9GSOtGwYWVz6QmF7petNt1UV/PLOgJrawaAJxeyFeJuErwoPPCo3
Od/j+78pMlnh4aJuQC4nuV52jp+7+6cICi9y5wJEjRZpIUp+RcRrGi1+dLCr28yi
+oHKVBPWJuHXtL+uvmkE4mccLpdUw8q27kqVaZbMWnIoPlrpYojzyWvNanYQQEFA
HjNdhAsJfzR6jgcENO1YhH18MhpxPocalUcnlZ6OGfrIH1hVGA3fIPjTJk+DlmAI
GpKqqGw1czHFCuUHDkPJ/vdKlAv1RpnqsFV0468aG75MY7mQEBl06JY17HqVSenU
0eNmixM08m12OUH7fJm5vGO9yD4SVd1Z5HsDRdNvEntKZxR93PLT+qiDRztD8VgF
NwUYzcc84rAsDkgMk0zKvgf7V1vq0ef0W1rvctZdDhTHsU6yfvWrv05J3Ym0XRK6
oeC7Uc6TtOXp5hzlIL1wT7dsgYXGLDnfrTjE1J1TrZZhVGKqVNZgubXhbt+Xn3Dy
ixCLJx4A2ivIXnJi+emQxyTjufnJCqGovNJM8lobRk4gRvF8Yi3b4JbiAh4rbWLC
UBtNROjtzzwu6fQYwdV25djQaw8hYhgwo7Hjloa+sHzI6DAudZ3ytDpsGZvkb8Cv
Oh0Z6O0l37nL8VjWhLxBh/PTsUcj2C1XvY8X8lV5RgwGKM4Pc9lUhMysuwEXdNp6
CtxmW88+w+ZKS1WYoWvEfrH22O48oos65w9BX4spawl3eoncYEbzOaeGe2OYNyED
0oHvbULcKtzrU/Kjz5WbazK6xYoLeFnE002yKR7foVlScxgDeWDDpfqRgpkXRZNj
vwsJkrmXyQRVHJymoWw62TowZK2wqNhwdRXR1dt16tQQohRel4yJe8yAucJXD79X
c5fOzGKog1BOPWQxdJt4hNORVeyhEip02QfkTNKPYizXSrzB2SiV0yn36N3oVTWw
klIq41xFv1tZZgUc4vxFUBXUArRBSW6OVNd9wW/WV9Dz4I5dH7iOglzyEOjeHCTP
iQGFnf8UnhqA20IUJ0zitq+XDO0qV9mlfH8uVGPkN09SSjdbGSnAXPuYAU83mQM1
Jsm5HjrvZb+Z+kISmvhRLiiTzmpv0eRISYRZ/H8kvEBu90KqrYBqejm01Dfgn8zx
sO9hEm1Y/uMWg0oQsA5JQNtgbzrLR4hB8VVZcacleDbmcVYzJFf9EKcUJ6R61wqx
/nEz48BHmIP31wiXPNQVrtVU2YTCFbBBNRpxpVi2L84s9jIdbNm4gSwkvuAV4Y79
qpw/0hIIlaPiM0rmy9GnTdgY+dmrRqM1S+3NoeusQcFVUEp2+etz6XUWbDcmTdIV
85cX1WFGMk2xji4WCgCpJPGAZ7AQdwDNX43crlZYMdJUJ2GO0RAXICssXHQI+yjU
2gJUh4sR6OrayKHtRtCL6Fb+yaII5p2j9HO+7HX3EPbbJjmBhcS/FttwzWThIPyU
aJFca2NEfjzL8M3vGUwyDkmgVdNfO+hUjgjCzbK/FA/weKL7oTGMLlfYLyVgquzI
dL/qACkq0NWkdmCNw0vc/t0cbPpE5c+U4F05Nl1QwMJr1SBojXNedIv1Nrww+hQg
DGMKSZHcGAoGMVMvfG57BQOPjRh/fkS5FV1rmsVFMEQHj1337JmO3DH8LR8aaPPZ
30BnbxobosoWzChnW/2TzQ0/Tw6MmKRGWYkCuHpTIwUkuu38ywmxj5laXQ6GQIWj
KtyWXAUOii480iSxJBlAYChr8ekSn/0XvXu8VSHM2PWeBXs+OlmfyacAYHzs8ks8
xESuZShnJlx1ATn9qEBII8r2zgU/B1KgZAhcrTWWwTC41oBF72TUv3P4iQZYciZT
uBE8Gp2X6OtOIfF6Xo5D4hCSGZvrQyhgeBmDP/UzbX3IXfDKYP75NE2ggr9DQTCn
UA4xU3SFuVwdQMGEY6LinYaolhM6/KPw8zm22SXIBX+oXG01hcLtJ8Xed4Zs17pg
aB9GaF+c4WbphuY3N9UX0NnpBMKkjIgk+T7bJq+PbqHKMrJP0Dgcori8hm/OoL0o
pwC1C8pcSCoeXJtC/g1BNO7L5sUmnTYDoEPVS2cQ94RcnPtGQTzYxnQ3FDhKbMA0
jYgj0eYoBOz5CjKm7mG8FJ8XbYyqCzz4BttJBGK1J0uH7HhIK/WiGe8x+s5Sz+Uq
HtiK85F6UcSs8KfUl7ACYubI4en5DGVGJ35cZC96e1FDj6XeVnZQCd9CD6y7nczm
S9NqWMAhmJ72oS1CE7V/uabh/yATApB7CLh2ZS2ifapLPzMzzqm3E6kMGZRwj7MW
RlfWwsG18RHHVb+fnGWZYM/TCcJ50L5c1w22x9JlD/Uda5zDNDidfBF83+7MqcZd
mUudEf3qWc9vbW9r8oc7LHfI5dpupVmgnbkk5yPk4nuD/OZsT55c15ybGPDn8z4d
q87C6eftmpHfm3YWwux6qR+H5iB68oK9QXiQzfKu0Y2pCAnZlLumMS+n6hu4AwH5
RZVbTcTDNM6R2lcPXj1bj3kV8chq6inCvTfhLmaTF5c0E9WF6XqMYU30fnSbQQnk
ymnTTmSzDHqkPfbPk5KbpdKKbJIRAqUUlB7ht51OTu/zkSMAjvb5oCr8y4FyQC08
+vpay/tT9OzqifF/sYphAJrqqgcwGsXTUiH63Ihp9IOKNgCN055i5vnh6XmGOKHG
IaSeoftlm68fkqTo4Sc6YyqD09EKqiAADTG/euBGlSYvI6vAJg6Ag9NiYyM9WAHh
XBIUmrjD/+JLZ8dlYXo25Y4TNqTTM+lYlUdXouAQlzaimD1FEslqjcI9dE623qhk
rp+nWx92f7co06YJf9YFYBjg6KvHspTEpA0MfbcezuqvBYoB+39UtR9sN3a5QAN9
PyYsA4TOz8WoFVWQYeiwHC6UgxqL7xRsyAVPVj1+woRF+GV7wFKcnYKy0rDo1Rbx
63IKdYyjdeQDuIsBSwjCmGTq/MsB9L2TbLxamnHMuY5+BNcn1kQk+CaEJUy5ZnTq
IYh8xDixfiIqfk0LLn0wttkTmhSJzIuTyNCpidqZzVGddFKxP1Qg7fZLAuIJD6Qa
WRKnpJwXNQwJe9md2kk3kUhWxpK0ZUoO4c2AecVDh9prXbjMdwvIIFG7JI1RUNwB
qLHVYOC/2xfwkDXc+qxqPIQqwj60Ya+Yjb7pcnWlgcjMYmk6HHhET7Zexcf3AMm8
zJggKlTiO4kMPTtEcE4GretdGeqCMTQMUcugb3E+cUg6xBEda3A2VFbhzVdg8brr
QIBNKuePYTdsKggD84Y35XFDX+oQoj1KPyMbIJZMJZEd8Su+TS7Rnyv8N3zNfKHD
SclZ7FV+KVCH6BUtYPUMfxRoBOrOi3qtFVKaCeOaV71eVzMy1hAuPsmZyJpJvqFD
aIfzWO+7Rw48V7rgIkKb3ZB8LgdBgiQ9xx3KD9Z4O2xj9nEMku/gFjQlDDWgdsu2
4mw8s98YTRCLgkE+mOX1TIQb5oz9HyRazOGRj6e/rf21YS0vt3byRD+YnHy8c7C1
yqyKxKqJTeP+HgEY00ELrsqbUYD9lZ97U6cGjAeq0rz9LexXyiucbB/SHqH3+UCx
Qe6iC3Teo/UYZqjpjK6QMmhesRrIW6/Kp3twNZaSeUfryk8q2D06DupVqTMxUyEE
15FmL8mq8N34gnIKd6s7XnGLygF6kOMyH1+H+ZsR+s0JCaa3YMcaEMWYaRHy+ufm
FuG0bOGzQUjRL8jcVDH/MnIzNDGaqdnDpoohZqmVz4jrHuhTeiCe09E7q80ApZ++
6WJ7UJ0NQB39KLd7oMcqWjgLzWDd7L8TPZCGW+jQc06voRbsKWf8+saJ+wChD0ol
loOM2l5du6rKTHpKeVEm1F90aK7h5HCKDcaoZjY1T5yOvdLoGVZzq7PJcBSjrNug
JqJz+amu54+ap2RpIrnMCkH3ry87i/THeebrvCQm4n4L+3DCJIQaGuiWw33TCBsA
kD0se2lnQeJpl0O+8kNzjrgg9yphvEiAyULFjph35qNt6bZDOKbWEI43uBdZlrIj
KxahugcpLG0ER51rAvRyZp8bA/mUsv8SSWc7Lp5FxvTZzD8ERXSFTouXj8ik8KIx
IUOXh7P0bLd8iMf+kA+Rr+9o+wtuMvx0pEf2RsNe7DkFMdBU3ak++KNmVgY4wK5H
6fwe9d07PNyc2vrcKAI9OItXJR/Xjxp2zPW6vuBEwIo4M6PeP/43raDQHiYUi6qg
+S0Y2l9siATe8HiK4QaVYXqkLI+NF4IK09ZDnXYMz9FvrHPkdXCLLocvMEMDW/K2
LByQO1NQIHoxIjoG7hVMTPcNjkHesHZtcm6XGJYrM161Rzakellfye2Kxk9xQNrt
Ej0ojW9IVzXNagTtOCTNwVTM36Sa5xeDHsOOf6hsV6cDSdCt8Pi/E6zimyfS5XNT
vvd+v40qhcON/67OdT0UapCNALAKXgUsFsoP03RsH/HOPPsN2G3v0wso2v9et19p
hc0zo1ab14YwRT3cagCy73OJYGl/jVFETBRdg2UJbscH06kPDT2sst1ER7Cs2gz3
HnZ1XBF6Vq6ygCMI/NzrpMwXFw45DUGIe9vl9uB8vgCvzcXBPT9k0YPE2t5jfwIz
QDMI+jqY7OUu4DxHk61nTUAgd1bTndpYuMo/nMmaLI9KLv6cp+K7vVrUXTaP7TFQ
bQ9r2NL5/+BqpA7iyVaIiYW9A8ktqJHgzHsZEpLQqIWuh6Vv764ohWBOwe/5TehN
bhNGsOZZK4kd4j5Sr8vWebuOqtMW3DdPVhuTwpgPYlISc8Mxek8EyDFNoT2TLQIF
8PnlAxzO+A/8tlEuS8XfvXvREUkNGXTL8dkl7KK+/PCSVW2kJwFeh7I1lQAuM6zq
uLysFfwlgkmUriehkjbK0jnYJOuEQ3075MAcKP3IxfbCn8e/QGwsTGbfGyBbgk5y
W2qzrcLLI14HZT0p75e/ZDYu8kfA4uHZ7YSmy3+XGOoQ0p1EBLT/AN/ETSax+SCk
tCJGEz5CS1rh5pEKnBNC+HFhzhQ3Y8iRhkls7mUMG1rXI+kUF+tqMlycg/Lcgi7D
MaDczi+2zVRd9n6y/vXOjPjwn9SeZoNbjpEbfsUEc0ZZ19OqI6G6VzcOOjJ3qBSF
+DNW2YXnx1T1Eo9ltzoVmdvyZ2UdXmQpTnc4s/hSS4rehNDufeCzov5Ze4rA4kj8
Ic5DbInKR8w4i+pxk9eVMe9qVfEXs9t9vanbLgiV1SDPBeh9Y+H3Zi5zbTWPDdYM
DO1eiD/44pUIsBHRDPlOwemYNrEYwhEo5HwhliJZrXNjKYKJuU3rI5KuakWLaxWA
Fg9Ko1TnfgotQgnRvUHJVB8BW9/4bkvBHlm0vDBboZUucy5noWGsS6H4wI1YKIGE
Ynmy1m9nokEyjBwREFcp92j01rWDUiFC4WiEtObyBaVUqbrXPErwEn1b1cUEZNCu
5BRe1N82iwGiuIsqi7Rt8tURaX9y14iiemana63+mVY8AVvaOIxu6WRb4JDV0IkK
d9KICIqpbBWoZniLTlZ0LcyRUVZfcdNaIlkjov/V5bsWCKApHFodh1bYNPySc6vl
mhHU1J++MQZPAuEWHvjIt/rE4FV3jL20bGqF4g5Z930qyYJ3xl/DzESLiBCpT2wr
VD6y6JmXtxMcepxf62c3dRMMeGNtedg5KpKF1Zpia+5L26jFujucURDsXAFLcpRr
evdr8tOgL0d+9uSVbUxCxCWq4st33xkQRkMPLDhOSnWs63R2Up88BxOaeK5iMqeZ
ZfyvW/fpah94ZwqqS4NSX42d8GGdzYgZ3AYOh0rAxgHSRNvLGjr5cjJtK/XCwntQ
w6lXKKeIaMlLF9vhJtLw5Qr83aNWqDm4wyrskLy07j6DBuxD4XpVZhxik8+Pp7Qz
UPR5I8m08muMy59q6GzmOqVTRpWSbm5yc72RFW6ldkDrR080t50LupbIKVlX7qY2
cI527eE7nCtg2aV4mLlve7vwDFK1grdAD59Sw+z/Gk8Qa4azHhiF15lJoIG6KdzL
CtXw2UjlP7PaCcKc/sMakyVu03GYECZWaiwE1qcsRmXw19ikg4+wpLnzf+VwUJSn
xiRSlNsWaDBQ73AIlZ+oZXI2L0RzTQLPxQOPpjFGtNaqj5swBiX5OgpEI6FV2uMa
+UtwcTQ/Zi1AIFSFM22d0GiTSoTYkIQuS/UGWBUVRwW++V09UezHGgSsLr/UFRiX
0vleA1OjatFczTz8Omba19XyrHWWleMe+9SdqLPJnyGq1/U6HhStaQrVONGJCs3X
aX9t1097KDmPrnjKh4kjZz+5+q5QMI2un3udi57oloEGuSnwlC5FwhEzyeQCmaGn
DZKKITFz6ZQyrfV/gW+3/Uz2imEhSEb3z/nAOI+fBNUAN/mCx456RJJaEW0PkMD7
r0ikp7DC9/PHmBF8106o1LScLTY9Xj8Fn6q0gnhjBrcFgaWIFXjCbgUMiLoz0iVp
sIgSd3uEOGs5VpqsBd6NhZa/u/kmZvhiz+whlwq8PVO5wEvuYOHqOT+JfWRRHmRq
glGUPLKhxgBLIGOM/2qulm5bfDfyVwX35nTOZwmRBzLrQ31aGqgWQH66235Bnmbh
M3Xh+utZUrupFwA+Jp767EoUkhxgwCIZGkI4YojaO2s0xdik+M5HmM3iPrTI/tdc
TYIkBbkOiswrmvqTGXnNT8RQI9zRDCP8nf6gf4Lyi+wdtfHikhUhXxwQsjtM6vUK
70qgcPDEieyVYYEIX43NuzfiJfZAtmzROpgOQDvM4XbZWIVrubjfPVA8hoGe5coG
0Ye0+hJ7tg5XILB2T9omXdH+bCPrI0ME+YxjYXsfFtKQFIPkmFiP9fJl3MuVq7Ou
3KDOsWwH+guCMV6VNALo30+Hlw8ST42rBhWhPbd9FUPS8xa5ZWNJ++TtjJWOY/Ay
UOXtrBRhuigZXJAwdLDDxAw8191aU7k3xJSn63FEDNb0HEG1B/YWq/G1foLoyrIk
GHocjU4lJ1K47Psu3S1Zxp058AdVF9/a2wdz3u1I7aZ3oJ/xnKohsSL6R9UykHDF
CbDKnBeupkggR0KSvjzjM15dVPQ1Pi6ThUVxAQxCgIGhJPPVM523/REhymlpR7gu
cAFkUeLLtC1CgUv3xn2naTScdJ2IoOv4xNhmEW98an+FwXlOZeetIeC6fsHZro3p
RtXSzx/+bzaTWogelyKy+mzjrENn3T73fBHwdqQT6jzzrMankTzRzHDeSIYphi9S
WgjnzjIWcKqLGIrftevuYtxRf2JkdsAlVVQJZH4uBNxy6OOo+nsXOtV993A9XHIH
Epy5f2fFIV4MoL7Om3lf08Hnd3WEZ3Py9yLIp48ioCzOg9X1uW3pfsFIgO1zxnKy
jy1WwBDW135hgT2hvdxNUIkAHQW1q0BrTH+ODgCib/lGom58oI7kaOEWDiXrxTMh
j/MROI5j2j2xOdwXYzI80iwMom21q711gfiLPQqDTLLqwxL4h08nkD/9S2Zxxr5f
oP+5pwrDg0q4ERBbHCgQLWqTbhjAnGmnuVFhoSrwWsv0msZ9PbUkIpySyuSqtvcl
Cj4s5zDoC3T3x+hzaOtG6Tl1wg1Farh17QJ9J+2Ufa5W7c8xFOhRNsqeDY2ggm0O
cWwBQm2w5ggdSovl5ulmhWRolSKJ8hDs/JE4M2AlTDU2h9t/SOfTfNkbZOEL4UUC
1gWm7vyvDzawtmhiz/pPhvHJN9frfLO55JRbhqk2HiP1AXScOA2T7T0+5nRLKFj4
E+KrK+U34SFIa4sVCfIZ6IJ+rzh0CQSeKhQk/1R2AmCgE+QLyHs2yzlDEvf299se
zfDxt7Qp+CVgAI4mbwrE6uj/jCNIxsA/lztVKZlqWrA3vxmwemkfMIZ285qIv+LC
edLCN3ff/XNMpKii30jTxa13GJOhJLgFQeaHDzmJWZDkKrlxk5NgRwR571hSUBF+
tea3n6fIHc/cV5GyCwB9gvp8y+6FmG6RtoRB2pgc676LqrNtgHLuHqx2IHylFF1A
PO9w3RyWOefHI9WNmvKtibEHVpyPqMIrJ5OlawyWQ6nCOQGU4Ktx7v78tBkwk2in
NnV8KD0FCYvgXD84uQlqbifFX1KSNAqc43nBt3LEoQWIUldkdboozVf4U6H3idHo
YNkKTIS6Br3iDm++/muVCsXC2ZSw7rnsUiDG2iev9hbzivGYCK4bMoIphLqaMKUP
R92hiTYr6cLW/JWn/5oIidpu3bbV+xHDQOAqMWcJULaY7JSEQUNjcPyT4xTjGAle
U0Mvda3bsKiLX/O7Z2upYMuBrMrJxcoWlPPfTVJ4s+nww7oUqrJEZMNCo7O21EQQ
5k8cBrgQVtqi26RMspS5p0QDM16FU1CXO3y6fDoDELJCRhbAd0LOfIO5cUAYltSp
3nrAnqA5I48PGGGGDBjOcfQ9D4LJmG8RXYv/jjgyvQ9bHBhZ1R0TsMdABUMetHBK
LNNgH1zhtQi+QyjfwgnMGcdjcFFlpLs2dYnXr5i1iwVYFmrO3t0vG5FtM0sgKqm3
tBHbHO6RedGE8R5YetnZaoLOTCAymG1X5gixE8BZXP3p0VDfhNt1xKITyFYaDq7a
WggZlAuBszNlZM0/8qMbjpLjEoA3wLBmoqUek0f2hN4+QVROWYeR0obznl8rDMcE
/+IJ2oEOZu+6jYEWeEJt+uniK1Kesyndf/UOq1dQps75qkLN/hyZ6yuE520+oml5
TmDjq7/coZHyfdTA7WvDOtAuX3Suf2vjY5v/wIlqHxCLy1w7+p2oBHexB1Z1B+kE
2uiKL8cGX4ZKkbvu+P62JP0jgjFlFjgtUdZGfdP1Yd9680IX6Xe/gWVEODHZeuNF
CT5y1HEzxrQr0jCWsLaRPTUa/aj27l8pIWAk4BnHamXaYAfxNGPMP7GoTCNprDZa
71Un7JxVw4Kumiyl9b8o+iF36ZnEjaEeNyJYCcxjWKhUnJYP/a2ldcYeaItd49sb
YTaK0sXayJk0Vg4njE55TEQIl5aoUNiimkRiGm4K9GnP6jmhez5XCliI9h/XkKqe
iOfnF36v4AAcDineAzdp8Hh+XkO4fHxoCtPHRgDhVKaI3jNojFDTK95Dk9Ig9n2C
K0ISWyEarM+A/rwqVVy04XpNSN/+9epEE5s2rAjtekiwzA9pxuhc/op/t7Iy2O3Y
7hEa1rQ85StAYb9fwDUqwoYxqK4JK6+bR7PSgWczAOsDvHqLtSgAzMhJPs5vXN3Q
Yo5HV/h1mwNFYu74au+zi3kp5FsEzHRKGAHsSgoTDcTosB9lNYayIKJWI0jWevUm
ri+ltLHZO31U8S6917aCYiReIkyensXMsZ7vgIBVBre3I1WRd52YdrSVEUeaNUky
aS+wxj1pRxZ8NIdhefLf2Qf6k3y7WvAp/fl+MPQ5JuAPiUbgUGIYCr5deSvs5Q9+
HBodQ0MxWQ8USMZ+hLBncBxASXrTQwKob2his5hGPSlqVP1a6grBp1MnlVHATlul
606Mdw0P3RuSOYc6MuS7z6CsnKGSYNyrQVheeWNl2dcy2hcZrNflfANdE6+MyefY
Ic6ZWH40niXq9pIVZunMqXZ+r7C1Adp5cEeKz4nXZuUKjADCqDboSd84lsY/d61q
f9otklUsAvc6NuALX185hLFcg4Rwaui73w7mWlwlkDvUA4dv7fHAtAJESMBpVl34
9DGefTPOrvXI7/G3rVrXQ/GxDvdjp2IJEPZJOBuY22sjg2Bs4L6rodPhSZ1e4+9r
LnNCB3KYFHx+F26Ss0YCO5IkH/MZ8WORybdcURhxK2b9U9QWDz7qxK3wMzmN1rEQ
/Eu7UPJXD4t6OpoVtkWc/vYWvlJVR9a3zAafwmjeRMwoWmiPXLt3ns6KfDFW+Uj+
NV0F7raA5JJ2EeEiSZQqONcDiwNiSedULVNQ+oc4wDuKItqjHXdZRiUwscHsDU68
E/UXheqa/aHZ7pnkCB06yJuPLh3bPXmOXRpaT3i5JcGuM7sLlFJgaZo5efUw6QTt
iILoXkCiV25GyNE9p3fqbI+VXNUszpLtRwwSwUYwWmbjXq252Me/Dv8BW2LApuJ1
qrZzMkm3Zn/R0BA/Tl1aZHzopJE2bPpUiPwH03c2qnmKZtFIGqK9JB15LhkJRtpB
7D8FXrpV3rz+x0ZQWY6SzH5wwllDp5V/ehtHmaKhEbLpkHzng9SeqtkntRR+BtGk
wLvVqpQWdd2tzz2NyS/EkSETUevMK28u+80gETnSs9B1OxskUL1sWWSpTl8DS5jt
43J7mPurTo4q8MRxRl6+rTTiLpKgj2lVotdlBTNV2Rz51q39P7iZjKReZ1YlUeKA
gfy6kZHLhayCtmccDJ994yCmVw+e5I+qFIjqJLtGPCApSrLUs43j9Adse+XGAadI
Q5KEB0MX2ujGTgHvrFyIboTq0IXzaitogzxLQnNgcjkzqwhe2KI3wmgZtpUZ1krx
xS+Fo9zmJb6E1HI4m29bE2DGx9aa4g+tY2Wl4lnuldN4sQVIOsLYqYde3Eng9Fd8
w7eh9P9U2sr2I2EjwE29C3wouAvxQuKj1JdtgCd2itxK2lD0IPfZRlt+OE4W8PWO
4cVVnCCm+11BAxvDHtBy/NIwUmLpEmkxopaFoFovogQlkcQ2sRM2ADk3cojh2U+L
V5dIrsLvq8cUvBBQB7ipRGya5/3mVVXFGnjEug37UoW75F/HNiXYmMOhStGYAzr1
WqGo5pf7O0TDXksFlDaacokijlSyqeXJ6dMMkN3x044fNiB3TfHGki0jaHzS+fPT
DvYjKMvxS5bU08hF7LpacXM+pXOSx+aQWP78MpxQK6pl4rCKGKY0Zun0agk3uYQo
22yCrw5YGc3wZqhkx1Q8AqAHFIVtEqVu9+PAO+tL+bNVoVuKW0TR9eUEWuSzhvgY
pBF8479L2AwS3id/thN5ogcPQgj/uDlqe7ScVEVz09EWSNeH1TAwUBU5rykSC24u
0pbi3Q4bf75SJZIQzrwgmvmh+wqhG2wkG9lmre73j6KKHapvrETOocwFBi6uNacv
u/4X6qrixxcYKlMLpv+6UKSmxGFJRo5Iru6DpfYteyuctoOTPOkv9d17kr5RDxiU
i8V45oFP9maULGjXThw3CB0kCOUb16MRUShvcA5s1d2V1KUFHh9ZY9VAAR6cz1xh
yr/ojfFQX0SiHTxVzffJZHftibiqyE0q4GOCpWBvP6rnskKwdtCjHzmsDqgEkyr2
nEMe7s3y1ED0p6+nIoMC4bTtroYoB+G49hdCfMy6Zs+ZW0Q9uMyqB9OjFZ01LUKK
RZkb5c8IXWAqcYd/d/zX+fNr0JiRPJmj2W31cticnHGKuHP6DHBwE8qg3hPTnIoh
DFvO1HBKwVi37YpzIX3shzldJqnSuICDVXwpyeNBxZt45gseedomxqjMUIZEe8eB
dxi2VXDjc+43HxstCM7f75iLWqQhju9uUO1C6v5+GupX2FJhFmfcvVRaLtBCebx7
mMGgcIMBkPiXkNOB/OKH3LJpXuEt7/T5o9C3goCfnQO/DP2fUdaPqFQhGmliCyLE
dXf1MUumNNEqJzJHjhF//zU6xdBsOjY3osSEOBEap2x1Si1dJBGCb20rX8+6U3co
C0kzc7qPliZ7xWdjMub/HyymF9yeGEFJ6u0vl8H2fLKUBk2rBoYoJ27khXkR4Cwk
LzFHhhD0TAPNDJ0zq1UFvtLnFz7fsfjq/VQEOork+zHOnzMilBPAKX3qxMT0mdPN
tIWM0OIECOzG7eaTp4TINXEnUHy6h1tVz8TZ2oe9TbrBhMoqH1V7OlGQNlaMn4Gm
/6pF+H1DuCcRQz0Vl2q7vQ7W9N27uZqW9cwi5ugOGabIO+7Yp6IzUG78Q+Xu15ZT
dYn4DYs7RAtYE6YdIdgH77nioZfzADhFmuzbid/147RKg/OWDO8QzV2DUW/CP8do
l/D4dnyrnxYOfaBnVen9zwymFJk8EgHjkR+0OiSZsge/e1uNXjjYl1KoB7FYiG1m
ORnUmYXsvgxfwgZCVQrItcmqoXPFEv16+66HKHpf4xe9qQpNZIbCOClIdTbJ1ors
EWh0A0BNq4NOhuNsjWU3KLAZhu8CNEGkLNiBJy/RLsbiIeuEJ6GsGvq4j2G9bP4c
KNJwWHvAJat5FnBniW69p1LXomP6gcOlINZmscNWQjUVBFYawdTl4y5kvMMf8U7c
uyR0982hxvVycG2SA24+WbdkFi/WGNKusTBqrG+KjWvYgxMrn8m9fNZ5K2MSHsEO
/O2m+7umo3VTFUpv8f0j2nH/uhhfY5h7VkLF9dhhd4YEMEorJWIA4o9TL2j5EdSX
QbB2Flt12tqUFKcUDWr4gSReV4pK4gYqJaH6HRZ0MVw3G+56IVevl4TXTJZmNpSD
0jKOQEDlysxM5Mhoq+M22sIfyMFSUeLpSPU5KDp85syZSDOaqrGEEO5QpbyiYFxo
5EDkwZJNXBDK+coD+vqIv1WHuzlwxbAxW2UmrtBG6AWWqEkSCgfxM77NM5UpGsdV
m6J5i7hCzzs7gUmvYuQ0lOXYt0yldGhdbAOe1pJSGvn+hcCm9p0Yl06vtkBNQz3P
+/BkXYaxqC5XUjBWtxK0fS7Im7j68TcdVmsLC1dvtO4WAZ5wJn2D2t2tPheec2IG
3lm99Lptb/NdEoYzCCrOYtg3meXH6/iEWXBWT7bszq6aC9d2pq9tjazQgHV6DzJ+
emRm2yrcBL2UadXjuYosfnPTNPNOXyXiC/CDWJMET+YlKpXetYjHCw/07qjZdJkW
GYWn74a6Lpm7xjgSUiL5ZENKh2DC/5qOD5pFfJT4y1njvAtzwn+9S5OvL1xWt4/z
0FVKKBoz1Bh5ogZzTTBXkh5F1fAUtQb+XpqJGLdWgcqEJiwRNDrbH2wUxiHB1aqO
SloRFj8IXKdL8BwvWXIYitWwlAn9dupv+EaiJLFhfdqzutvLfQpB4+HJDiVvMrJ+
Uv+lq15bieuqw9LbkO5WEvZP05LPHA/pDk0StJXprChO08+voN/P1S4Wo0gv21nt
p0hR+uQ43OVI3Ih05Bhh1tuzZGCmJH6wybPdqP0/U1KwXqa40+AlnXitVePD4ilF
6ORO65uTWxmYJ/p9jNRKsHA27xHRbfExIx+j13SEznSibM5ITptpe7KAXmKtUcDA
02FURxTaOhi6OknFtH6qcN9vb3LGA4TZu8IYEzIYXPSQ9m3lTZhvCnBSUdX2cIqJ
ZIUo2LcGShanw8DlqhNd5nNkwjfLsSQGQCrZci2xZjJts8BBlDSoMxEgUDhbg17D
ijHfDjNE1JWBRAecla3LIAFR3PCVHaF/MrR+7d09DIWSbIrvBQbIGgSXOzrK79kV
XwmzmRyr25wBQzBmy13+fPXP2CIdSTqz19Xb5S5i5ALOURWZjvIQQg3qLwqK7yTn
l19UhXaMUkUZ98Boy8R6uV6NcCOfJy9wnw0suWbKD5NCm4mAK/kZLXubgL91ALkY
SzswfWsAiOfN/2fAmzCRki6QoiyGxyB2pWt2XOzSWbURHZ5vXrvXO9OKZYMf/bHm
vE7OUlmMP3MynJL45B2UJdegT0YW0MOBZV3YDll0TdV85v52N32ffKJtWyDamvrc
ZWCoxBcThEUQdIcFWyYSNzLpZw6wYFHNXJ8S85gXE5j3ezbWJHrN1LwVHuNGZiWL
WPLJSeAht1FlFSmRNP/Eut75rqrELAniHBtxmD3LV41op/POiQ20Xe9ZNhP+YW+b
XM7eG96ypCTYjZooWwQbg79Z5rVMgrLPmAsFgLjrTbmQpniXZvE+zJvyzK1Tmxlf
X13lDdWtfqpVSzu2B5RzvWDu9Ultn+i1xi07pGU3VLVPw8aQDePdm4XgxVsxhGnh
fwwspyWcPQeaYfOl5cAGLkqD0Ejk67h9WwbDG80Ek8Qtv58JuzD/ohxUSU3iN0PN
ZKuRicFsIzha+GmdspXwWBpeshKWcusDOeSam6yjAOk/hTRjGyWjtN7RhtWirdxF
zaJKEkvyfc54eD69hkM4UpaGFsmHoaQHe5CyZ6+7BN1sgjTXBoSxdWLZkQ9w/r2s
19g2uy2c85q1wonRuW/dG/qxt/xktYRJbi2c6gGbzXJULMHA+R8h/Ws++qlSgoo1
srcuTsAtcWa1EFgCXgimolR0BlFec0S3XTBgAftfaU7vZs+w9CLvD24LItkt45vU
2SSjUgiaZKyWsUQezQrXQKazhndgIbAMo5JrYzTNMoBtGkfeaiCu/K4r3vEwVWsz
J6b5lDt+iJNA2JS0/kDoJNKSsLXu0NlS8qQpbIX50h+NJ+Npo+cg6DgG+sktZOUQ
vw6YHtmdcw5a50uVCSckS747tMVJyjP3ZFJYv8ZEGSOHjhAPn4XF2n/4pxRLhAfN
JtAINMW3ebvoJRCWjkAYyDXmmUEAd+EpdbjQT7nRq7FQDSpZIN93F7Jc5EjGPq5/
Axbi21sQG1vGvU0LocPTokj8zGFy6lHoVOpt/LW+XIMG7rYbCedGHHq5+L/Vb9nl
z6WAqPaOuLC+zwM5cI9Ovcb6iw8UxZD8qiB4bT53MnvVsVfHQbykFyXYClbF2Kdy
QNmGVxEWPTGRdaAbP3uyknHQ+j7A4xSs7mhOMZKmTE0jBctxg/tcBrErGF4OxJh+
Y7/cgiDzQg4Ku8J9dO068tz63FTimV4Q/yvIMU1CQGFuKXID0ag9v7oSMnBMk/HJ
3pbADQlv6nCw8I5ibAT6JPo/mjgOBaAmoxWwK4g3rsCj+N0Q61GtAX+mErwWjbZv
Nxfk5Uf+7wTilFZVfKqhFX8kHF9a7NEZjfE5ZPWjKGiRv82IwC4AA+4U7eUh6bTa
u+Qi++3f1C+osZ0rJzya1jKGKFvQ1Ee8NpAeNQ+hiBxk2KIDk6w9x65sYrJ5vmkV
SWXP2OE896btZVD3AIJmS7gbP9JvDPazM5Nv0p9ZxyKR7dUJvaK1SbnJan/EDFyk
SyfZ/XAmEk1bQShWK22lL3BHXgMQTAavQ29XH5nMj3ARWsBe/9LYA+SKP1fbxxpb
Sy1omEY/BsyU+JbQac3p/lgwpZr881ln8Mk+B3Bx7NEU68AmNdqku0elcd/6syoV
xNKA0vs4pzfzodJxYqnfS6WlCJ6z9pNayASP1Z4b1lRrfei2z6+xQhigfuD+mGrH
wHIwq8/obtG96gf4kyC/utSdFKRn7DerAML7jWvyU8yDOfhctPx0LiyV8OIGqH+O
oM5LRc+BaNA8kSyOEPOWRAiivWhXB2S0ma9CgQGvFulvpH5koi+W1G/cBw4qKXja
Cb1L0wMg+dLjsYHAtjVJEiqid55QmnTuekFoJplrJmpFAe1Yj6afcBbuTFAm3HgH
W/hcs62CSG6GMX7vQjXpyS0WPBYS53lHFt3eAITBpcI+gaE0fcobTymesCXh2HmG
Glij8zHpaNKrzVTwrjaYOtEtlEBXkFOXcEVkkAoZ4HSGM/D0F8pavAzp126RXhJW
c/Q6p8EAyaseAe71oGIWOSf+8WYcjBtoznRYtXf+BCS6FcUHt58FfIQySeKHG0NV
b+7Tt+ZnIBDEdKPWgh3GGNKTHE/maZHs82x1N08IX3thTTpV/ufKx65vBd25Jbzz
QZrP+jI1rIMhiIG9DoqDJvS/cuvbiLcvBT2CGbSW+RCD0VPu35r2dxeBlbRRI4HF
IxmWIJpWEwiVndbmno6ABRFORYpJE3niRanMwBRAQTqxUx+AspC5LwTqJCHxdHDb
L8i+U6pUZM2pUA7Y6kiFdrZGiatoZkgWu7+5ZlFkTsUb+FeUM6DuKRT89q3Iqa42
JE2uf81QUy8u+ZPUsF5nZR1Wr8/NoYZEwc9cgmZeXeQhKwQteuji34Yndn/qgIp7
RVXb3IeqbEDrPa00OH8FsuwXs0Bn7pgGqY93qkI/xUHKHMWaCHJAGOTlWegwYs7y
q9E7MfDiiFoVbrU6PMSww1z+x1h6EIdPdZAr0ZOC7bKc4rVgRh/c4alOsTGd2xHI
bbW1ZJnHOrSN/yAAaBua8MMrRbyAHMVgU+0y+8D4mjb1FxzeQJcmb4FOFIdvIJ1V
wb6MlVNIidNZcfMmtH24LDIel6am+eTEDuHIAkJChtuN9lvqANvHFR2eo72ApO5x
zo8Bqwc9vmigyrOl1F6T1i6hF+coXEo77CCfr6LMXlQyBdQs57s2pd2gxdnQemFB
0Vaj1epaoyX9wlby2H+aPT4XJNXyNIcOD+nz/19Ds5c+B5G1tnyHoyjXEHnCUwQ4
iiC9ao/8gcWYFqbi2Hwmjcqq3VTtP2rirh3+D4gXK1mkOv5Doz7AMOHjokqNMEZC
Egk6+Hn7EIMu/bmDBAFr1+ZiNOwwzfYfOgl5gSVeshTQkYh+DM8SRiTJCwVrtrCO
goLJdYVZErR8gxMy6+ZGCFhGo1Gu47asXnndzSdUa1lDwOOELcmdtcf9zv2C7hUh
/yqdiTqy0P9GcNeJleXR7IsLEU+n2Qscc//SpYwcnfUsEfAnSESlfYgTmsn2gTqm
IDmkjoKIuo+vtsVgNQVdPa20Kf/p8N99urPUliTc/MDkJZyZKM97ATBGMwBPaQot
Gn2Q1o6P1oxydnU9/MMAKf4IJn+ruZRmWvTOg/AW6eFZptGvmvOZ+GuFDsSw2xY0
VCdyY/h2t4Y/ZEDFgwW56GMKUrQSigy6drpNDyD+57ZINUFVh1VhU+V4kqFW8j8Q
neBB7hx6Vci7+Y6WJx3bLwr/usM3hBf3wdOA5HgA6obeniCfFlZ/KzT94QhEpmz6
5mxx/lS/Rk/5btD41SHluJfgbONISqBwQxBwQjx4mwUDnvzvfGmgdzwfN6jT5kA5
xUvqGl/6dnuyhSycpWME+AI5zaOKrKSxRSR3lvxMsv5iCsTjUJEeTeOMuQcm2Y17
gMeFWzdBF1PuDohMB16g9mXCIwJf8/X9dJcqURZXGMjG+xY71UpNow+Pn5czt5zb
TZvTKWCtoXp90RbOeUUbt7C8sN34Eugx0c8uC3F8phMR9FZJPBmbu0JpQb2/VjgY
oZOhvdd6TtxwE/t2qJFKkwo+KagmLcJFIHfZOe1GB/c6RnVk/EV0e2bnERShTz+5
LtA3dUzNnGbCGoaZ544WQhoOvL5oFbj8RkLhVMzKzGmgJQzdWQQWKb0xLDINynJy
c7IgfgO34szuyWdMFaXuD0/0qkvVNJn4Mqev9PhbnYxlk0RJA7WsEyiDoGRvflWl
3hLN7+Kk74m8t10QfcV7AMW8wpeJGfGknU7/9eSxutGkrdp6N06K6O33WP1zItjv
3RmAJUs3VSKUNER+ooGYIFS0O8dNG9oVtcROt0xc+7RQ3jMY2Cv3mhguCf0A9anm
hE5CR2kmZPiNxbXi3nTRgy8Y87vHZaNmH0OkjIwt/QkxK3RvYImHmX1e3tAj/GRH
OSrTbLq4uMb08JLIsgJHrjkc16s6vEtumt7mPrjMT69xGJFXR+gpp3ad4r9+Sq2s
NUhgmCylF68rUluJ02hQwtL+X8dwk0mDk1O3w2F1KHuDHqRKcWlA0ALSke1aP03W
XKm/O1pv+TQPpx1oLG/JPgcA+r8ZopTH0kZz9K6evLlOv6qYqWLAcJdJhAPOeKgM
hVDwvnrDAM2BKCMjzYDB6JGyIGs/C9bwB527+EoInBkYVNPbVa+tOhEZEYhHevcv
dw4d6MqeFi8mt/Y6vlWAkNsFsyJ4+dz49qRqTAf7DWs2swkmncTRQO/al7FUFk0C
EM64i41dRn9f7nyFOQH+dhys1+TgiUFyxmSIYC+Ddnt/JALpsVbo8qpg+6BVfouC
aiy+pt3K4oMWNJy4qkW7ulfAb+vdy+Lfi0HCoqT2a1hD4c+J9YA5aPX92UlWB8J5
pU4qM/fNRODQ+16/H2yejDhuw77yKY4J4Shd93+j/HjhUhJYX6cYjyDRIm4vKBKy
son1wju0+tD0W9JCGCDJ2hV/XKOnMYwjlu9r+bFBsaeqjuNxrJZOrjpR1yWAYBRn
nANvWRRoZnHMdHcqgyr/7IaD+sXzaRuJYY/Q7gSe4q9KYqRiXC9N4UDHmNVirOpQ
2owDBZwxpilsRggydlDdFn9p9wXwLhEIH4RO+FGd8VvavzSLMGSLSYTR3dVB/ReN
WaSQUYLbAIXP3PPSZXkM9b+parSHiPCu6ZKvWZIEjDFF9HcSo/c4K0G4c33AW8Xr
1//RXHNrDsjtFfqWHlzfdvQrxrqudMYKAFdkyo5WyX/shDsKmoECt4gU7qVRr1+U
ebiHrpYvekQeZBkx0O15XvoD7ZcGCokBMjcuRqjlOsNOtPFgw30ZMJTK9G7LK18m
HKoN6+XsAibpzJN8sUcUhlvNP4gs3pDV1eJ+wen6hrgkNN+Mt9leteGU/X7AE2aS
4vmOsNYL0kz9u2oJptI7WrDgzKUViVFprtIP0AYraYMhfhc4Gu2cCHhcdN6EV6TH
9kQonckjnoTBjKLGatYUN5k22Ih/GQVLCPA5by1I83lZ/ws0StSK0YX8QWjuOYDX
PwgOFthS9+Z35CDYs6JVW55OnJCTaHJ9blxv7Ffj5MVGWpc8Xq0r2s+ykJMukj5m
skosEPuS+nJFVcM9KTVgtJBeQtqN/ysunko5MDj+veXenwIo2tD15cLyzxVaLw4s
VpHs+t6NQBGbzvAOsARKryemCyS8sPCkH6hlIPhYsE3KQIOY1ZqgG17p1lzIVid0
6kEp4c0QDhwvp5nOq+h67eNeOxMHjQkNIUYuXco/UYox6ayFfQfMVOnbm1q4D5LO
deVBBKIAY8nMhQ62cTVpmk7TDU32S1WdNxDJqoU1xTD/HorcC7Kuaoyx1E0voS6d
zTuCjcTSlmniaVjjNNwenymf2f6m7mqi6eo/Z2OQPYGkvenF2M+w+EJHtTMwzcC1
Ie1T1H5o9KJy5Sp2l6ChXK5P37OuVudv3jsRt+uVdgb1wRscJTFgQkKdC6dAJJ+f
aiubEdwh4iXg/YyNbxnPcQJV5yxNQJ6Xh1JcmsY2vNsw46oXIHwJtMU7bi3kwsb7
hHcpwOassWaMZTVOlz0j/1HJApKA5qDT34z3P6PftN+ZLrivGo46MRG+FQ7RvxXc
g3yBF+KPsInIA3zv3Hch3QSM9zkLdyVDc+V56tB4LAc327jsSsGnGb49iBMd53dc
lcs71QblTc5fABINraSud8oWuxTZbbrY8uGNmuSkSpG6pm7aOB5iCibful/u7xv/
xoU/62EFf/R7bogceCckH6S0RiouYE9SRKoRTOa7KSpVaMxfnBnjeKeDuK7gt6jY
UbouCcezWnDfa/SBMU5ukBcoEjLrPBCvAKq9JdKRDFDX5s4L4yYhwfppFnqmayHy
r6eBRNsyII1ySTuzOCloWsMyMoywppgaGxTMVKeTwbhvsGGBa9qKXcbk9tTfRFfG
NuIa3CekADGhKOVr5hsCQ/PuF8Dmto8rDm+1mmVDZNv1GC8nVvWD2TsRvOMTcdYW
IK7CEdg73gFCZTquv3xDzM0Di6fLFMmW8ZZMLnqgP8Hry2f5JT4s3ah7JYZlQSGV
eIuDxab0AoOLtsJVkfJ7RDPCdXbnZzcwYm3mwMf8aM5YQViknZIe2GGaGsjnVyCP
tNrboXaT0G8OW0dH4w0vsP5Ravxm9v5k6vGQjCmf7RqqvvIZZerMDaF/pR9SJ/TM
KG6IsA/XRKcYWbHEpeVUxLmLnXG4j54DXTwfM5N9gQTZgD2BwNbvwECyf+E0KYkt
9dblpWLo4ISUcVIUI2mCjMsWbDaZQycBVeZ59gRvRziLMrU9SB0mp1jRsuPkHDvG
WRbLu4iaqZTpsrOxMsgbBqc7Js32ofBqMVF/QLWGdhE53U0X9McQJ0RCUr+fNPn7
x1wbOzd+/Ro6cov0jh5cJRNgxhUqkDoZVJR1yzhyIN8Nkjl98SHXggVxeAA6C5He
YvP3KDZ1u+uy1ytwTeGdLTpPrjQHU8P7jch8cykNbvZcWO8g1zBPxRNcxRinzcr7
lmXiukeCLo3NYiEUKSVPUg/WpYsidp4w9Sc6HtBwr9AFAdJSwvb2d2aZFwj+qZgy
rBAm2CP8Hss9AbuKjVbjXiZRavwVBmtJuKFJ/wdafWnZlH3/Sa/HyPF2d8XkqnDR
AjixRaTcSzpNJbfMmqeB2CFTHh2TfRJSBZXDcEBZ6kHCFn2MoUyG+x3zsLvg4xX6
1Fn5hRVWynAMiWDIBLA40Cwb+pToZ0BCXDxR2g82DQuwCWA+dZ/PNizWbL4nu0kc
6d30CT7Kwpa4Cwq8cAUPPLZPWaHltv0GfeWVZiTUB1JePxUSy/eS7QJi0WiVfOS5
ZU2EBAeoSKxiPceetquez4QIOwo7cOaxm7+tjLGtdfh9qc61Vj3N7bewHA5CPSZD
bTCQb6EMF4XMd5iX9OHrMdDHPOg9bQ69/sv04Oh921YlYEdhfJ//AdJFvbms9jFv
UAVThtNcSKA8cO/CAAr3FCo4GQNXsi9i7ORQDzN7y78HK3RkYN2QPxZSvHEOMgME
aE20e4MkELU7WdPb2VfZbB74eT3wKmv75RDyHmRXsmzHEFuUMmHpORc2nEUFN8gJ
NbhcPHzEqXWo/6hFMmXCLAE78V3BygFcRiDDaq5Sm0uYQ3t/Jr9ip2QDyD1xhwN6
j5n2aYV85e6iirHL+M59exA1uN05sE/9JQnRuKlqWi+X3MTx2e24RGQQxfZTJIrK
/rdhXpikt3WBIoCt7yw5bW7nVhOvouqO/E+qLbEqa7IVxMtu/wZO4F30VlPzVLxe
Wmd2uPbC3MDt47AjwENoxuu8Qi2oyjK6HaxVT94vIrBduICfclQdbWTp+rGeIlAo
gZQM+Pu9MZINpEnwXzJOkSHjuoEc5O5EzG4QYTXPFuj1O4xWfoYm7UAsx7Nz6unw
Ch09ZFcvaC9A03aPW9cWuzTXnZtRpLR6OtuDDDHXCGHQ2whGWgmc1IAjZvnEBBFJ
r8sLix0ayWeEM0phAb8v/fPl8HHseCy/yJNGjsupitQdKTi36RmeSHF1xyk/BuTE
EIrRNGQX4YS+X7rn7O/L1QecUxZ8ry4huGFOci03+6vC1FtLXnCjm14GZd8lBi6T
fcLA8w+gMoqtVnEoOa45HHJIhDUTNrwTG3XheDNrjRI9UkJq0ofPJjqGb596rshK
r5Ka3znb8mTrvVDdI9Yuh54IODXXlueqMBsJMeAQShmsfmUT8PebRHTk+LVUjqhr
vnm2NPHFiCHXMjHrLgeVAOCgFv3ttXiUSlbG1ctiN3n+pXKxTRSg14LewtP9qedK
YLBB/QAyVj8W7eK0nigx1NBuvCGqLJAu0vgeChrDBXzWKuFlrWhXhA4E2+vNK4TY
vqSGwiaczlcKoIz+UhEfXP/O6RdKxAK9xOLTpWTeHnRqNpYyOAyvN3Bi+m/kVBAk
QpjD7R+UnRfPQuFH+2G/8DPRymRHYE0iC9RpsVeA/6MS2fB/LD+bSjggYq/MchMa
ciYfk9Sto3HC3CwXWaTPy6SKEFwrTl7n3oMH+Aq+ayp2MwVBre2OBXBIIThXRE/X
+I0iZY31dCROMKbDUHF6ILJl2wVP9wKUsPLEnIy4+D0rxZBhMSv/hZopIvREwHbP
wlwUumKZXYzLmR71k81L2g/ptz8vgGpkbsJExHl9fE/cdPFu63rGH/so99vloOQT
bXVnHSGV3Obv709ZB30zwAbjr8ULXSeLoq6etv+l2S0YQmeoyDOPshJgYIOApkmp
TkHBVvDmy78M+I8uH0qXT2iKpr+llC/YxRM9/GWHfrSMy8+bZGmhlIpB1ZOEyE0V
T0l7uU9a4x+j9BmdQBAFerD+QXUVUZheTr+ClEKw6RR1VP2/CGZb9k+oVsKQ6Dvy
+E9W7K+v49qnJMSQn+eG1xIzE2BAJBV9sZRLABMqXCATZbfACncoZXWUfmi6TIWi
8OHD7sf52vDBXzFPCbryB3HakcNVvL41Q9xIM1FhPoylb0HYeAKR2/pr3Ap1C1Jd
whmlzXUoK8M9MWk2xPYiEs7Fiv2AXGE0r1kz6X0CFxIvVHYYxeyYQD3b/vk3h+eg
D6+P6cPwD1ES2FKGolNeOJZh+wD6/ViJXJOy0H3Yjpkv09QS5QdBk71JDGfYhAZo
GXr0mvhj5FroXJ/K1bi2Nqd0gSS9YdlOg7Qz7d/1nYn3COmiVfn6NxZaTOaEgula
VSHF1aVMue1i/QkNTOtblr0Qnf/hq+VOzB5pKkKQsnyX0HH8xTOD+4gLnxvwHPUm
HfzwoXsBtS9tCTn8RknHIjb5NqAy4ibBGAqE2m0Q1E++n5M/X5Ic4KWyKhGnzHeH
vDb8wkA9Oplhhnxm9ZOvEM9+abTy7oewjKc7e1ZWA+75miyseK+yn9DtHvvzjoRa
bQPRmXPUwEPXKkTdj+CXmIqAjk7wPHCwieffgqyA0sx7gsQQjb/gdH9bnzYaidQ+
87jOpookij9ltR954cNZHzQlfDzYj1WTyQm+9liSumfXC5fpRjRJnmcD6j4BM40M
zyUvH/jEE+PauGruh5mZAfSE5XFzxSrfqDSBkgI0i7TGbRv6STKPwVDHg8KnRlUm
vkn4BIFJPsuUKkj0Bj8p03Zq0Rq/8EqcT1SCkcHLPh4KuKM4NuZ7QpqWjvdpAms5
MT/1DYbbhGzjLJTV04JKgS814Zdq+RI7ynfyrOwk9z3SV+xufKwq7BKkPUP78OZF
5bJuTzY3aQDjsCYpA9hnRNQo9qpDRMROQLFlenseISP+g7Busns871fL+9VcccFD
j4fNxXHlF1n7tYGxbNUnqCeEpfv35UXlQcIoqguGM4TIlxZPcjTVQM2PlF2uyv2D
2Po9R59v1Jo0I0gHo3aw0hkugt3iiDad2dA6mvlQOD7ivdUTUsJW93W6G5NDd44V
umrQRNrdi9Oa3j/X+O7CAahoTdZIf2l+sgVjSCYBRp29v2NcbpMZw6mN9yMIz9aD
d3S1h0q8Cw1meb+6PtH7SpzOGwpCmMjLh6P6cDsU593nJGN++NykvtzQnt2hmr1o
CbVEIostVjtbI3VSuc6Elqry8ZLU+0fVoq57Of/J6y59sWIWZnDYtjgQ/Y6+ljWx
hvs19sO4iBpfdP5kQP9pY0ykUZSqo7PYsZU8vz5Sn2ncNrx81bpa8/+muFY+4sRH
4YFWIk+eETZyC2Rk/Rw5pbptNsNo7NCw7nxXjnngjSoaeWNiHJxHqUeJEpPQedOd
guUcKWjqstw02OpX6x0qhBJaMSOvnJBV+y9avCDRL88Gy9eQXY0RUxbfECboL5uK
JnELyEwSA/SWuuXAu/H0MXm+hrks9luH/3z+Z/o9mMae4u7NPyLAmFlJqrHAphTu
l5KD7kZZ5nWDzXrNwVmV8dF4oJzS8y7ILqBIx8GWHQb2fm8PCQRdl467oOSIbSZQ
NEdHKk7NxGsEi6epR+Fqri62f/wIX9ZH7nk1gpCWATvW+x4tDzpa8yIhDSF8i+bZ
KwYxFzvPFnmeu0Sm1FgEG3nClZH+3u4TInWEhytR0lo+YIyL3gwD53KGvjulFpQN
wu30duX7RgmkX4KeFgKjmvlwCy7LE95did+nUm5/JGB4kFuz2Phj8NFibI0R2Ndf
Kwa+Hkf1vVQ1lQjJ0gOtwj+lB+RiszuXUgEgCKdhvtUqPmWbIbe5cUFVAX2nMnTQ
HrlRnauDUI1NaoJjjf5VF7LZPyIRW33L58EKJq3kJnVAx9TA0HlE2gYkFonG5Fe8
z6LwBnWFMMm+1rUaMPAry0ZvUngr2AYmi1SJkpeyRtcHF51AhWIxKmvvperA8Zb8
4MiCpk2/YJAOhBRP6vZjFickWUOQsFNSScrdF6VSdiFQQuQ/MmDj0l5igX6ZSd0Y
jH7DDynqd5j4YoFRnIKUcpbx80lRjrVe3vFyOjsGknqEtdr84rNh9JJub8yU+wVr
jxsjJxSes2GrkME1ZeGx63QofkGtxLN4NvDISXJYQsa+oNcmGmlL1BirjASONqD7
Bb5XybmcpmptnoGFSA8A5MvHvJYcFSfs5iH3KFmnIfXzByERo3SwH1FiWWQahzNY
nGTDufz8k6eoo/szfC7NuOIRhFzXrkF4EM8ZjSQDKqTT/KfiP+6GnLQqy1Wrxh1g
oMZWUKnz8xEOZu4YRzMWZv/kJqL3zNJkdnVQMvdcYXKBeOTlzdB+S5uDIaEnnv38
9zaZoKD0NdLuqc/uqowLgJqNu7UFZxM7IAeeV66Snd/A0kz1PXdCPeEI+X9f6bJk
Xy0cm/wSl8nzpyKDrDQmpO8yMU5GWsgbWtNhJ5Aff5fr0+mQQeeSEvvhP3LHJzir
DE+FvWgbcxjpdT6gL33a9xLQ7gzGdRJ1/ra5DegWUqH/r6O8jty6pfKXaXARS8IU
TQJuzA59Wlukll6BY0niT2MkpclcCOO9eY5rQ9t26oBopeVKsp/+v3Xw7CyN3H1k
waGbGvYk972lf3YSq8j0CBYs5oT2yGGrcig58iGZhKXLkXeVdsGfY6Bnfck/H9B2
n19VYrDjO4vIAQhnPnO2T5lM76m0vzmVrsFv6j1u8oVhDkgLxckROcf8aTIuu3eV
BG/iuUE0vYoPVhw+v6gtpFV3rUih9mV/YNzYIbyvc1n4vnLaI0OaNvRe0PVbCTN4
gwQYWm1xnE9iuaj3CWU6ccNXQuNnQqgIIyIBLy18FiCdjs3zOhxf0JPW0e7BO6q6
GNcMU9GCEFHL74/oCfYcuGRUfsVE31hGZc/JL2BhBB7wQiiEGyqn2s0rIxSCQ1Bp
fXxvJXJ/Kyq0ezhbFH+za0E3QT1aopAVDynxTkaTtHrdHGc8gO8zNKmFQd4723KK
oOcti3wojNk2vDfZeOTX058fxDy2StXcmlEeEC6PbTPdxyKGtIhKOOC6zvugp08G
f/pA9e7Ga7Kpln8LSBm0QWNXBgtVdewpPufu0hJlqFXIndiAOvWJvatRuDbciCZ3
PPZd9ekUusxdfy267lto3ZWcK9F4XSx42EW7YpQIk4eTRWJEXaUWHoMS3Z5r0Bmp
ZVNXUkieR5CMOHGfLaoRD42Ym7U+8FBqr79I/G97d1aAoYQSVu8oyuEkW8UVf5oo
4JU49fNbDQvXBaJmqiVOMEN6I70v3ZzGm1hyOTlefRzQffpqssZgh6Eh6nKWrtOl
HLOXImyVzb2dp6XksxrX80kA5UQZF3BNu5PWnBdyFhfmGBVyCvTDPl7KG+zbzZ2p
6p/5fW21OTFK/OWm5Ms/alb+pGt3wyy9muFULfYDaLXuCrIu7/PNOY5XoNa1nSEd
No6dCizm8qMMFypRbEVmWHOLktd5f7edo4qU2ZZyhE8LaUPATmcaiztH5ac/H80z
Eb9wdvKrJihIExs3E4AND4PmQkDpbOhFBaX6ZF3WoNf+DbMByhX71esTwZWNREL6
9wjFqGl/ZXeSJjJ72e5JeTwV9F4bSoanVuTFP1xTTebCRBxGMMkPZ/IE+eFUDcT6
Ca4ZQkAHJfWnJtJNH5Dy3zQG5PBeLwRkhB0nOn99K7vS3R6d2l43fS2MLETvWqo+
ON7hOOPYItOfwLa32KUHBxivu06v5YfwHt7a0Kp8bCgvwWwKHi8OqIjyNEq2Hvy9
SoYrfitKp4h+dDpSUMsOWfINg0kWaP+7R/KdkBgJjXDXBRbRr5qD0QDj5f4TEJNA
I7JkCa3mbhb5l2POppYzPA25evIDrnLrb8+V7Ea0tNAxQTeEbg5broDGJI9jGfQy
rQF8PdOpdLzCXl5jRv7RR9BHvPkEYvwACabSJdvKOmukt3S4TFE3854lztStbhAf
r1e/1k0EtM8eacG58kgeL6UC3eaQ0fGDOXfO1+2qg+yehkZiEoVA3SCDiwA84Pzf
S2mg30hI25cj7/WFgQZytlPnGxnxNIVvuHS2YxEoHR6T27fPNY/12r74SibeVaNU
1cAlctLtA09DuCYKBkdwRSAxhSngNy5HIwaLi13EsyLAg3hnlkjShq2ct2YxLL7/
S0MreXRrdH48Pf+ACh4XpbDi+W2jBznDAN6a2ZBN5Qsz8JcBQ1HHZ45sEmDdvWar
cslBxd3ZI8yTDCH942KxM91OaevM8en4RktRap1NsIaUc/rF/JU5upZDAcBw1gJV
bvaZZStBKc43gPVOdz8iyU5LNdo0Fe/p728Lz7luQiWuot0D9H3Z99XoBshmSfZV
sBM7d3wkw3f/IX7VB2K7iBlU670jK7X/kslzbRwqbspmr4kFBJXVVgqI2fceUdS3
UYSaErUIbZZyjFxRX7RZ3dVQDet4h4JPbo0UDxbOh3DEckSB6LM4NeC5syNZ3zB4
tzTFkzqC6zLN40eS0VV6Qq5PB6C8jIWM952THgkV8lxKK4689D0rO9OVhOGnxoFh
X1TDBtRIy0vxVtxp3GOtVQJnAaKxspx7PeJ97LQVRXb1KZXmqLwrpfGlsQGKI+oB
1gZ9GlWuTh2pmd7GLAfFg0LgsKsKCFmgu7vH0i9I+WPaUWvP5fxm5Qi9UrKe34E/
KsU4XwwxCs0NujdK1W9kp3FF9lbox0mbioT2ZqoWPvoJT9h5UM2ALNoA3rTbhdIy
/ry3u61hcK/FQLoxX4qN60Ov3P24Qdx+DZJpEY5fwE9kNG3sD7gfxePNdoQ4wfFt
FIbnS5G1bLnBTF9D+LNInZaWqx8e3Fh9qGTPi7rUEzyNc5fP8Rl5EXsev/KuiSTX
qxa22I5kEI7q6FkBm38jUGbzgYVg/n9DfgRVFRnCSb0NWLSECz1bmCtbRV3GnTVo
3QFm8/BurvrM4bdCXsrYHxvrbZ4iHw22iX/eXV21Yx3EYMuoc0PQnGQn1hoUADxy
zilEOB/ml30GkZoRjvNOXo0vDzaYf69MNm8m0TI7E8ONR0HiTVCNWF/krf7+JZ9H
FWZba/A4YEGGEKjCaqZXP/L3V1TuHtnTijZTE09G8IflDlloIgh9rYRxLhV7oltb
oWTnQZcnlBFEqWCZDZdYdQ4IEyhsarchIsWJB2voblEEk+E/Qd7wNxdiEOcChiHK
XtwIFz2X0xifSO5R/RY0QcaxWxqOdpR2jZCtX1ydveoeJjk7SRprz70uUxdQoJtw
qa/nWybXqcGMr8Z/t8pdom65Hh5CSCT7yV2N431RuuOWifPKNLl0pyB7cbH3wDQV
YmOG5QF/z4LqmYAuxIwNd0g4q3oFvknG2qCCp3EfVCYd11MMXCtnbosaN4f4J8Od
/v3lRQSWf7h1BEetW3YBHC0E+aujXXOR2CO1AQfS2KgbaEwUI/Gxlw0Tq/3e7dcB
8t0gctvEhvtXb6tFc3mt9U8FOWTHBgCEusAXOrKgw507aI4Sghi1iip5Faa5CXMR
hnHgwSg1vfzqP+sph2Cvv6WZwzDqI6nwat2oysWXTDNFL39413qpcFg2eVjw+bp2
glNTedFvU3YlkhK2+F4ZS47TT0HZUJmdwbNTpqgY2349+lO9xl1p8rBJL2ouSW0Y
YfVgDA54XtExkC4FysdH5Ku67S/T2DqdPoHCfKgfYDN+pfqBgybO4nXuvHKY6cnz
NUukV8lmoa8t0u/QC5m6gcRHP1qVbkxMKdf+S4jpmbTUBOeYYvoK76lOmhwguHGD
vqLy4c92lB1dP5+bJ4EZ7DOCCpZbGH7H2dwLPPR50DGuADOXEbgoCmj/VZE9f5ni
XG74GfkY5v4RsrWCtvfJ3hDX1TSFauZXZHAjmpxJz2AIcfHgsi7JzQgQNyzEgqov
qT9FHShoEhvgE/VDvTqQ+AWX0NE3Dlon/AxePiTroW1NMjy3wNhB/8EXg/1NBhdA
s3Ar4YEYM/wWzY5fOmfnfPhz7qJK0zpuKOKOm7NGKXXZqTo0p6uUzD6U7lFros4V
6RqTFz7l8FAzaL4tkwVYJB5yDjkaDia56lh58C6LqHjmxsvH5G3PeOUEzDK7eyg9
w2GsOCz9lqjyAE7bT7BEMm+oyt1mqdVmcRsLu9xMj9EMktT0yBzYv+UVn5gwUJVn
YTn6Wliw51sSKHzNndq2iTq0xyhqu/kQBNcnmI7IZcefYR3epFqhsQt+UW2bs0+y
NKI4adnR2q0uV/hVhOGptS4hllhQ6IY/bwuHMwfkhc5P82JtPkF1MN0I308Rdx1x
hGvoIF7IDsjzwZf9JT6/JbmffomsDy9g1jsGpGQlhRdhBw7yklESJUnPDxAkVHy/
oS6mRMZM5v97cRDFerJcJqEfTaM2z8izen3Sv89LCbnMZOEw/IWSKTiI5q/emiQt
avZ1XI2wS5DKc2F/AAkVLVSjCH2c7PAjD4oDwwno+9G84j2ccJjxClW2zynbVRX0
Tk3QQpDhJdIBCaAepWiWie5fPiaa8CdtLlk/0CC2DyS6rLQOwC5lUSkwUgzDRlr9
5SmmsIssNYvFvpGlCaGJe9PCGgzApb1HVQoA8qYUE6Tf8VSMdTtkyZELtDPBTIsx
kBYETkAmHtUBaYATUbRc7A1W9LzR5pR/WMVXRxQOHDijuYX+xc6VJMxGmfeJnHBB
/YtRaoQkYpFahfgsM2l2txIzU0+yULf1g3F/DLjHd198DP6ENRphyXrigoSx337z
WwylUvzZOcCKHFCxO3/YSkBNgh8ZIS7bVTFvZdxXkBvlIJKOt4jd8+nPf48jTHOz
UbWzY+ZB/BJR07aQmMVhli1VN0ZvRQq5jebriRFodBInLMvfEK5BJ9/ru4NoQgER
JVvndt0MqkK9kAF3NeRMZrJBzDfCtExytslwW6QP07Jdkgr/J7KrRF44IonDc0tx
A+Di/wVcMH9bIVwdN7j2MSLowNAPBVW774su0fUD36QTviHslxmX/pJYFOjjJd5D
HWjVum/P3ewUjAD6hTYsqPZ6dI3NcrV6l/N+S1gOBMiYI5HX+laFrVtHVg+CoTt3
uglVuhEzPyJVmckyqENnF95vu7/KwPsHzy0wfpagSa0WGbHZs4h+W/iYWu7reFZi
WrMupGKDdxDW6wLACxnib+aYsiXH/uosjX59PRalIrZfl6te28PvaoBrDQgfe1KY
x/OkX6CNiE1lYGKzEjkSVqfwGAMSgZnsiJD3rwWVA6XKpy0yULZvOUkiKEhRZ9Sk
/T2FAZ+WksbBHcJ/NhhNtyu0777tMlsxk2yEO+YQtXf70QtbVKSC2e+wNdrk90CV
WWeLNXRF25/x4RGCL+/+WZffjamt7hQHpUxFbnh32L81gu2Rg+SYBOfFsgZRUJ5K
fXgf19/P4XBM8rF2L6esX7JfR+rn5hvlF4fs24ogS6q3k7fId7P631mizdQZpg6Q
F/u1/Y3vssIPxugJ+OKFrZhLMThPgtV/3uSW5WGt2ogdTA5C5jCKHfjpg8vl9Pct
zzmPVmSJPqLeBgg9QpLWuYvulW6noG7LiNO4RNECYaG8NLluzjlA340wKXhohZf2
XSTvuMxzXoa+6RGrxr+DeP0AwHs3lyHZXuZjbD1mDMcnKt1+98x5OEogDtOxdfoq
CWbdJYBksDk32sbIOdrN3FCQ3qTcNKgvxkCujpmObUUWyXvdrZ6zaVoCR1ROPewC
irOKyJq1b3Mv1YVixNDceySGObHmX4dtdCqjwCUg2vVLuoWSGusLT4nLTce9+fnl
1JiXRfFEvY3z5ykm3orXIEEGDFBJnSVFgbx09w58hJc2Bjm5nQyI02fyl4NKOMzE
jn9d6G46GYhbj6agv18T5Iw0s3N98gBAbGe1ydfmy4G0+SYWAmNczjL/AkottBPf
Z19qqQKSO5bwddF2w3rRJJSqyQ7xg7UWWrJHfTjURNgjZ28GlMMxA0krp6PG0ASk
YPOlON1rRGTrxa0xODIvMA/NtNJMaR4c4wquDl5yqXZWwCjcME4kmT+5cGkRuYCI
KiGngS7G3P4u0HROLHryhJ0eNkEtk08HQF8afLMuTA8pd2PFZdgZC9P0rWKvUIXY
x9Z+a7uM3jD9cshTqROdIbDP6GbnTRcnn3sxEvP64Q47gHEf1WAqvW/51cveaXYi
xkCNFvYTezkq4qMxNOUXVVt2jl8vrAgT4qbpI07dhDA9zGTK/hBMp+RU37DuyoKa
z0gK7BL6UAkbtSERyIa0GvcXeGVeyuRhuxvgY0PORC0Xsnq3aOzjLxWJn6gj4Del
7iCG4GCrPoY3P+60HY+91Fyeb1ynA+8szbGUE6Qsg1kavcChtaaX3bqUjbu0u/Yy
OuLx2OA9Q+Zcy9yk37Q3zObPaeJjGCnaTYRNL2aTiWh8m7ufJVYSmtl0AwXZBzcM
pocnUie6FSoVa1Fq+zOeFYdm0XYopJY/r/kE0hRk0CfPYvc0a+KCgV2jElTOPwa4
tcTswdwjLikSosGzAIxHdajUAEa1XsiNvj25syV9jWbdqe5Oqj7//QVU8+wj0+PL
yZeGDP9hj4e4NhuKXC1bR64Nez3CzhUoX6ANbumherkRIxZqfHAdAVbyCjgSd7oy
g8MulOP5kOWqv8uhdgTVi3to3wQNw+Z2nXg+PHYUbqgOa1vY4BxrNU+YcsGDrzxD
9FvKXoPvt2w30+ZmBL8Ixdq0S7K9EpcVDO7u8yC2vQ/2jtsF32CU/HgWIBzftBN1
pmcu0zPvo3IaUhlosRrmgo291CMSsMq7G0O4ML4LxOtgrfsugMKjVLBSR9QRDUIy
lfhmpT9HP6+MCWMXM8WJW/1GBF7nHSjg+r56t9xPINzaxHwp7HNRptkabyBJk6Dg
3U0FFqqSw73xYUib4t+lwkWOSAMxZr2Zh3+4mSMn/uVWAkT+wP9V8ZB+/Aq1d8Ky
d3KGWuA0yqiGHmEJf6nU9Qsj9jL9GPHDPAoZRbt9DSXncrxGAZspdkhMEkwsMl+l
+GjcaCav0YQDDAxlSjQfSgazj0rl6I48Ia04abOIwUn9An6OP0tuSAv6Gsr22hZM
RVcDz/ETj7J4POjO7rdv/bX+1ngyIE8xXCCO45LPCPN3YzrKo4xj8BjnRKdDzMup
KhX2swOTYRpL5F5IPahx6GHZtqjUS/BkdSO9Guc3OXRlVjj9KjoK+2xJRGOXW9UX
i93FrXPC2d4d4PIRWKCQqWEtSv0ODxNLtJcBsaZY8ObWTQ4FMlIYZm1KBWIQ5q1O
4HkfJ/AvBC5smqcFyHQ8GYsQm0aHqxawRrR244gdinr2I61mhLq/dGuN4GDY61Me
EvaeBZq016Uw0FP/54QU4Izp94daDv1CNDIUS7uGasZzpE2ldB1uqnjK3G7a1/OK
U9UzjTzPEPWe3xFvIWtmApEJ2o5QNBf+pcPqPIKjA8JWzE08nAQJBZY2oz6wMDQr
J4LtSJ6P8PPy3UNWNczqASNrgV96P+vltY50nFxEBG/oVm9f8YfWTnstEh78Ohgq
rrX4VGCW0smf+JSIhhB6N1BhLOalxGJPRrBPpXvMPGb3AsXmiRruAxECPQZkBJGY
XepNk3G1foK8NBAE43jINOmHEWqZ/Kdnn/xaeAWimtadoml1WE1Evcm9uOWKV2R8
go9DJdTRtzCRB7C75t6WiZSG313DFeif7ofS2PE6Jx6cbqGLSdSvEVFb3hOJdvGH
z26+KJR2t2WqjPIlS/g4mgaIhk79ExbSp+8L8KRIRYAGPk2k6vjrGitAvW5Wf11i
KRySpKuVVktxUV+OLSu9FfjgS4AGTdRrOxz14+Ku0G/uNcClZ3C8FdW5KfxYNEtv
baBUPUUpSvEfqRGreZbWGKBaSpQo+Tyly+bE+rdeNSQXUDme0V8GxqfN3LI39Kj+
63wrGXqnLdm/mBCoTEbuCMQ2GSI5nxPQu8LYbWqPzsvnsxwUNkv8vMGvfXDxLBIp
nUjtkIEVK+RrdrqQj662wNfjH0QiF7WB216HQxxjWAqJGVAhNdWoQfadUNjiLCWO
REkkkqxw2ovg1HZmauZve0twbk8WfC3lQKK+VGPpCuOOlgBIsUxwKJPEEATXmUo2
uNPcfsSP0VBzv1CDH35SrTuBlQXrON9zeN3ITQmiv4Ah3OnhDB0Nige/UzrSp/eq
4z0mnCEJdajoPvhOrteS/bWSqv4hSy/iv1QkBtTw3rVKSLDkxomaZ39FlKct5Yk1
J3Ddqjt2AmbK7t0xS/2v3D1Qpc3WancWgjG/M3DJb2wEzmYGNq+zVedk4geaO0kx
7nUw+dOZ6kZZf7ZcpsQf4qDAyuDq/CVhB98Xvf8OIdU0szpJ6e/5ohL4mfOx0LVZ
K1bzmktFtAVxtY9J4VWSiZ/Lw1XSkBMwFs6etEyIzJvYd+rij+Zam+tO4CvOJ/fn
9XNgqHg1q5R1K+JadshlFMXynaTb2SVrjcGZNKg+dtehgjU2x9eYRjZEI+0sVqfL
0BvS74JAMRZ0YsoCY6j1qE+fdKppsmSxHwNTFh8SbGeTPloyJn9H3Eq1tem8tAxm
tnBndw7J5zbj/bLFz9A5LglexXEIHKHoN2r/XTBrx1MJyIGf/UWt9ZkB6zwyAIkn
65ARlcegJC1QrvTiTeAHHXTzreZY9lYDdwzerSsHgnRFbPX7LGi0UqS5s8U85Otl
nUkTR6Nt8mW4fy39enerB+nFJlxtlSZZsxqoxiKuwVcD5C9e7sTcTEYTNQPD2JTL
W8li5kSf0RcgwW99GHrEPq5R03lZ9Gxv7eU3Sp6vCM6nwP93J9hlZaMv55Swd8WA
uwuvmkcVF17VS1oGBBZPE2v0mviT+/t+y1/vLlJPUrR1guQ2mULx6eMI2Y4Y3eZ4
c4eK9g2IzBtm0WRCbT9cXoWq5sghnokOU5o9IOu+vBsQX/SKuPL+kbyg5janW7+A
/SRbJx36hIUWz6qFz4PNBZW68q8JRwZfeCfHJYbR2nOb6LOQmw9s+TtAMvGGcnp0
e1p4qLXJaRTM8P7kme9u1t0jeYF5JBTrUba8olIMH3LMCmyKheFcdkABeAr+WeFV
dX4bM5iHw8Q85L/h5FdW58tbWaToHF889W8oLFGa1tc2ru2Ict3kjTDSX+vCJkNO
EcT4bTlnRz/oi7BowIfuzVvdqIgr7KjG6cN+Xh8WEj8IRBuqGL1Hj6A7p0qgUnzh
gbfsqCgR5NqnfNqxqg0fzZzlCU0WOjTJ8jELZW+z+GVyl0qkgzX5vkvrhbHBwY0v
oFFQYCXl2HJYgsOy8+yX4wyUgy/r4RGtCERCnflufIHpaNb0GAnUNSV6SOdxee5/
IYZGyKSVYyLqemn0LJ/s5Di1tkB3K2PDh6UAW6qJdHkr6OMNbmuL/DC6IGVltjW2
kreU5uQZ022Go/AbF1gwPfU+e0kLn2CNxO4NKyXvC5KZQBuPvEZ6H5K0hRpDZOf8
ojHlMrNx4bh/lTGgRhTZHzso3uYkPtE+icmmYaREr9X0JLsZwIN+UKcLHpFcmQxq
PFh0uwYsJjWUjqRomxjEEs//r7jkr5ion0iIcfTzyAbhpc3Hu5DbNQoDdrZWOIFy
/GW6WuyxIrcEQU/M1qaYUX7t0zAs4tOm6yDAIMD+YgTjRI1uhCOsCCQCN8lMxcZY
bGGxHn8vqPWIW1362UlqqDiG5Mxi/H9E9moHjrdNqRKgG8Xp5r457irrR/b0+EbD
+wvUvKCoDmI4iOJyjyqYJNRaDPIppuUqhOeXVl2elgDMrYrC36IpkyX8ij0mAJ7/
EDuoQkBh9180uVkM1QURPzq4k+oKNXPJfk+8neh3BkVVM2mqREDteFlvNZPrL4BZ
2s53q0CvT2bjr+c9UZDcR/B+cfQQLvYpVoBgGIyq81YZI6hvT5Bn9OOebQc4TM9U
1TpHqMcZN0yKw4WoOFM/P3UtjXwF7Bezqaj60gT9Yu9M7xHqqzfjzYEIdK6adszk
nOJAgWJBJXCGXw9jYbsC1ur/84vqDxdB+wsChMCD9Ssv24TBFCH0Ki7+nh3VpSIW
DxC2Ts0y5dDGUWzBDmCNyIek4HUX4Oa/lzvYtJFrMPtlllduhSXuDYJQXJ7xVccH
C6lV/Klkea3BBd85WskNQ0CgnwoHJQxxGweIZAexbHKu/PxdF6X1+U5FyhAczrBd
z2HWjU7cGJogOyP1gE+t5eOirbEpaMB+SZDYByAFRrXiOLOud6UZhs+qxnv/bcrY
i60P1krHvgb9dABPWX+LZ80LjeE8JC5pKI1g8gPOcxGecPYKvE5nzdppCNGB6Rq9
xNiU/zmk1cWNF2w6PHrgZZB/pwqPXv4ev4b5N2NHo9xR8eZFXQRwfM8GUzGmQUW9
i1HVMAWKBE3qs/GBuyIhM4zhIox0pTYbtvAJN1hExl9FDsAFuNGLpy6beI4xgtfZ
0xLrnvIlkctS0DLH7QK3vb9XfcU9y27lpsKjC5la39PznX0O2INF0oQ9hoiPZIYG
pryKCrWlAjLA1NoEXWIlBhG4gNnsRUYdI/Rfob4FDTyiElhGG2Iha4BWnDZeO1+t
4C0Z1EFkn6QCarUezg4eWyK9I83iFnLvN5L1LmOJhRaCtX6a+8SAZL4UK93HbLGP
QkDfDOoe/2Y5MdUrshEvOlkf8JqB7UPLHGZfCiDycHkTlWGMobEaRPcNHxmmQxsa
b2YFwT8/+M7RG7r+1/3/p41ChRyp5qE+Jk/y1qDvMcMC8FQuKM/xoBOzvhFmdDwc
9qG0/VZvwUbhlvWZaE7axpVo8sCFeT2UMXpd6yLoSK5o4aoOwUYGcZLLtaYIpBoy
qsX+PqHKDAVZKPr2+ze9CwJitUGq4sfS34P7Aqf+VGZmdCRBw4ObhlEM667tDboI
EpNuQgvxzewVBG6PSxl5KjE4ev/zQUEBaM9VDII6gMQvA9WCf1NbEgJcSCY1rWWW
aJnKbu/ZLpQshyxTayZI9tWBFBwXKgc0Iu6WP2vF/rIJBm2nCS7UgwfFVdmyEq14
4oesy7RrWCmKm5tQaw/k75DDSmYOAsA0HK84T4q8Gs7bWttnzClfkIQVR8y0PB2K
yRX5lvgPWe24pm4Gn4JK95/5rkVbOxEiSSaaQSmQInjIa9M3ymXtFyYBTmusVvEc
fmjOMhrmplrOA7MOz+hxQrNTW89zpDpQbBO00o6XIsikSS2Ua2NUXqHMulE136Mz
a8VkzJF/f33eP/R1h3/NpT8U92EMv1RbSbQgKLIUC9SlsHTaXsvhrGGngwYugbaJ
7xGq7tcwVAn6WBfroOPVN0/RnAqQPM0du89KhK7e5dRmGdASnaRb9aCffLcto8zh
gANo8G4rQ6tlaDc0Z7DtOQCemIn2WHc2y1DruFPAZZz/p5q4KCuBe4VLwJTXRzN8
3VGaUcWP3BJl3bup7KTlU9di8V/5/Oe6GmgScGxXNg1xV2OS3xzjENIVcyQHpxCm
kU79wwn2hf8xd6Rf8eMIZ6IgVXibpHssuvSoWEKj0JpZJWUehE88N4eXMtzR2a/R
xPOIh5M7+k7LQFo13xVLj9uZm4Yh94RqOMQSh67Mv2nG6ZJS+gXyQnBWFu7b5HYN
/ZEbjZR4zcTn9TTgH/Wu4Ba91Jxvg6J8vcJf/kLnfrVZNHm8XoYUoqthGjn5ToYN
nj0COlFgOm8ybWbvMTjVjoumMDii3U6kDxt6bk79j6ut5Yu6lNtadznhVLxEXiIE
FutnpDexgDvLaX+FH6NOreWn5lbMb4lxL+3nOc6a141sNHB/DNQPCaldz3aQ0uov
vuIN6Ni9rM6GFoctZhzK3ESDwBjx9Xx/FfBpiw5aEfOndkwCCeu4XI+58W6xwGRf
5jZ6pMZkxlMVW7942Pprr3XWy2orGMXOg7ZPemQhRQ5YL6p5XESWyifGATlrCxvt
Xlb7CL+7LMII+/hmOTaWIsNRI053bnA8AEOXfAizLblINopzN4NQFhlpNXWfAi7e
N6C6sV8MyxmyF82Wv1ewyn37ttpyEur+8HTZ2DooZ2Ayirf5wpZH4qvmWTzmfBpy
JwFffWNLduCbINCCYBBUVreaio+NVahJRsN4gBCvCHaIaagRPQKp2Z+0nLULu/XQ
QdZeM3shf/UuIX2HIY1HMglWCIuz71VpTbY8vt18ok/m/nRwpR6rQU+X6RSTjiga
ezNlRLgdurs3JxHHd+8HZwKE33MjQIZSk/pCz2TULTtm03dDYJLqjmq9pRyft1to
Lxtgi6CHCziEVzo8ksIJvxM9/zmGQXm1MikQZiKq93Ws59BHZI1HkSR78JVwceD4
ANDOyak/FtiN0CiPWbNTQO9rockTNDcWt1O+TL1EmNJMs7aUff5imJl4sUbhXQaA
wpqLGgvO12OsPS0dVrYds2fwX6TG1XMwHlTupdYGSmz402vdgHspcyg7lZOdxE6d
7LEq4zA1a3l97ES4i9zQHFjl8abDrDmkq/QXP513WTOR6OWJsDUai5vdlk/m4nY3
f/GtWgdSphDCQqJNAzYY/T+2JuJ5s+GlS/6uDfO03ejgaPYsw6uX8OjbjFWhGnv+
q8zFAiv/H9FUSHRkoUHMlx1Q4OfTWMwGWoSE4D/FAcrBEa8Trj96K7Wb3jjkwVy0
dFU92fCDwu3CG473JGghUKZAot5vexvlv6RC0LX0sXmu8ovsvgkq009Tzq+XVxDk
0QopPxYshbh0ueHmPdfPhIjiUGBIvnRHW8Itqx56pGMq171IALlT5zxLgHHjkrer
i7Ny53XXVQbdDBkIKdiy4rnbtYN4O4gnE9wgXRXNB554nQzMtshJHwVicIDkOmYI
0LS4nDr4gFocd4acu8NXMTIlqnV+4kWTz1rLbFBMN3o7Z9pzTfVq9l1i8JbDO8sM
wOSIfvroc1k3rEJxrcYxFUPAafb8TEX05mROF2MZFUhfS3fUO3V7/lBtysnQqjQj
+4qpZmhPkMy269rjtHgEJIpoQfrP2gffSoJbvWtqp0U4npCK12NPgz2VH3lWAlK6
nBqzwjkECSjgT7c0fosKHMbMjx42zyP84/vfgNUQN9W0co7GB+BjYlpkxa8/36bE
VMg5Kx7xwfgNqIHfYtoBhhJdqTdvtNIE8Y3Tg/JFwq377NI6lpvGFizOui0rQpug
WK+oZEkNmb1FHBVcFTOhN11NfDK+XsnNOu/ynsYevBX8SXWaOItI3fntd2SG/yXI
70z1Rq5ORK4U8S++qTWb6c+5hkWIGIssJMFaDOTBtHerIO+kLzd6mhiCeaTG5gHd
T02PqX0+lbF2uxF0NqahmkJLxvMHhHFqJS34nR+iD1+yfz+bm42Z4gxPnxiHB5tv
Yb4Adp2KRg8kPYIqnzjUXL2pqna3n78ooUpi49y5cY6pQhBYDOABifIUXLFuYjf5
S1OBHgm7FbJHm4pKCcSolUSuQ81XeLICnUYWzr2UL/aZSmZ4WD5J1DJ7Q5gMKEML
rXcoeUgxF5MpXw0JrjpieJEivbblakxsauoaBIp9oWfg1fUOZGtCFrRgkGme2WhT
avoKQc/vrTN4hsIiYGhEH7gZ9WinTlTdQTSnn0Km2oS5MNef5E4v7ofeshg/jKQg
2KCqojba6tqO0cBUBiz/BAOIN7S/KdyfC92pj/gc7uN6ZmiaaNyfSkfkPUpG5iDU
e70nhuyJbnYh/AV9nqKznX39qK9nWlYD6Vaw0MX0DKIVOoc0BVNsQiu8mRJxiuDp
mqApXq3rPNJjv2hF42yysf9ZSe1f35M3Mm2h1RmJzJGef57dH6tWQ9k+8geQhndF
0NhUxwftlEpYXY/ubJj6AuUZFmYHURxQma3H2spkkXilcWYrLpynwL8yQuYbJf2w
+rEGlW15dblxlCv5PV4rB9ZjxFUwRyRsYOWQk5aNUzYSJSy+i2mFuwmz8CeVaFB/
l9b2ascP0R4Vba+ZG9TyIsZaj3rzrCtS0W47oTL0rSqwah3wrZ1EyjiaLMprDFbN
fSzgVFSmyEHCTS3XPqLuZJZ09jAmhfABdp9ftPKISqewmN4OIrBI6kYcJkV265kw
zxOmdyklAh6rJTGtDImk72ochd5tUdPzftiLBxSCp3hjPZ+tmoFWdtOv40Gv1BUd
GYPTLs8TgMIidj9qehSHprqboleLPudehPrBuicnKQMiAvt/SDvajQGnKA63bJBr
1rOSsDt+Khv8954XX/oMZsnqoIrZeQYWHbcj71/S5Vpffm8a+lZDxxvumnpcbrFB
8CkMu9VmbvC6il8lmHSHbN2QOxtKKb564O5aoxyBCFgcxD/pu7ikpgO9UM5FX7eH
/KHAcPrPVAX+SVAY0oikSjV6jPPEi28tdYseLjf6bXHoMX5+an9mAzUUrO/4jsye
a8ypQ0miQc4CbPG8M4pBsvMhDxipPDtKCYJ2dXfDeP9y6tYMeAPZ3UDroWZsukJX
pI738x/UCfH5EBqt2NQ4+N+3lMKsEM4t6eZseoPz5rSdgHRbmguRVdF6MpEsK0XE
2XsKHWog6nCm0e0pWRfOrJ+vHVDwDz386Z9gPlWa8A2ABGRfbi6ir2v0xq/8JAWL
u6Lqyqmi7leq636vR0lOyPveoa2ty/3H3GCnb3j5+JWJ7+CUxb4LVnWF6tDqEI+x
tUtsIdy4PWEda40/6KWzXjsOjMLk8LsBgkVFXKAt9wOv/CIPDsha+WS2Z0AXzXCC
HCvQPtoGj8HH1IbNfuO/9fOb5qraXeiGdSx7uuRClyuwhDmNzZ9LperxzYJHQ6Ze
jUyifRv3qkaK7Gyb8qM66RyPqbiyG8to6ul9WT7dzAJNf7DAkP/f+fIDjecJ94Ix
eQgfp3p8lN9b2Vq2eufyKAX+nnUITRYoCf7Z3rh/zVi1Yu/VSPv8MwypyI3qnJGF
LywUYFijeAhIERnV2P3sVOu9T7GsiOc37vRM3qBACpn2yw0Dqpd8NdtgWgNtgK7S
YbfW+KpiELb3Zl4R+CG0oR0TsjJC5fqN/uHy+ykttnVvUgbBkY/R/1PEKCY455UZ
+JRHemGMdt8KVF4fLxCQjh6mNy+iFst0WoYSVeplBL4THFfGK/nHHWbiNsBRM0PR
dKaQe+NG79UKINapjJP/iEFVzyqxquoGWklc8M9QPlpXmI1TBIsWh6t/cJb/33PX
3g7ZeH4HmTficf3mmpX17QverLYKnr1phw/9VIuj/Om3T6WmgBRUVwMG1pjfdC/V
zlhKok6V7hQS0t2wwD+hVUeF3CsnFJAppScS7vwuf5twy9cmtPOVLbR3rpf1O71h
ni6VjYkI74+PH1ciSjrQjHNA0Wxk6YRP+/vqpedZ97u8VHtXRbf2JFj6AAwKSzj1
6WIR3EIxycSZ9Asi5pN7BTVl0IN4chSJ3oxtKM25p56B8mG6TWtHl2nBA2rs0jR1
0+BdaAQc+e96tG2+lYDvw+YryIL++AoL1rifzfOTfubGZP2R4rP9/TW3doyBoUp5
tzKzD+AjZOiUjAlEQrNfGeGlb7wYetg9g/LP5xmB1vI5tQBrXuLZrAbpA33w5Xlc
t20YAJ3GHX0rucMFPFNFVLuaPOmJRa+ZAP5MGymubXKi5dTtrVzgtf3lnBBsdFHr
rElYwecAaZjbs6UTjmRGuM2JJDh8v70xVGXQlpxSamsTWkP4le1KTB2lBgc4vZOz
As3vvWt4NYQe7Qa+ByraRAjqJk4B59bEerNDjTEXOXlP60GCPSZcx+x5J5szNuJw
rMdM8W2Io5ndSf163UXjPV7dgxUQDqVFoiXVo0qU7t3nahOnyEUEke+rx5fGE3mf
75t9MELJjb9mPt0Fghw5/Z2ctejSvwGFCAfEPiTL30T6RTuKt/ZYJQDldsKHHSHN
CaNlAS7q5cbAeDUxcaEK1kv7XWEf/xmn9dkFywiJ4X6iO6iBoGVHtEygVtTgPX5+
4eZ5MSNM69A3QEzW8WIr3a2XfnowGW9gQwQz5l3Jkn9b56fnR/7eFRM140DUiDQf
VpAmBYbGOWZXMtPPrrn/4ycrkEVC1GapCItMxkmRaST23htk7Qr0ofzhqV/Fvniz
h3yJirpM+HxvDP9WvSystiSgMF3Q0cJYuDpJhYAap7i2Q9wQIps/+Ah9qZx7XzSZ
EQ5sULZWtAaaAh6BeMW86AgbmHpTJb5Zb/PmOGACdskK7Cxm83MYPFEfdRtc301A
QnkoP1HR3Hq1CjhLEi3NI2vAICOFk9zrMhyoUbuiaT34y3Ihl2Naj3J5LeNzu6fo
SBIA3ie9LcKIxT3apCKHZXGhDwfqgzXYM2ouf79/EYeJvpdft+fO1VKosZoFhTA+
714lANSlJ6gLoyDkjAwAtTojYslEAo8Cwbh8d7B+tg04trvym3O+Z4FgKTHZbtYn
1a2si6O0hXyIvN3pE6SK1lptbLVfZJs9L77wWUEzvWXFORYUhXEtwWxvq/cVWtqt
ECCpklsyKeJv8UKqh5G3gVsKdkzdf95zLEX40oy7UIyUeQcASXCAdlPfCpALEs6+
BZJXrYbtpElrMO0pojgdQYWVbbULmbQglxcCInSKO3EV4jsBtm7UBM7Qn3A6M82x
z8eVUOckcYLrZLwByR0yPePf2Zn2beDJWmL1KLIXzBLLamcBnxat9LCOVObRNWoC
UOFKzM16tjaFE0ga6/ygerrdbbX6Szjy7M/Kc0ThD8lrVkqLb3TqKViA/Uc85IRB
qfl0pYyNzuO6pMCDyAvAp28vjpbPuvzE/Fq1jXO9XbqW3rJyCZvSTq0gyiKAb/Tx
cI0LZjHuMZFkuIiZrreyjUMz7qgNPz2BCEWKaYtdU0Qv8t469QOId3FmzepekyLj
WBS3WtsumDf7B0NgX2wrUZWHcJBdn762I6kNDoYm/yAuUg78BUxWFqjiMpghXxJy
X5naGppQF/Ov1o2DNEom7tWTD7RcBxaTPMLL5rzYtxaArig3miGMhzMteogvMyIL
4D5wOhvjbwu2PGISU3E76bupWKEAmw/Yxqupac1y7h/bXjloo0jLQLRqs4K2QFu3
SLmd0aBmH7selKpcJZmssChZyRQkywfvQS3HX86ejxR+jbtUOpC/MYemxcMq06U6
oqfLC/Y++IavXAzuLJoKOl1QmtLmjhHiX3DEzo8LxIKgAqzR4NPuJ5cqvvDva+wZ
aUCfbKO3fLfQvozAYqDoC6XXnJWNd0vhuFd7Sse6xV7CIZ3Ty1bY0K5ZtzoyfOGn
ZYBudNJHEqtoJAvLZmCfSoabXTJms6d4Z0CBlSnUjM1oeZqCg+hJtwgRXW7wcB0z
ygfGN9ofiTxWRC25fVlvmF7UTM6HSMMbrM599D1y3o+Y2YFiYJ0bwWvAPYOZQfQh
cNY3U1J7Qt/ieQGhTunxApEQfzGm4Mtlvpbk7B8pkx0e5lxZYbCwe808W1IeRL53
Kqo8t/T/PCm4A8Vb4ulgiXR+JCOx2fh/CNFvNcbzP+aeAOBbyMqevXnyrDBaaPT0
2fXWaPNlkQWo2ka6Vb0Y5T1iIEV4EfDfplxSw6i7ehnl7lNXE7qhz8Oads9rnZaw
Q9zmYR5wX8mPEumxY/wfGRjZ8H/1t8iZJ21dYZPRFIoriMMhlwmDolh1m6AfaiEw
GcSynGoJmBejmihp1uRD+oZxnYoVU054tWbbbDYQNMlSITvwYIWdYz1oya5zqR3o
3QcGDTTgB+/lv3OKFfWjH4AgRx3TAbs5dUETC9+7c0YvR1cKVp51NwtVGyIXzgk3
tNhIFXixLhSDYg8NXwwA3vkij6dD9OGjYMPBangfJjUfaTFDdnCRF0kxGUsw00qI
Djp/0YoDKYJA2pb9w/iPNSRqFwaqZGCkJnBtlojobr9ZIk5/sMzDM0Dv6Ys8DcIN
drFy87JgJFjXssINYCJsv8EVYh1zduTWKxVoeTqeJ7+YNC+p60mRMipezVhjHuK0
FyoIIaTxqpZBIzG5Ze/H65K6ppqSDfvPx8kvbzQzKEz27ZAxIDvd8pPDOvU1C81v
dxH2EtUwrzbElHZCAuhlRy0tTfx2+AenrIyX01D1I/u31FmB7cAAI2oWOXxRUkEX
P5IkcBthbyumxUlzkVV5hLJ+OcaJsLVNSrxwm2FHR/h98K9e/cEIBoE6XPVTxSK0
sJCvXpFB7P/3mjf+cpEo5JttmUFTfn7+IlMUvfLwt43TXSrt5IGoKVip5cpA58jf
Ks3iLv6mfvmBX3XCreBvQTvHxFy9c4R29pdb8gz+Zq7LTNI/olhOhlpsucNoVOq7
aYcB9oSPCzMDmeDGjLXitnnWtVOcN2voRO0Np72t4uwTvBX+M5mzpaY/GYOh1Zje
k2/19x2BGE7m6MX3X5GJXvj7noTuZk4XZnKKZ6Fb+xCtdsPLFhmx+XhBRccKm0m9
nt2i1E/ecA4urRfcfbyF6nM+B/C/Zw+yhNC1Mp92rHDg9cJKrlkCQM8E2KHVeEn2
LCgY6jSr/deISExgbJR+uUIPgvks9SZLcXxOJ0V8P/VejzCIa+GAlByz7CgSAkSP
KVzQBkmcQrS8hw+A8DlL1y0xS86L0+TbJC//5Y4P+/sW0tDdfgijYImk5wQMrfQ7
5Jn/JH+osiVxv7ONTfYV5/S6yYPkkoqqGEvP3CaZuAiJtqsS4YaatNRzG5SRmFfZ
OZj5po4BenRFBQHLj/VGhlkuB1CpE1QWSAuKrPxOsW6u6teVGHZTmQAjPQ9a0W/B
yEcYkcsqvohIBy7Sp2RhUzvZTBlPbHyctQmXQ/RnY1FD6grrlQrrxO6GN0A0P1IC
wCN3gB3umcwewIXyZk9HIvxJI8gpn/nZSO3yFtEIT8FY8rLF96HYyYUHU0kRCFGs
8RsH0a2vmEmFoonv7BFkiDjZlj2bI+lccO3QBcN9r/tapX/P2bXARbGK2D+PXdO4
jNWxUuKKB6bSIuG0eZboFxzShEufwolTjb1rXKT9ZjxFDVMgP0OBUVYgwxVZiXNY
+MyTQSEyvnHYDrrN182x+SZsf2Bv0dw8/ABLwD9S04vVhPnRVVJFnJJ4xF+FEefR
ca6Fg2i2y2GAmVI8ioQX5NkXVjezfpahJ9CY09lkhg2b9JjkPiqAwAFSwq0a5L+O
OEOBWIMjOGvReIDBHSiDV8oGYMSI7yqbM9FURy988MXYcjIrpSCn6p+XwFizGCrb
9h1h8wNrMX7nIOz71uaap/cQh7y5vw+wHXW/hVUqEQMG1eGJocI+oyncuK8r4CN7
f6TVJNZ7XRZyaluvdLp+WaB1sI85YjgPAf4bvp3jc7ut7sVfXA2Y4SU70zQsx7qp
jBFBKhEs21NRY+DL3jL8KhTCo1cApis8Og3sWLYkXqNAO2Tt88FuYQgxE5sF108n
9dcank2Sd3GEKTHdYJrgp4VjBFSaC3BNy4FWhlJT7emFBm31aLHRuMmBBhMaLOTf
ZDdWhlJZSCjtTfcS3NB4d97ju0JHyaKtJerbpTAm712QYcIlRl/TN8p+14CIoKNa
sAAy6Ff9T8vgw20JQeMjrZEEWDue0dr+/vZPHwtTkQcT8+p6tYfMF10yF5efSmIa
ipccgRti2yNNqexS4ynxuqbYoKpr1fx10zUVunamDZRIWDpWPhNZ0+IeOPoFhDck
XrANhHlF1l38ldO8qunp2W0kgSvj1R5HEECA4M1kK+B0zQLBDWjaO6iKV0HWtzO4
TURFiquCEY77y+OPkwgDvkwgTjHDNW5bj7mLAG8HUuk/aZ8uEdTOfX4SWs+m1jLM
KvXjpLWIO2JAyi6eYjbZ+L2/glQl7Oem5ClL02t6HQFZ0hTUmAwyWANuGMdRTj6j
ulmvcWv1h3gxfC99MoLtJVeHUlxKtVSVYAXUhiaUa56quAdu1Y3ufLRb6YcWlCsP
ztO/z0IAu8dHEULjef3VR7mfGtGkEqnU03BO/TJKb9HvmgZ/5WP/D+bxytcz2G7A
szbkkbBvhn2Ks18fi9noPwehjYt/jyEFZX7BoTgDPh8+9zR1MD3Erslytb0Kyj3A
TxLvR2i9zaY23iXK/F5xR6MkUIzw6JySeQk3mZmFoiyiFooLC5cLTnMcwjsxcbp9
WvxWl4L3J9TOgE1/9ToSzmWnpUQrNvn/kQEP34mGl5wGeq1UmdE8prfnHzd/V+RC
/cxM8RhHCaPUbXC+z9nUAIg0wtyvKRJvHAN56xZTI2S0s7yXiNksRP1zV5hBOiRV
YbqxUKq+gMLmKRb1ayNl/engP5jXQ4uwj4hB0ieNljqFnTLT6tevvDEJKHPEuJkA
QOa88COPG3+p7DYHtAAZFqtWhwok5XKjPcbCxYn3Ebm2V9vzm87rf9wB9Xdq2hKs
qr23zEaYUVuhdwNZb40RW669IjPvFx69IYrMTlewqHSCB0hwqxdH4nWlzUNryGS6
oZWW4v0NUkb3QGqMMtWghqRvgo8NQ3i04ytoyQNpLLNvFRee65drJQ5zQxgYYXJw
u4vVP7b3MACEz/Uuwa+d4N8abXL4JCQh/dTAAl5fbalGGiKOq84TkQ+WkA24EVds
eQ07+pq7qnoYB1i4YViGiS8oZgJ6kAE9LxRT8jq7badu/bR5Kphwes4359Mnlr+R
CxmL03lF9PjWzjiByUD1tfb7UstS1OEMtcFYIX1n7e6VAm90w628iVRGU6SUa2h+
GhibgW9+JRxBcuLJJB10VhOHrFsnwRY8+Fk4UUqNYXXOu0bXE7cdIpqN2XocMHEL
VH1//7+2ObxJKS7Oy75qp8DVKyaiytr/jyEOIAXwSuyo2fUZgYX7hOUqpx3zNmrP
1aDqAJNOjnadtpnIwDK8Evs3uiiFzsUWJM5LieQr0pM+tVQS8L8SbXJt1DvLyvDT
DH/QFW3W0ENFQ1IvMs44g/SFjKFjSYTBMzz/e3eDn4dRuh0D8yboJMIHPNC7PytC
dx4Tnl7wkyQM8vlqFH7Ea1EAxr69OBXjsINpc2gTNvJ6DrCQuo78iy+WsyMd1YIm
AyGnuJUoy46nDoX6hZYtV66x/E47SZfWUAGbVSyq6dv9XcurPOlNxQegeotUHM+6
RZ87BHLWC1+bkJcckP0I02Ix5a+wplIOSiiaJFmOH6Vuw+wt1Pwvs/YAWbwVVwHT
b97h/5NzS6ViHhnOn8ZsUMgALuazysbP//VUHy3T6hVhEO7AO88Dz9kgwuqTCT/3
5YOL+JI0rYoZvwySTrTpKCa2HcQhgt+xJfg+V7XgrIkM2qpG2tuW86TB/9J4R/Zn
dUWEVyUOiOTZ+XYHGpyUcmAVRlU5d+80bpWH1kAooNdIiDnJaaDDQQX8Ta2Oi0ps
qEXo4yIRQm6ns3fP0g+Mi+VtkJAuwX03FYPrFRA0wa1yl1rWZJ3cw33A0Dm16eo2
isMbp/7TYW9j3D14M6v9OrEt2M3hgF8MmYHyrLYPAj2EDuNAMouzwdNllqvoe2rR
2T752Tr3aOM+viup9zjmqqMojQvOwLZ0kxKNAynz/3VeaKUMvE5CprGO+0bgz3Hq
DiN2bn4DEYAWBoDbm4F+fBwM9TW0zhhZnaIteUM3atvyebruAx209PPNJw6bBBdz
8h97R7u4WeMo1Uzv7M0E/KwezLGaT+9V7JIhu7EDxKARzibPibIYhHgbMkEEK8mM
OOj0/kAS8OShpbNbjBh7MQfaJKttpUFvZSnzU2Nrg/YJQe074FKV1w7VOY5MDfTs
zFwlrhT519CoNSo41yLRFcA0XQcblHmYJ5NFzLEVeWJbxHPoxR2JL04r3VaAOk2k
B1RpHpu3+gLOf1ew9s97vCVYRDJ8ygtcNHhX+5xM/+qZcrCGfQZFlDevMvWj/mX5
RpaE3due4JwIjhV0orBiCGlD7wW9jFn9cjlte62QrzmuLe4Yd8ts6JiKBQbHeUTD
cdfVKJg8ZGsdCNDJEV393izK+RsLKYaO3BgtbIrMmL/inicdhT1ZLDyo9wCInTsz
+k/zIKaAg4erLC4EzlNWkADE+t9Jp9a7HampDPNwnjt9Ybr6TbfG7yG51cysv1er
t/YECJ+EQPOVBKVfiz+VVuhwCMbLiEulms6TAzVAx7FVDMTZ3JSdTBBHKYrwtAQc
qrKwN4x8oL1uiJ2nFV6pwaOHbUCyEVERRVH8bKfprlNRtl5dnG8GTE5+YEN0sYmt
FFQT8chYkEo6F1WuwE5jX9ure0nmQ9N5ER/Ul/EsEZGaVF8eOUZKhOPKuez/4I+e
bUonWlFQjeEjeWCrI8UaYSEXKSUTdrReKQpjVoLXCQ62pp2bjjC/pqcznsJXfCYu
A87BCqxjZmStqLF2NE/HRaSqtw8c6Owqfm4hp2TJoDxYCaLKKbFzEMepxJbF2jc4
JumvFkjxob/98mJGTpQ1bCdQdk3psfim+zLvaJy/FZ7QPT55XBjJZ2a1oNmBkxb3
n8y0RShZyqt4mclAjte6d93wcdztJprblLLPiks/6cw/07gRy5ewtZ5vRrfe9srv
TBhb82IvHD7qnzt4msJvop3QrhKlrVnJ9i4bIrFzluUuz0KNNNowUaDHYGyhm+Rj
VbeIqwl+ew1jiw8vSiP3+EWrhjt/KoA0vbLAxc6eugOhZdJ2/2Ai6JlinBfIGKV5
aoJEnPLWmWwv80uNxm9dR1KQH7hySOzHevaNtTzKxrC97e/i5ZNEEfLkFBOQViOt
xFSQM5kIp7Z4mSZ7vGR10kIn+xK6GLy0fLtT5SeRWki90nYuvWDs7EY4mJfaaVrb
8CwHeMDB+qmUvb3I0dyBxnwp+rwGP3trbe8v6iG6M2D/KfII5fPhD+KhbXnD190c
E/lD8Imii6UMtarfjtTlKLPLv/t+m34swLfBpyNZML9Ai64LkvvzlVMbTGTJ9DYQ
7iJ9PESIsXmaKBdJA+8R3pZRa1CwFETOu4Xdin3leqeCSIaBypgqbG4HJq3NheC6
ajP23wSKJnI8IJelc9gj99pZCP+bRlzHTZPWl5Q926JpKNQBrvTf5hlfGdR6V0t4
g26zjEGpnTdmRcvbqbth0Y52M2oEOFgQOjHmNE9FvIFjGoQW7oYs035asFfLSNGX
gnKCvh80mIdfPMKdFIJ5i3cvUfW7DnqYb2nhfUxzcq9zwPDopQSyJ1KYjFfvTT7T
7IFaw+r+cdtrN70f+kvvMu+P6WW9kOKkvXN0qPDtVKG1jjyEDjmkTR8kGuOJppFB
E3HD5HzdjiuGKGZqQD3vm+LCn3oi4e3Q4iEIbiy6JMF/7r/6+ZGiDleSv0z6wy0U
LzdL888SorR1ghmMYQW5jckG5Z9oGkxNV/7LcGzKTBb1IoW21KJuk+dbqz5zUzNo
PXA3R5UYcm+MHdx1vEfk9J6JFYXAmw1vtuvsIZzK9k/pLHK8T804Xat75uK9Q6Mc
gOAbtCl3U3sPixJ3S9tifHHdip1xsIE2gcotYdjfOhGQNXmH2A1eM+D/6NDNt39s
CPmV7+BiTtARJ735czsqEBRpaQMY9jMqStTTsPDJrPYJ++d6YyyK6l0K0m6EKVWt
zJ0wUDFw4UIAHodWGObz1Ye8JKgrCRJDKDb2IKPCLkeVSlixBD+1+WxXuMGGrqaG
DxL1tHsb1TLS/xEDEFr+s4FCWQu7x9L3Kx0pKaOq4uM4fMzj6xhNeVW6KEMC0AhT
LMw1BQ8oheLB/t59GNjD7aC6lEEvwV2FCtpDzUAdToNsSDjPgQmAht9UtgYuwFBZ
QARxjU/GpVmd91GyFq+CFXNEYudcH0V/vXWvAD57O9rNFvSPtM5WLSD7yXpXJHQs
tjWbKx2YCPlSY1Ontj62QufR7DOM86fSzJsKxBaJEqvEcZQh7z7eFDiklH1dOor5
yfrbd/pqTNBK1xkY4XUV81vr3wZoZ097xd5WjbfRwZMfl0VuRGFMkdBCb/Q7hadI
gLpcofkScvLCfkH/7aA9fxSMMWlDXtycx8GJrwhse0KcFMnNIz0eLGadruRmfnE/
WryVOw32hrB85G6LXELB8KAVZQwH+zSQ9UB2pNrJ5LrAOPkYqBDU6acxU27IyOIh
b1rYqr8N9hz5mTiGGfLBBKbvJ/jF194843iVhhLqPirk5v2sS43S0Rhmnarj/qcA
ePQX+se4nmz+6CgYNPWeDO4c8rbJS0TmjlSiCFwGh3l2EoPoSe6ObP9Yx2b6Vz/R
ANqFf+TuqASlqRoOY/YlJoD5JloSHqDvlWrIGtk2iz6vO+UCCKLV14+BH4NYkcy6
5HJOI3nezYdOlrbpZeQiJXnagYRRBfkmp8l8cJhF7zdzVYI6unScWgx8Bk6+swuh
j1Nx/Lg7+ykFI7EtS3kJwkn/vQdg7+uFH8Q8YbdWCThulvlTo8H93C+5IZqcZ5wD
8tM6r/RSSF6q167CRZPAgETNdSss61w+gLuCDbd6hP2UUFFTxZQSGjyaSSpKWfTt
SlxxUoql6liZ+Sgc29icODC2lKqxqK/kLUHFszzmNrcDdtTa1P8HltiG1WNGZe9E
GLNx66puXBxAbzmYgr7VviA6i1Hwad8a4jYRcNQ7mmQ8CqEiqp0aggKHtQ707WPu
BGA6GvO83x3kfAXFlI3LGyTpnKi5FWBLjHjyAOFmzwCUdaWUIcktd3psQmNMiAcT
LnYPUufdkLvaIdoyY4hsEMIaw3aMTcVkOxvZuQg72CPz2lHmx9U5WE2Pm9uL7c3+
dhIOHH90F+cXxbLrlGl5iVUKlaz/Ao7j9hIHKc2e10n18bBjl0i2Fjw1Q5fOlHQo
ar5PqXZhsvZH5JWVNuj3yEGdTqIqIElXdiMCsnid1yyAl1gtaq74tOrkmZpDZVum
dN7dQvgfwIbS/hTFM9qdqmHF1UWm34wta9JG+jsRO4gPAVyE0XPeaDYO3yNDqIUC
KYsrpcny8uCrktaKUHQtV5+wMHSFhuQtvfPGFTPiX7GUsiAizHqXXZ8J+Sc8o+Ny
Y6dnhrxb8WEimX6IfAf7917vqbO21JW8qwXQbMOECYeTVinv4LBAkgsP+9P329y8
IxS/zXwZV43Bc5oTLVC4i27AgXPLFIccGPE6Qs0s+bEv0WQMGgwLcfQLpcvu7xYJ
XnAPUPdXkox7QYUkPVslOYV15ro8Xd7S7hyFviGR3La7gdLCVWu+RlOMcoanuEif
BshmRc7Zfmk+anVavHdC5ovBH/b+0BJqHzR86f/AWpAEfq9FysUQuZiS0IwADzV0
NvtwOk+JEPOSKTMUSFaGBucz8WSEeJWKdUtibpC7C4U3g2ifamTBrc9FWZapabic
Is1IJblJVVY8d1yicsvIvewtrUBGOXH4Z2uw58BCNYSqJlQdJIddgaBQuV5eTVeE
0NDO+16oAXuaSyHGD+x0Knj65K+9OmeNxQGPmZrJnwVdclwHuEBqbocl+A/koaKt
UrymPzE+9KXBsDGvtv9SqJC+4DeQ/qg0JyAOfoplzazOTpIepeN+V6JbjX43yBI2
kJWgCJZsOWcubp+iisY9FrK7888lJHH/UXVqX0BGl3YICBsZZkgcmXvLqHuFZOYI
X/C8H0UH60yrFvf/HQznWX3pUUtY0K4Vsn/1+ZLj1SDIyL0QhHCTs7O98oYsAkaU
/x+b3lWc/kof33OIjwR9dtiJuJPkI6AjjsnMSuiCGr9CLS44IzGwBQWvbS5gDbUD
5KknGjtjGHfV7Z9NjKa9sFfWE3VPXr20ASotDrxspYXPrJa0zKHc4D6eQZFfgUPI
A5rzN+/O/3bk00WIl386tFppLnycy2ttL3ILdb/bVDKKpLWfEQu5FIj9ySiv8ywp
4TfWoQzbf1aaCK3Nlpq/5m/xZvTzF0U7c3p4KFznsOJgzkrJld1VL0ipFOQxd/M0
6oH5I5PFaqjYuFi6XF3WQ6TClgk6ufT+3cnnhPts6t6ntahsiCsgdaraqc81s2Lq
pogCooKVWhE2v8UE004qKS2ToVmNMWj7Z0VWXEm3Y9ZotddiNB3yG7CLmHABXUPt
Fp61WSpCMq2cBIyN0fRHkb9OoD45wfgJ3TyZgc1HAjKTYHsJLrs2Dmogatw+HNNv
xGShA7DgoNuA+b4+8pGtQwHiiI69keTeUi3BhWOKE0ukq22QijH7kb7Ve3UxPqCf
j9jtuPfJ8BzSNNM1vAr8pLZkNryuwXuurquQ1qStL04N9B1swmLqv+J3gEPji7DW
jUF5vp8GAv+ZVXH4stewca9u+EzLedWnN20arReamEjUvuZjJsb5XBMYbbOSwtVY
2z1QQVGoTn0xcjkC42P0oTvaV38lXI1ZC2Ss8jx8m8S0tFqOWabOWVv2K10q/bMD
CkpkzJAmDfAf1mWyfhL/O7pJPHFzv5/UzKcLFkmLsnVIIUlrWbcFOch6x985TwXf
yIP4AXhMjO8kbejx8eEyStdqWhSVYVeGzlmzjw6n2XdUglVLJkOY21YXdAzUSEAv
geuQfy7XMyeB2QHlZCdE9niWowtLjv0IUro0q/vFuMBv3Bbs2AZ180jojomi36N3
eJz8eEjZ+2NYBOUBQGNIfB/UFisCGgAvbWiCi4aNPn376oSIP3XSSmA68eLFrrR/
qPg1ocMa21T+VCwDNA3zSVdfkWWxgMV3/IpASXwZh97jRNID3wfGlZmOzGh9R9RO
pa/sKOGOeuD41BlK2yyONca3jtO/om4LFp8bhlxLaXvOg6gCacOBd5aTMFhchdpK
9MLE5uV4hBJgTd3s+4beHuhJCLfWthj7nEQ8/j9Bo93nH/GNRqDio9aiRiJxhwAa
Q+Edcn3NJi2bCAg1zZDULwRIyG5nB5Ld/2lN/Npmb4q6GUB10/2JezkWA1KEM+Zl
xZRJm79nRRCvWzx5FpYHQOiBk2CLTNbdZuNRMwK/FKarlLHRvXDZUlImepm0XLOo
I6m9VMv5iPVHYaoIDMoaBTFkmE/R0zCpDGkPZ9O5aTyowCIPsIGrXynpA26XtBQt
QUtr6Ybv8Fs5gzj21WFUPd4fF5+p372f8GpzbVdw71DT2NzlTsbx5k+buFJhiPqO
JDssNVa04jdLrk2zxmy72jD0M7A4TQpbTIBL9pEJaoIHWkpbxxpZv6b7Cs2X8/xr
S3cuv9QzXTW6eEF0E0CvRUq3ZgAUipnWWai6ZoxYddgercmJ0MTGMRcGA7cN026K
DbHRAN3aotqNtknFiE1O4Rq9se0pz5gDs1L/CEAUI71ljpB44guRfB6176YFqmB4
x0tRymLC83gGeEN/A4OXLMnrq2cvwoa135N7GoCAzmjyAvI3L/F5+LOUtYEjXFTE
4+dDdisFryOKTMkhY5tjTKIYKBE/rlmBBVkrbEaZMXn74gbOhSJoBBa/9VgUGpka
nTCbuxjnt1aoKY31/cC8njjg5wg9Tn9Kyo19UVPb/sIyrJQnE855x2I41dwNawcG
urKRmQznPiAatAv8rX8PRMoDtohByejndc+6RlaDBxLZ3DgzCMOzweMb43RTronY
z/iIj7KWFDW3qFyI7BURFn+THTuMy4nF6vA88HTuXmD1f6ZUlfVtc7jY53vi4WC5
dbkJ3zey1Nh01uaj1jfBru1mFVJkmnrC4gjnEmCzSd01IUBsbpqkvwqsg+KQNmQM
jEKttGicrz5w1nhjRP+3dhC+z4IcCYV1BaQp1eq6swrwrM3JaOeDjlsuDZqGZ6Zs
3SRlAoKGk/iKvsSO9RGmrRmuJ53c52SrnJDRF4icYvB2U/x493o4+IFyuirk9FQV
sEAwBUv2U5yeS9aF19kqAy25VGtYW9CFPUGiIcDugsINOAXAbnOKlm8ERUdw/hWA
bQbkp3bUok082QI+MyiWp0eGvuduuflLSAbHLnToGMlv9DIjBWoMURSRfixZy+/V
vLdJsXZNk73e6r9RbK1kQj5u7TyLFNOY+k1jP5cxklexGIQShMbrsSnNxkGgrpY+
uiWJHbV1Dpe/OuoC9p2SWiwiGr3GtjR1gX6gwqyVJOeAK8ApyyYsZQXFHfvgBj6W
bJuUh0VYr6sWqil1KmFmFYEHIBOM7CG3QsgnoFc7x+5T3cLYEovchqwPpR142YPQ
qQ0f0ZLBea1q15S4G8ZdcDGUxwq/fKm7BycqDgdEk3hMdSDthIIG/3ROndwRYYRK
HPpnQ7TnHPBFn6NiHaMB2/FYcMn4l11NwXUEgjd7IRgx3Id1M2qvnk1w5E04id1I
EQ/crEH/BQQ3kHaV8Nzhm1Tjw+dIhcxnxPvnqWcXR9tImDy2qzLGTg5KuQSkSNHZ
LB8V6voPDZiAN7U0ZAQ44yMu12QRnQCkrboMpMQtjZukywZMWDMGLlMqxLw8upK4
MjzANn4ncxbW3JORjDv4MGDtDudo/4veQ+2MRiZuQ6kJLnuXwl8Q/639p8ThL9oE
/8QWC4SnIgFXEEZzblNy0Us/502sQNRQ9p+ksjGhYMR5HGXLZ5/1UuTnhtQpgEkz
VaWwy73Xj5t0lqVqC06PQU7h+OyoXxuHtxayAnzv9Un7vvpiyVuo5PsxyGfdteGr
6E9cJUFG5dD/MnSnENNJV5f7mIHmzQjh2UduqXfTTMTlsSZcPyFys+j8S6jOWKGH
I8tGzAa5prqoauRt1KSEMmU77zX4ddgSmpzvXx0lHZD86Pr//1pHzhoaqlM9cnzr
Y5o+puUdvj+9WwXzmBPmWEQBCk4/wd3Q33yIzyHyvQ0G8z65jkSuB3IQKJW4IUoB
AJOIZg3AjBs7L+CJCLUPZB+ty7CEfBOT/CJsOMjH0svrIgK0+ycYYlZHIW/F0qXT
CUmzoRC6J86z/7lyq7bRiOMv+PDb++jX6neILAnjDkvSgficqJY27/H9/bj5V1db
M1xoM6ojBCGcWpC4yGrNwKk3TEsbMyFvVjqM81UPccrVk7sxJD/NL/zGL1Ki/5Rm
XMlUC5IA1FdRQJjStX7EFLTYaVLPouMQsTDQleeg9olYVAkmuT6Cdiv4vyR02aaY
kelvfPWPPf/6ew3UXM9ugQ7p5v+MkR4q/S8xzfp/7vv4HU8ZAo7LQRfR53HRtTPW
MO+NfrQPKcMSpyr0/bUSqYzzvTP38C0SAdsQV+Fx+HemxPO+LDEv77+UZp7RCqA/
KTdwXZGOmTxsxwyrLtldXp+eRvH4jNQIlBDTOKkjPCc2gPEgbOeIogxhZoAlSjOU
PAT0NffdZcW/fOmXbwBQAUQRPULGf95UyGlbNPZhvoVmT1a9YdjSDFfFELSrhl+y
wCZtRVUXCFFtUO8TqhNVXk4BFLFzOvzS7bAP6gxsmg0JEoTxdOXJzmM21xq5tmvu
Y+A/TI5R/DGS14d4r2FWcY7qvKu4kBPcgCEgFjL8ZgLL9Bt3zzREr7L1jQoIuUGs
OxNpMaUPoiSTrN7fRfv55XjYaJui+n0pjR+pdz1yY/8bvtuLA6Xm0DosLHig4IVI
xYv7/fS06O+eHHX5bRiitNChrTDSAMspmV6QbyaKCAewooyGuQxm4xoRDvJNuXRg
rNKh/mphd0Z+ASqjWPVwl2EMoP62RfgTEomaG6gQ8VWuAhM3g/413kxgDnlgQ+Qc
wgRth4WBNTk5syYkKD34aCVUHzK6nHss1ytgHGh9Ih7/kJE/qS4k2WsRd3av/pDg
/n6BJuoXAQCJSxBFepHXvQ0NXkz89V+XCi7F29eJmhG5QswH4/HNREUqL5qO28Ke
N0RIv/TCbpq9HdxVI7Bxh9DIERJqnGNxO/jWjVqw+YXAI283NbPTJTm2eLu1ig5y
QVZx6v0Ctl8SMqWDVLIDsufqAglQg8V6G0stxrfrex7t8uW/FxG4V1k67OiHtnV3
7zkS9lHGHSEuXMPK19vpmTOUUAm29h+8Z2SGsJVUgX8blD4a6cx0QBoLmDKyaC6b
0oiuvOL8APBqkQX31wV+AV8RsYM+8fygob+xNgCfAt6dffLYuK+QsFAfApV90amt
4ckR3Y8yKWU46wprpe3YjMHNCNOtd+4oMOZabAEiRwNiEw9003MAd4YGuESxvQj1
4hYF6lZxet/ha1hmtsH1OKIce+MxUzIQx6+Gqxb6nhabiXv6kReRWdWKF19JSqSL
nj7SKJgd6rs12Y7Ze/+RpfP5CBEBXRNrwP7TYQ/S2yNUROYdoDtwHXquXI9a/kQZ
fNrfkzKoTLY62iu1xeetX50ODfHqGPCJ5e5TiHyZahqdfJGCLcP1aYpdmSP54OsM
2FOdZ/tV17zBry2ie5slIviPHOLS0n1d6SE5mbUGLclGQJKqgVJCoazNDd4qIIzf
4AB5EGA9YtTiL37O6/YPqOFvMwQ3YEGz1OeqelBhntPw5L/RZP2uF6VlNo4a+/OX
l8elZbbfEZhcnMcNECm9sTaUrqR+cqNl49oAecnec4fGquR2At0KIV3MvNtrAdAf
97kEnhhu4lEdmEJp2/ofKIIBvvcpSNbpTJsQAFYI8wjT5C3h0HeiQOG0UbrOvtAn
6QBGR/DARTdPlBDdt8hQzNekqlLBHhW92fvpGknJbVv4F0ityObcVSM4tKUNoh5Y
cC6CJGbV1SXWbJa9SAbsaLxHpwjOC1tpHXIVX24A5QCyXflLkyJqkBPlG/XOuZ9c
NlfbCj9iPriHUr2OSH1vVOIkmJ95PxjzZdLs4pC9eLzcSjLPkdqciqFoKErKBGYG
94Dy3Sgn9mq468OGcm3Q54h1BvOXG/H1bUjg1h4MgnEli0EuIlvXLUgF229CktUm
4f9aoZuR1rdpbo9wyi/TazqsoJ4pIKlPZGC5Qmgp75innQ6/Ify84GxtTdQaxwhB
lUN+qOEfFKRKdGny74ehCBaPfwuD0oSyK5NB0V3rQcN0mLFyU2jM60UAU0Mo6EKm
ly0TOIEBqqczMdolcYsk3xiI106/TlDyi4ZuTLEEr3DM4GysjBVW4s6muQCKwZ+U
Kmg5+D+f2xcG8UFwX/5AcmGunG5sA0NC6cYOAYs6067mavvD0lT9Z2rNQ4TE9p6q
XTFdzTYETmrahI6xWhHWPRyLNRRX85DJPIfIQYEuvvxOjta/5SCQadZD1rrwBcXd
3j6mogsJujEmx305EZbPC2pRLYKrUr1swzeu7dFd/fGe1IVulX44OxG99epmZeWQ
BbTlO1hV9xb+QhEibqbTTXRq/kEgoH8y7mcy4a8DAfmIz18OZQ+kjUM1Cz5MGTQ9
sROLdjlXTPQSqGTChUHt7Ep7dqmceY/qZLK+IbToiiUMYB4B14irKU1s5nNH+ApX
2pd4I04hEU2ccfWlueN1I/smeBLTiDXwvjbnKTFGaFNfP2JNI3PEjAFsla/rzafY
sETzTv5G0U8+GnzsxRruM1uIxuO5QrjtGJda997xPT+WTNQvhzifPkG4AlG2PsSo
h+qkHsb5guUbJv4BVX5/6XoA9ZR2W5ygcz3cwQRQF5NhjEl4BS9OUfussxu3zSHC
M7XD47DsnAHtIvowVRjgUI3qesIR4B0QwHmAJ/tv9pu7wvEpZRXp5fulksv0DMOE
OBwPOUklHCJIvzCsPObxvvm76a3wC9T0rO/oOgyF5rdHVgvRDaQIfGBVtxZ8BwU5
J31pWdNYdCnFfxO2uXw1a4UD3vYV0TBumK7s8KUx1oq38ldtGjrMA+g8YwsooayY
op4NCsR7NX0weQD/Aw5ZWqvl1g98g6+1lDjJovTs5OTIl+UylJ1qDAjhNXhbqqdH
kwXVKvwd8KlQOSugk3a3BOq+dYQPKJdaWIKuMt9J71Lmvkc+Lf9sKxYrNBUbV7fa
eB7Ub7gb1k8BL7KLGmszjgv+LjdFNXZYrwNRjCl2DJ97NwEEmFNGK9DqAQI4mZ6I
v+zqEE8BLQ0yc7PZBTMk1NmPsCqTwmI33o2KjudRl0Frlk3Upjk03WOwbCMe9rtK
85fNrCVhYWbtozeCS+UzF0t1vICu4lJPd/5tKM/P/hyi5hLb7S91R6RcTaLoAz3N
4ec2mLJBzdFzEKs0o2b8HJ7J8pkeHVoJvO6YIZS1ErFBmoVAFu3LJtZx8JKJUuUv
R8puNgHloYLD0tITEpP2xohDLiDTm10++Yt90CaSWOyZkkdHyz+zqq6kt9XBTSKR
x6GIt2Gti7mZRpwBq3DI1goW1Sdb/ByYcLcMpNidTNhNTuEapijJVEOx96fZcmAj
wYu4HM5ecBnkeUelQtroZj7y5MEtNyt81I4Mb574YhtAhH34OWnmQLEsSuo/Av0M
IyqjsK3qjV6XaA02b3ILhqMCzAww/3FJp086owZrpQZypJWrNUltn/1BIzroMHcB
tjAFJLiLgKw5sY7sX9jPZVhjO+oGMtgri8QkEd5qmaqvShR1MIoJ5kZJaR9g25cu
ZW+UMXeyjZbqM3aFJWzcMANbBaRhAdgvdsUogFHJAnr3zFgb9cI3vB54WRTi7P6W
agnC9luc7HvrfkbrcSw5gEW7zxUxNVAH0WNMTYVbAs+T/afQ1P9kIH4b9rATRs/x
fB4G8DUv77zGkzRG2ZX46Rxk74lykWxPsJxhjiyIpn7afOf77labqLltGx/MayE9
A4RFf3ZA2aWsP3V5zALRRySuql+Hb7XNaLuynHFcFhuit2hTrr+nmSIjiJW/lxJv
ZJCR7KVYHUoZcPmWkiuJyqMi9OO3YdilBcvnCQDIH2/cUqttoUFe7h19cOeHQRYc
9snhU60bsaSL5CMsFPTNsyDxqrGl+FIuQCLwqSDE0kAhuARhDCvIx3Wb4NcIkOPU
U6+g+wblOnY6iDLKLrP8MFEgvLzCFL+t7l/tiEHudDlp5cYywFQhtA5eKv75Rtu8
RRva2v3wA7+NaBjXLXcdL3N0fS4VbWdX5qu/chT/jmtYG9HeTnmptIOGuF5QlHpC
tzme9d5Cg79T1MrKohp2kgrCvWfS2DOG1keAMkIP4j/h34DaWmB/Cl6E77GjoyNE
Rz0rqmhFilmcqlw8Q8iOGe3DiYFmkP0VSX5BhaX+D2ACcHUBS1gB/jJrxBXAy26L
Yn0LwyMAtpxRO9xsDrZ7k2p6TmRQYGbt2OBYkg5xN4ej/su9dDpvWWE2FUtotGjb
jYzOHD7wr9lntC+2H2wY08vuyALk94ZeD3ZDtJv7TPiH9Afa2NhUXeeox2w2gb0m
Rqhjjk8j7he1KIGhWjM7dGb955f9YQwOJRDh38i7CumWbYdW/hb9fklrjJK+HfWv
y/3JzkpaS/xaaT3M2b+MCO5vL/FfM5c2TCh4TnAErobSpp9/9wc+9qbq+G2H0cfv
vfYIWKUFy/8dcwV7d5BZ025Xp+kNh01p/N8CItwXBcZct0L9Ye5ny2bFc0P6mAOT
YaEFMWahOAvEbeWQ9ECzp+gaEoMLCL0KYF95Im7cxc8MXoL/DYe3qdvQGEFkHuEX
xG/rjw73ilK1u6+1oGGouVb89f0s4EKdGrXKFCbQWaTJZji/o5YJ3/dtqva16zCv
EfUMKTWxnd7/alYaVbYUARerUbeipUfxA+xH8BsjsMw8zAxqa6aAdMatQBpL+YfI
jURPPlWEOuIptpaE0Zzht4Am6iQmDKU0NIRBxpgPSwAZKV4/ghKjYrGQ3GWyf+C/
dESqvX+nen+LbHs0ztsOppoWaO3qKpmjtyiksnizFVqj7cJZfecjm7QU6hb+PJ/j
h+2OiTnOtOARoC9/2xkfN4u+HVkCaqzJgpU5G3UunLF3NNQH34V4mG1wBW1gwRiP
WHYE5KRx62nAT5RRGIbOHTRs1nBARZsfwf/yQFxZwcstJ8FpCB1jimY+tqdZrdUD
23eKQjGpEHXjh4cQt6JN5ITNGrP6HdT8KpU3mi6iY/e8NnDF//Vm2mybZ7EC2Qak
zJ8xewxZJRqD8xJB6iOMU64lpkgDW8TUP/r6asfZwhPES14KluzqQvOsyMvfDNMl
Rlux7Qu5iHuP2QW9BvHwkrJ4+8fxtnI+3S5CbT63t5VvujGMIQwCmoNYiyMti8qs
XrTCww5KTHX9rD+Xx36wNmilNpJmksjRDUKmYhArZmizSUrhEQ2VIgQxT14Ik2ry
YvEhPieNquiqUk2aUES1jYSBhP/bK9ssv/djsbpLpmkb5gRxnpYzwn3o5uT2TFI2
Hz+Nq0sfr5SZhSbMAByc0y+pNOZCnkpqN3LXCA7JLPmlAXchT13BdthFxguXF870
FEqeYJTn7aVfRxmtPzs+GBwLGZdJH2FuQ11nql6ydOfT8cV5aFJQjPWJwCn00V5Y
6xmNbh+By+GJxxs/43msZ3oTBvQEygHJRpTZkqXAEEIOS6WuLPwepH43SwuD9EN+
d2GXam7iyXHJhMsANt+HJuu9xGSanLhhPEa//amHJf62wvQ7VRTHrzRR1MP8GSuk
kRdAKy06FhIQVUMPI6lPtqrO/gft63euRBsMJUhaI/AvvquAmTqbg31bUoLnlOA9
94sEbuOGtHL9rC6a/8kF80DquFY2+1VIkR9kQxjuw/MlLpNBuB71ojmLOseKS6ju
eSTkXf4Lx17ln5hGbgIdMnr41D1SQB0TOevcTuLt4A9fALzALuwWCBdaFbxo16Yi
UXqOl7PKobczqsn43mhc93bBFScwx8Wu61G8X1nrSh5p+i7mgccZGHfj3hfeDnbW
bCv6+gT4ZrpaHx/98NYawFLFPEwZofP1XzZUdIvKqFUhvtNsVzHPaGl9lF36ApIp
0xXuQ+VkVBRRj8KW6OqkyYNjz9TeC0nEs+TLTq381w83NsDuZ4Rgsy/DfQTDYxcy
LB6q5DT/wSOyRiMRgPjbFlKU4dMeAU/OiL9fg19YQmtv4Be7KsLI7iE2ip+be51H
95FSl8TYtcrKaU4ddgdxs8OfuWmd5wfti/Z/Ev0TTWxXXcJk4o3qxso2C7VS93WE
fu5YtxeA5haxJdWfCBlOYf3wXLW96friKGeiF2kRfmMxLXkrVPn9rgAlS5k+SdCy
CJKjkff7hsj/wjRYwV3OG1iv076Rqykq6z9EYdhZkA+xXaF76wH0q+ZvZHbAHU3X
Lk3mA+COnnWwewUBqzvmX+0homJGPtW9Xh/M+BCStbg1K6bpqI63rdnkKRwvd+4o
//O7bc3Ol+IRejMcT2Hw6Be2qVvlTQc5VLRzVnwNIPoV2kD+G/HU6fyaco5wVuiV
1u17lUhW6CAGOxmUR+cBbHhZq9whrq4+RgWMroLK4/a/YoOdjciCI5xcHNVXW8+J
ySMp+tboUluHCiyKSiHlnGeqyzsgziF811Kx9Ti3vcnDstUi94e3+gF5FRjtMM6Q
vrrK8mTpJ6MXtxwlWIbQLGage96R4X6grvGp/GTVpdG9udhNIN/v7FhSzYCexjnW
wQyrdpHy3l43h2BIvqG1KWMQ0Ohrv+2NSlVXOZf4AKGv5Hld+Un4Ew65Qg0/000s
JwjSWYRTaFGDyPxQitvacNI1AMKxJc+w2pAs8+5tQHa0AOysQOboAy1HXnExoClv
0YkoGOuMjzUOcLfkwJwpidg+mSQg02KNqBxvZOcAX5owsXNov0rZhRCkhfnLo54G
Otm2suv5xEgicyclAmGsMdgTqtHT29PLTVMMKKSCn9L60xnWuOSTWC/yFUIob0Wr
G4o3q3b+SqZs+qjj0HB01P4KXUayT1Ht9QfqDMi1NItf2Ts6XxtdkVwIuNHx92tE
TJyZNghB7+HHzrF0VJfeuyv8I9fwfhZg7JOvy6y/lsNB1IHHCAtc4opTHSZVBMR6
BGgCV5GAJEOw/EURuo5xWjqTX1JHMMdGO+5pjWQ6K87tw5XzKnzN6r5dO/xpMIjX
1ww3jmQuPhXLlL/r4NQ0aHZR53brMAsuckw2hRxokSX57nOGmLO0ZbIrkNxTkAOG
7hxod6smkl6ITJHq0LWw2B9PaLdaYa+vyFCwCzbRrn6r2mjyqTZsyE0wfMIvb5iS
MEI50XCXppt4CkHESAAgdABofIij936vQfFSNxxgizmKTBi9/JnjueJviWVvpiYc
zWo05jaGbRL0ynBqlKwyjqa3tJFo5MZME4MOtbuKnC8RcdY7y6eKSC8N6BJWFau0
pIRHxqos7LY+3uGQ0w9EmWFRpUBexaU5h5uOzXMH/tfweOSV9yX1D1DU46wUZw0Z
PKN3V+ZNUc9U/36Wsan/9Vj37B9lZdZABY0unr7+6x1eUuWN/niS1ZAhXw+adz5b
TiwykVhSCdksCaNl0F1+Vl/9p9oU89L3p9XR0GDNTURtn+f201mAPeUEbg3KfEcK
qwtaxDbkRW0yM3xSjZPdA/1ILqdDxHlSizB6r9QvpY6W4nfNUVL4/DAr2gjp5qNq
w9bsUCnGHuSJtrIsp062QOMCUTZ/SGIqSP2eZeMcOmBIaSBJogpUWdYKn8Yfhug7
CE7hw4sF1K1J/3xCmxE3o68dQLAXDSpiVYD2StLjawmVrOv3/GHUs6WEo3Wko6s3
3LYqzQvEY2TnqAaqK/N7vH+HbqSKBXeOlLgl/IDXDFE5bsZf73QxP1+/ajgxq4Lo
aiTZrYClK5iWOi9uKdIT+8nCpND4t456bjnlNX1DlECU4fL/TLfIIFjucAtMmXcu
b/wL/HDZj7+sgLl+h9QmGNZR9hje42Qp6RIfGyR0b2TEX8rbx8x62EZ5InHy2D1p
gaZlI6yMNRu0L+OPeQTmYZbpdtUkaeyd/F4akrCaGloMkRbi3gkYDy/xesxfkyuD
G8CzdAEAInVUrALA3WuIncgcN7KJgVJS5qnlp3DvIOMUgkMz0XeKESCb/uxuATbj
dH9rjZbNc3W+YsWqNqEokgoUnFSVQeNupvc/6RtttVvknAa/oJoqwLDH2N0xna8N
6RnP7nFBG2DBLKV5PZnX3gUk2UVAGolQY8wKIp5uhfNZBOOK2CM28V7SsWKcAqy3
ClagosQmoK3nTzzrPyUWex542fX3AmPeYqTU//yJCxCtpzx2ke//x5UvtKmYnI7J
X+U1AJespTloxi6mBHPUgEBALW5nbBNg1KmF9bluu0dFzOcv/56lZKvK6C3Wb/AL
b2DsvDnnOIBRy4Hk2IffyO9mLAFjie9qCs70Aftsb2Sf2FrCxoeBrlzCvUy5QSEX
K4AGfBhza5NOPZwek6zHFMYjjRarSoL2zu4RmzU1UhcFwiHqcVaSa2cD2TVQgBTy
PYXjNJ1P/yxO6uNN8yn3ExuWW/KZNEo0KnB/Vn23+rbtpMs04MS0KiRoDenqah4R
PofAyQZmk0nzdA7Q8MnelfbAbtXERIJ6da33MnL3z1sgo+IMKKmAKLB4GFGz5PBy
OWYEXkLDIkY4rF+8uiVm2R4Y84uhZm+YwYC61ItnZ9kccsBFeRz2Fd94K1wb6uZb
I920ULQslpzXS071PKhNg+FHBv53LfudSfp4/+mLshoQq5v9R/blCw5djDuwsduS
Wo/U8fSLP6Bc08cZR5gEoogu4Ogzd9M4E/5HI2tsdTMy58df+cYrxa0FIn0hT5Kk
iYRAA/i+FfCtQNm2DW9RXmncqxFvlPOBtE0j3f/Q5HDqIdOxuRxLJRrDQjZLhmLV
os1mqh4SK3B3LnCAxXroIl5UrrBK9qYzruHChHnKryQAOTTFl2mX75IX9D1SecS8
Om82pB1F5vnFb1G+nWFNgtnLR8IKckL9/TYbM+bo0MqK+ezcY/6Lye1dg+UiPC2Q
MatjUoFCkj5UZZXp5KjrStuu9P8hoVP5XCgh1BYtY1Im5L0tpe2rFDVSSkit9A9N
U5EsB3Ty2xwmNgWO79H5dZa3fTnVR7aOXhp1HSWA9L6b2hnzbFjhDSgmzWd8TxL9
9WCxRomSxcEsc52npDGlQOOsFmByYMuWG9qxveAkTd2BN4UCrbJYb5gUy6x3VVbC
J9BvH0Uigyj0+zMAkBV5R4jPVEqkHLrAMoRp/7X1CK+rD7jEME9LntwmgfSHIkZr
pEu1Kwd2WUdUizgjaxbSht+BWtqisTiBoHTmUdzGSSr+FhS7C/h1MXK5ElAHmmsg
vh8FCaieWV6ccn36fvDGv/vGt9CCdfK3W2xZ9E+iChYdo4yJSe4xm+W5/fABTDMx
XSuuMhH4fBWUYjyrqIUcE3Lznw5QchFaxIcBzkgk+8P2cnxkyudMS8H8kJ9YTNZI
L7xUoLXnkWkyPu4Dg2/X3CXqLiYz6R1H2HRGsKPB9Ii9hdSftz7ljpIpguhj1CJ1
6xIEOhTwZiWVFvNW7y/+q4gt3mtddAF2h3rvk0YMEYDzyPPqEqd6IeJ7VZm73pT6
2ziUBJ5MM/Pni9fzqTjFtBwe3eA65dJPoWgsXZkWejTdty1B+bxeqhJKr7fhLv1l
y3sd+ECv2HZGTANZRv6CZrMDqU0gN8eaWW7PNUuMRKSuXuoI6uAX/XqWiM4gyKFt
wzPs0IZmDNVoqUkO7BWb95BiO//VmL1pgs4pz9rsMVzkgM+i6Ow5zCC30HMb0Xsc
tyf/A7JK5EjzfLtPDCpzsXoWXFxMFMp1MnUksc//FlTvbO4i6JDr6GrBk60iSZQk
gYsqMn6gdyzDEeWHKa3/MTpM9bSjtdNyeoY0rabWXIOlxVyvVNpogTUgVbnwKz9K
AbGQpk6TSrlzD8CtCCxePVneuHn17fTJmO9IxxCK0oPNAfgcJMrQA9I3KPRwznVw
KuK1RERQ/OHuOheKSDmNjhYVPqYHe0L6AfpPRU/LPqKhAZwTUOmvuUIKXE4Q+YLD
ZdZ1sg8JwubrtTY3NseHSobf3mebg4E22LSaYX/BfPsP7ctKBsSc96m6jUILYdiD
gMNfN02Kqi+BQEuFSlMTTHg+Eho7PMtTdVI2W7KlBZxPw3GRGxVRex1nHcQOot3F
vGJdjElNg5uuHiRnXqTs4/6jqdUn2FBSkUtuYChT17M5/BMfRn+816MbJ7ZTdzVK
1uTUOttZ7/SDxvnuB0/r91Yr2OgiQ9UafBcPqMGmMipBVGsvqf87KdZrouEYmbKm
FB6xnOsgZOyBRWV4AnTuLOecqDTWpCaIsGygf0/9I9RYRenosnccAszYOwTyIfAZ
8JbIzPcYDfYs02oBv5X3/kiegpqQM3lIgJEIukl24YS2fDl8Twls5vxo8FbHM8TI
4DWIzcvjPSQ4vn4+YlL9+kiAlCO8N9LQx6XitjTVlYvK7qCa3VgEGZnTiJIGzsf3
mW1AtgmAIlpbWIX+yRqJ25ajSGidnH7ZvV+kQdAvsgY3EdR1bod6evaFNFLpq133
eKlYyKZpceypk0B+NA+5oZvTPXn9PwCNdr+LMarJ43cjLcPfFUONuwhXDOg+vtm2
S0BYbDeJCCUzX66+7ienFY94SrSjV+Zejc6mXTiMXXrRtEtef94b4t1n0ye359l+
24HwsZfJcyPp2Lhk0GgDH8+hYj48m32Clz6YkDy5JFe9wP6Qo9h1hG+pPT+AeiXr
wECdZ92PKQlUGzMKXfvdQzGEb2v5oRsL+3u4t4QrTMwbaEyLxwn2M47tRpWm+2wo
a8N1QVmMSkzrmvHJ14iRGaOObb8HQSnhtBmNhmSe721g+6YNcGrc6S4Zsac/0qsN
4zbPCrzR5+SKefxp9Y5z3mdDGwZRwM+gzP+otDuGozXJDo3N/YvJtIERC5f7CFxz
dxbqqgMUztE0OBByZ6qNO1QRJZ0ANtSMnyu4GjfWOSVqe/89OoMakJswlB3VakhF
XT0YB/WeU7h6can4P4VjKZxLLebolgGxgKLL/bhQn7wiObiQDgUbrnP1r/qE8vEN
zCCAzCyxU4tIkP2ISnb2SeOoP6KVl8VhjtYsxyAip3Bup/qY4DIPtABQfzY3vpVE
OKRwrS/Kuhrzdvy1TFq6WHf25P+FJiQ7l58YUHIjNHdtHd6S65k5F0ZhqG0+UeW0
27uqxL2+ribe3XKTaZ5bq8kSiMcAtDrPovNuqgoPWbfvTWXDxmPF8RkLMr7joAmp
zEnStHxVY2infGZxZsX7hlwbOlHCRTcNJsUnYCFUfI5RzqAcnD2aZtQ32x/hsgvy
7u8qea5Sgz9NMMnpBcAYK1JYcZHClXC9IDmrXyxq2FVCGVHXXbfbbEKgrAqzKXkd
I1Mw2/1uHT1vHLBa7kLdAlqdnLxaWKY4jvN8Ax/FA2sGFOTHQVAecMytivpS1MJR
JqS6zxD8Nw2rzlI0UPR7eGGA9sZAfcoIX+S4eH2z0t0YRJ/M9Lps/wXCcHQ+++kZ
nFpJ7D0TTf97Jsei6F78PgMA6kr9JFly7FofFcdIt+cN9XpKNMlT4iu1y9vJl8JB
aIlTBmgWe4zUlthFaejv/gWw5GbrfaAzX+u2HfQN905U+10OhfW9REheavI3g1Dt
7FA2yqLBB/cDr9YUMBGwCgNUmi0y4Hp7fZcou0WXubBRYKYs2x5ZyA2f+AS85sHd
8ctEOBxrvlABjKZjSJMpFXnpxgPb61X2hVoCDmpMWVTCenu0FFYiBr0IGYnoQR0/
76N8yBoWhW8oyyY2YINlB7sHW2bOF9XMcPQF1XY4zVfIgq+2S1yuDSPHUmChCS9X
TPpG82z83Ql3EEFS4WESrvGoq6cn6mWpgvpS+vxLBJnl8whtMtEEqnQ+/ODKjIQx
5rz06qT0QTtDzXZ25EsWqdiR6KqYT7BKrjw8IZQObdvusQqHzRlh48y/Yb+lhCZE
wms5PshViKQ+3ldCp1uk1oRI52vmNEKwuYY/Dok1EbtZWk4QEe+vIDj+hoaPH/H6
0trH/4HwD5/BDHscbgP59AgUDxN1M4slrGr6SLaKlwqlRB9VhkuHWm4F6m2nyLkQ
RwD1k48dvzUb9cKguQzhqmJ6HkuwIZ5oICEND8tU4kov11YGLOPnuh0V3gKs2JOP
mG8zmhG1BbKj8vWHanE+gdLHn22q/QZKQcN/28snHU8EMn+ouBVvHI8HQf5fUivC
+2LBS6kazJmhkSDusC3sztc/b91AYizaF4voYVvySaCwAkW8/1k9NAQJlaDM+BZA
4xxvdTFIJzYONqdpiAt2LtyuSQ6a4tT3+0hxb96rmgdTzuQQltlxM8qhTpOeJ7+U
fkPMmTp4M2WYz3kOohn24HE3amNnpOMyyokOY7B86Of3itKjHm0dl/vz1e0gU3hW
2dWi3VbahOx3M7PijNlmFkTISGzd66xJScaFmlQHQoydZmYmZrAzJzIaQve0wx7K
4MCEQWz3vAz/qonNewC7xxhmn9r35K6YScU/zmNtv6rc+RPV0sEGsyMOA4KLEI5l
hFDMiMCjiYvcitwIerLdZN/a1JjNevBLGy2IyfVeUDjH+nyT6xyukEfVShUEbPLZ
l4OLTrMr1/Lv1graXmmkZUSudRHb37nllS5QfXVZnb24QfDoI2KqLIHh6K2+vW9G
sNOBPzGphFGUQisQgjNs+k0hHeDgLrCUc68G0+khgsZRBGT13PHCgPaIWLTLVZ32
8pa3uMx03bTLo4rn2hYv0e7GFP/seYp07TmNe9e/qHMfqNnvnAMnNgUFKt04yNcv
GRubVW49FIiD/rlInX85RFW2GWUmLA15n7AXD6V/MwjMiwYeOSJwDnQ0mceMdT7k
LccC7DiCxldYbSHsWle0tQgGoMPs2bk9JQDVdNITFDSc8vIvywjKpmyHfl5nA2Dm
XNi+4JYIa+hTe0nwUbBj0DLTHDlrfzYCxAsiYaWdu9NgeispfEm80lMa7vnnJ/Pl
VqddyWjFYT4nTbfgDy6G1bcwx7HeeTD1UNV+fjfz+8G2lcExlu15fHyiMt8jHvSK
EpG202IwmryJyHgezPoNGGjEDVOzKx9YcGOZSUnpfXTHsUjYLAds8aLg6L1YDJYv
Wh+6USa+EykQsQJGXsdXbnkormBuOPldXVcYONXpDhoa+KXJTyPnXa4og6FmbTtf
ni0sjDAkHXP+XZucKPgS9n8mATcb78Ji0W2XvcUWjHjTRCqbgJ/ZkWR/Z0zpxnK+
iJRFReQc3XW6TtSLQFIZSSg+6ZoHxFIO7mnBnw/iXtxY/wjPQAUZIn844H37f29u
AzOnuI0ZP9tGudansEwkybCvfzrQQtirXVwjg4A8m6jQA+yuK+USWNTAl48/p/AC
yu5nvVshMRPqAeaZ04X4j/B3QLk+nlXmKFsSkgh98+kxte+xTNoy5AXo4dbT6j0F
k4L2ZKRUROo4fM9ZyhwIKZlWRCXHhfJODG3Webx38DLMM8uP0yxWRcFO9+c29R5p
r+sNfRd887veH69B8GWEZknEzzU9fOO07KUMiag2nhAY3wHEr3v4wtovQRjKrp3D
BHpkJTvS2UhC1PkIPmXAx4jsXwsshSNJahgGonq6aMXOcOJ+9iSimZKYJGuTR/5S
y4SCrv0xYqp057cUV2+dPr93WEjHvyEepVtBxMbPxsCS3fUd4PnrVDnY1LEEvFWk
CYMlxAscXYu2YpMJ2Pqqcx6bGuamFu63ONaf66NAh8CzxA7qWL4B9nEY3hENwktX
YKAunJrjxKNzgNLSWc2dwXs72Ro+UTzZEExxOxhgHUcO3RuD8hQ/ipziAMjCEGSW
EiNS8ahVvoVh3sTeDmZZ5IQBO4P88s3qxcT5oTFyZoCwfx1sEZrX/eQXS3yTnjcb
xNo9V8/ql68k0Fn+2PxXYyJhzMnlUsnXosKus+fpiMhRCR37wFWJotmoza2BHPjU
Lk39N3ZJOn9QFUzLBwNRje1ECWHPoO6AsEdUZ9SkKwr2eK0AyiVQAxEZzWzEiQs/
HYr6nO7Qvts0dGKMDxMa42BgD9DQPQU52BDset8Hi8f7NDHQznVvPC5ikj4myP2+
Y1gq64XyiFSCuo6HUbBkmw3AGO7fb/2zo3JIThH57Uu6FsBmEH7DC+a7BUSLp5dJ
tjAueTLmFFqlNwdGvlI99k0obJHoXjFzBnvUr6smZkTqbiGy9fYXqTHtQ08fZrVQ
GId3pgRU9u71s2WCnQsP/m1M0kxrdXEvv1pEGK2ALa1L9R+clFPx7QodGe+l5lC0
D7tRnYTpoXixHe6CVj9Y6CAbQ1H5S3y1/JdCNDKptVZaSLlBNU3LAd92Sq8H80qM
rvLdKrCU0gRuYg/0ZFE5mMNETEvSuGKrOpDku+Oe8iMSLjb10i5mfUIslv6mWzzZ
x9GclYyXi8/4+bQTVSezg2qXuxpGKzLp01q7jBVRTacYI1HmDMvWXvmjtXRhpzsC
bdH5dNvKP7gGSDPHda/CZaOUbPT2Qiut+XvuriMs5ZayOshH5pTBXAcAxMFvm+sk
LzikVaS9QsyxqZmCnwjea95IMuAHxk7oyaK31wH6Yyn1AZnPvAN4Xgx7P8Bw+U9f
7yOlOSgc3kgNgGWbdJ4Szmv6uqdO329s+bS8d+lAnyyUr7o5rxKB7f80AfzNCwlm
JuWNUgArzm7hgbm7dZHttjpo81oPelCN8ORorFqUwqxbAUOmw6rJsvlG18zyLAb2
C5RYbT/yGt/GXikGs6tZg6pv1FcjHboFOV2e34f57CVlwcsz0Gu3QuXZ65ixVTJI
WeBB+K3ZtRFIuWF/du4oXmGKm/z2HCeVkdW/maZ5LtM9bF3DKy8EJUonhUcYUOUp
tC41lh3ZyeEjOfDnLCpFrefpzi/mF68663JrpbjAotXajZ64scqLpca9WQKWNc3p
q52EU7v2g9ZrRhQxieoGWXxHxLv88nr2Z1UYe9UqmkzJRmaAmMPldndHuhCZutNy
Kd4+OM836hOGMgm7R7RyOX9kCkDispptLwAqG51aTwA03+jvOcUM4FEDpjos7hln
3VSDGpg2ef5LEfehRsJL0dsIdyZUSdmYre4g4mW/y4yZPpbPTvzMzsz1XRW7iYXJ
KPqrwGqstc2Lf5grUrqiw2u3cGlfjD1CUozyjldKcOsmYMlFnOI48QK3xp8b4Mjq
seGZmHfVHNio70zodo4zOzk0fiSoOUZLlu4Aw3klNXyQcFpjTU0FVdzPE2AET6Ll
RqA2/tayKjxUYVaFG3L0gsGSTLogVndPvJ/LnGIwkqQzBlNVTqXjy/vNa1jRccJw
coWYugGX61yDzgJNHTvTHnAdNj5yrJyFZmhV0zf+bhUZ15xAQd7ZjhWUGI5/XjG5
25qLwDPDk6SwWriWk3trEVuPNruQ8OlAQcUqSiZaOwFZ5i67DJVKOIAjx85itTLK
nr6Uof5x5R3zg3ftuHvxYLC7YgWb/pcMS6SMEaoCrljy6MFtFbHMMELeJ0WWThIr
fYtV6prLOEdUM6LL289QbB/tboWUdsqS4poMXA/6aT/qRm1pnR1D1Y6eEYjkhnTl
oYRblIJA2764bV4vYDAphckm7v50NFfU/Itm13zz5aAUQTD3qRFEPmp3BUisrFd3
0hZxKd3/5zCnr7Oxd6VSZavc/4xyp9c5Z+p21pQ/rLFQpV0fz8ZucWdd3vFFz+tZ
Khg1jkjNibqMe18Ht86kEKqVn8S4SeV/Sq3yCyhavtlfYdbgk3wZHKGQas2KMFAu
zN5ZazYiCAaI95jVrDPEkOE0KfV6bMIVyIni7HYD82A7nreSleKwYlQAPDi8QJcv
arM/9IUXCUQQ8Sa0JsuMg3OF3ocFEAPZdBJlAZxDnWdzrtlgXMIuyzgPMISfhbsC
cm7cILSZ5ObfSu6UNju/foDrVJPMv0W6o0k/UWc6W5UoI0+kr0sadWlSasGjKdi6
9EFEa4Su0o3cesB9sK2VQfMr5efyqQNAPEGWrB1eV/9HlFaj5U8JKezVYL8d/ndV
PPxOtqd57WmQc+0dLLmECSoFgMUAOIkdVgrMDOq0aS1tK1RoXfJFOIk9hBIEJsyv
fgQ1fS0X5IE8wU/UpHALMnF9L5AMBZiQYaDygGSPaHsYEKdr8UyZSqWnwOcrGDE/
Ky3MfmgnGdp5QaGyE/4Bs6lU/2mVYFBO+cHbgyduwA1L8pRbkU+w6h0m2XJWVXvW
mYiaQJoMKblXyka/qWtBf6rmnD+CdW65YgZ7y/OrH592M7xa8y0dmAYGFkdg4J32
89xRGhkIbk1WdKCaFr4gdXVhKu5VCctQFd76HGA4JO5LXLsbii0+Atg1+e23Bbjy
NDCKY2KzISKIT4l+v9WM/YrL1Q0bwlI2enUY6DPu3lg8ykXl68V1JFbVhLPesFYH
Xs/d5VLYu2SN7V/ddH6kmYeZr05PnsEAJ5CZjbfGPxlnofyCCGOcs9M/rf8T/ma2
GCQ3ysJHXyX8agxN3N8qV/ip4P/D1Fh2XeGRdJPBrkT+zEcmyx8WDusIg+k6z+zb
0jJJtx1IK/vynE6d4ay5383NAcdJKcy5bnQYtbPkBTJweYJF9t1K6Dv624e8Mbdm
OprembJc0oGiMSnvGc01zIwtPKJP75gG58jXrjSGnySbCMzwXh2ddavmnWUocNsY
fV1xybI5Vo0cJ5mqlSMschehR3opM7AvJEiDvXCz6x2ots0frRCkWyRpXwTnxhy4
HS3+qYnFIgOn2m7K+xCKuJ4B97TsgaauMGGiEOYDZW+dlXAGjKJ+3LFnqtsqKpid
EXR79VYiy5h5wV/JcnQl8rJ3w5bYFyWk+bd9dUO6DyOr+hsmLwTXAHDyw/3aOoEj
3TJeH6N5eSDpXqMz4dqxbtmm6JovB8NluSAoj7rDimDrTlg4+HW9qvU1BHANcQuM
Vgp7uuyXtVJRnEEDp4sX76wxZj5kSxH/bDhSgKMwsgg+bopkTIgMiYWoh5hLXCis
VVele4FiMPgYD1nflrm03ASujESTjL425jjP2zjE/+CfEXquIs67WARPVDSUvoaJ
SXmlFuTTyE476Etv48oh/bTn4xOiXIlPTlYdcR7hrHllQi5ml4Gr8NsDzn7TwNGG
sWe36nToRRPbascyS8dMJ5WgD3Exuzk2w1gXm1/ObDOJX49QsmPU/VAPWPkhvllp
ScD6Au0TpsnKPFNST/os/KUnzR/Y9gj9lon4tCGFoPFNVudAQvGGF22BMtUNw7Gh
BaKuk5o8xS15AGOPTBgQ61Qyo6KqNlaoypQSxo04rqBodbTU97yxZdWbzqvJOJ/J
OXQDok+DxkKnpRqs8O23MlLCDD+K14GgRh/7j7bvq+D/oZ0j6emTUGYJ3wZJ1GLc
9AwfeD7EcZkc6C/N4YYnIYyWvMdRdZlUFVVMbUJPQBHDMAqlqvsebLOXWJFAyKlS
lENVDBrpT0Zh3Gcp4fI85NkUzdICFs/fFEsjVN8fI8csfHg4t7O84iuhpGI7UllV
OjC/vy9FnxTZhLuByhPc2MgpnlQPLtzL736FCtVcKolhXbUTKGR5PrZH7BE+khiy
GxfjyUuod/b38wp9axAxoQC0TNopirngp7E8lwvceew2ru1HwOZmSxHvV2Uqs1er
EPvPAm1rdfNrvCcwx7R2kEWRH7soXfSleIxzybLtwqkHiI93pUYvj/rrUilqWH7Y
aLsVS/jc0cRPpCpRjnqT9plYVfeCRCSGx9zbekbvJ5wRIYOKPaMCEA4ney4zrPqG
jAxp2ReMAAwkTTTuWFznkD80PbbO4PlOVvCwa0bDUjsxcdY3O2wWYp38MdGvL/GT
Zekm16KBmey4FiRH3TJfoO/Z3XaAJcw4AhaRhI5PmEkcpCcHhsOs6sQRPGVgDQjv
sgSNA1jJhTMU/TFcfKR7cbJgSM/tc1n8f0dF06+VVN+vPXCr7B8HIDv6zfdyjCVd
BLfe9UUsRIyBK1yzO2V1gXZkUU4yTvdZ4GgVeHMh/agzHrlFGw01nRApHWDzoSou
617NC7w82g89JPKspBfxSLYwMMwMu+l4Du1rbdInulTyba5GYBhJwvCgc97/eiEi
P9uFbd57xsBJ2O5YvMV9b6M8+XSKD2ge7OgHyXxe/q+5fdLAIJ2Yb+MlS59OsYxz
+1s7ykDeS3CdzYjjwZS1772TtyFFjtMdE/k2KXmr9EBK+ymwI18iZOotyouQb55b
sbnTpMIROgKjYDyAjU4IA8udPBywQkGP6gSw7F+M7YUgJgRdwZz7eVG5q1BR+Zkt
74Bl6t41O7eiKdCxSNM/t+3eZPnuONYsJbFu0gzmExfBoJz1H3Q7+ry8/Zlyb4mV
0xODPhvf8IsLW9zWh5ggc+yE2Ah5sfcp+uAulUaX3aeRMPbqbEMduvzGfMv5mdPZ
fxlLBn6PWa+F8qRgKhsegIPUx/Mv0dpFJpIyYJMrSW9+CTECzIrumfa8aVyjcUp/
RJgEn0POd63YlqTy+2YxNonqGZAoWoXtukMrgWm4Ot+r9pbxtBjrBLazRL+m21EF
QPkEI4uB0OzGVKiGG6oNvO/ltXvszvxJfpWFbtDod7InYO5S2qpEqXxMsh4s/sGK
R1SRCKixsY9Kgg2s5JspplDG3MkjfZ/rxcOLJT1hmTMI00YpopieCNXlOHASy+zC
zx1Acfq2X+pGM2Uxzhn9RUauOcUELx/XRW2b8UQ1lXyw+zckcS/7/pt1VmHH7wt4
w0PG6LU16CjqDdQkG5SxQ97YXoitADiNWbIB0mvM1CuZ9AkYiOfBnPSjkA/9i3PU
uGvpUTFirNvq6iicIyVcW9zPziIlh5+05uhPhbFc+oQsT5E4GySXtrgbb6eh49aU
0vcPwFlANybF1ZxhmshcticJeyxRpidcJtPLXMkpLUFYl0n7tryeI2VeUgWQVhtj
EIxhmkxG0eZE23wAfWZALFhXLk26YJssNxztqaENvc4M+adDbUhBFTfy4xgz0AmZ
viZGnecIHRcICABeTfz23aAQoX8bv/TgNM9SjEQt74X+0DPDWI7TK2NT089ojldw
GSJXAHOuZSg+HYRIzQ4Mmnr5D6/cBdZhsfVl6cYX9zH+RZsBZFO4BpI7gJo3fkKl
ftel30OUzkETSihRh2/Uj5YSx/dk0fB/whcTESnImUqUGxW3KKuFt6GwVB6ONBMA
pW7dQZOCW/P68zBXOhBsndmdfcUTiAvKk2VDIJF84rns52AJ+9RGUTZCYDGKJO+s
FUgGyYFeF5h2HZnPGCdkLPmvzm6s6WCKUVV4XRURqvArSuFYcqCLNDR2duAx8Vjm
93KXpslQzZIr2cITG7gMkcZxIOf+TT7rF5oGG1W23pD607CNSLM2621TVxNCiPeL
j3StTzZm15VnQPlpehUIz9mwJdrL9hAj/uqP2Fm+4HmyoE1o+x82Eo8DIc9YbDfm
35gwlSCgh81QOlmfFXqFkuicH624xckbbW6XEYoEi979lTEOGISeapjM8oD6O0/V
ani26GADpMbQIuIInxXuVYsnscB/ggJLSP6Ax7GwSL88m1GPKDzaiiOUNTEYoIc6
PGzIqYoLkz9QVaP7D/tqWPF3sKIdbGCY2nH6ZxuD4dgk3rhwKZlLIBCRkvp00Mw8
HIXBTw6E2JG7jPjUQxt6c6XeTLch+jN18OeK4B/mNeUZSLPPPfVSVxfVAF1QRKU8
GjwOgaGota44EIcMgBM2BbD1/UOEo543/yGE7ZkbuYC4WEeRDV5lWSc68D/q5DST
uHgdcp3MrWDWd0X9gzjGvaetNRRt/8litORBhObUhcd2f4w+t3P7dm4qUjWpRENj
yosIkzoVVA1pin6SMw9wogpq2HxSiOdJwfJtLK47aIPWe4U9SukerxsEOe/0UNiQ
KmxL0yWqson+7APiDmsYLrkaYwOT33Irlw9cVw98t8KPYyuQzh6+VHu29JZEA+53
4ZcxhzWmYApOd6F5ADV5c6mngEkt//fKymWLOiA/k4W7eR5s56QW/DhMgwuRhqRT
Ri509pe+EqoFUOBs6V4ZY+wslwRZBBZyHCCrYqgVfcWRXQfBXEeNAzZ6mcQfXMRM
NOz5NokjPTd+5gfafsiT1MlU/Ghn3R7escPoGqZclaBanI4KZN8a9dvm1Sfdr/MR
koK9b+0KBG/8XpRmxWRQjNHRB/N/5gZqTwENSqnOYKk6CcB5BHge1OJ3U9gksX+C
0uKQPTL6+6uKeenwJfv43elGDTwmGsJN2d2RZtu0Tr0QiQhF6zfG7r4O6P5D8NTs
XoL3Xuzp0UVZyRoxhwkXpTcD43B4BSW3/fnqoMOF18azEeiI3MC8FHh7moIl0Xm9
WdLWZbqVjCgRX7/0kOum9DID09p9xu7J+iFCnxdnJXn++Ypx2Juno0/J0lJgQqSl
FKxGADM+3u3SUB5nfWsdMvd9ILCHhItEjMRlq4am1wxFFHpACoSvW+AydF5Q47xj
CybCW05MN5WcciPaa70QwszC3SNX89nGtceo9aibtO90TjKMTZCsXVu9HFuBBfWe
rhrK9GJJ9h4gqzB9+NHBuBU4Q8C6CC8BhiirSFU4PJbh+VAa/II3crpmfqFgjdzh
mmsBsxiCO+1qQIgy3IWjmtGce/RCDBKF+JMD2QbZiYvlMD3tOE84o1hAaoPFhhId
vOgFANNLaJUfYguH297cWSjNz28Zbi/AJNvHfnC82JOAiNjRuya0EFe/dWTUQv2S
Yg+8qcZVkOURZO3D9ukgkC3ebOppu+13x2+m1228spCKlZxt6gyRoPw2uHh854IA
M2vYULMusOyae+qtFOwOYcNfWzvxfKPJuB7dseowObdl070vFB1lungM7pM1QFSl
4xm/bBk70MpmCnILBETyCwml8cEsy5LUGwVSzsfCRE8pQV4q2LkwdvCtjb0yTvq3
eNHX3w1BF8xpZIjhgMUodB9fOdeEQvw7vtW5NrxCsf0vloWmOBhWaa13VvKAfoaS
qXdIZqGGnBH5NxjdSBBIvFTehxRf236rTIV4jI/XS15YpYQvARuJ/Q9PJ2PcN5NE
i2EFGYyvUkWmbAZb7HclXaSDgfMOSVbj8P4U/tTPiJfxaCWbH6Xqty9/sK2e6ufh
nj/DXA13w+TrMHUAthXwW7LQTnQ8FK+9/R+AIDI/p/YCIOq9KcNLLB70AGun+GUZ
2wbrvpv0oewC6AgSzdA93zSZK/zjjwPjMLdUGTNW/6a1maONdJldBtCZSlZGvE39
s1tLpAB8aB5d+HPH6ZSRMSMW9iMN/syhIS8kAeTrOnQ5ixCMd5RUnagM9Mwrvlig
FbaaTiwXOqCcKaz6OD00v6741IKQIomoLZyhyFGJpAKBPMtQoYHYO3Lc3euahv3d
eDdaPase4dG+GRfuFbN1hHsZ50gQDeCblqjLJX3RwN3PfA/kNTjXfgtg7AWJsjE0
SklBpyyIP59LVkVp55M1uL7giRLhpV5nZTobvl6lfLw4Gph/FpNgxqq1MxFWsWto
fEfEenF2FUxlTXPWGUuAJJTE71G8KiAknT9XbpAMl+Uxl+lUtFrGtQJ4R8eU2NeF
G2tsGtg/MQknMuQqR9VSRGGwpaINHruDMyydhSUsCZV56EyAA4D76WhEXgOmuecZ
+2eJxFAts9wTsCD4+FWTD9bHe5jo1THxDjl2G7qlsruU70CGO4owKq3wNUX+PA/V
KI3k12Va28uJJyRkScy0FliZxA5HOj4oXfFbjZG3maO8e0FpcPFLkVxu1gEuVU67
fDJLwqoxJWE0i4m7hneHl/wpjmKlrLKvsgT/07hQfr37q+xaPWUNJLPuz+ejmNwv
gpptyZgqMr2IBKohk09vfE15NbDBB0ETwpmob7COgcOUICahYzN3qG1vCXX7kC9q
CKdPKn6qoBl6sM909oZeZQfXpGSVfipY4xEQhRitdrfFkOyZYLWfxOyYkqE0aXzK
uK8H2NgZJ1+oNFgpx+ByuSonQW/scZWiPqr3XqhGgJWeAVv0agmiwwmA8QwXTzCs
7KBDoQ7M3L05n8Rz/I7s3ztRPdy9CPI3UKFzDN02cd1k8JsFsFzN8fCS5lWpyX4e
NzKzYQwmJOJZ07uOneKBXzDiwRdVVmJk9UJbtuDE2n65JS8Wpcc9Qvcw0y1Vwc3o
V8/v4JaS1ZmCBJTxo/nDQwqts6Qo57pO0LAlDHEs6IiSKR2geZraspgyKOua3OS7
kcP/QGxF9hlIQqvIq5q6Y7XTO7NZwSo4YD+BsAdCb9LPDPzrZlwKI9cUV4L1qp+v
d1UaxnGfw5RHO/4H2XeKhv8SyD3jY2vimbzN3aGuVnmhNytKFEivPytbAK3W/ks3
VtHljgDb6HArsJ/p4XaLbLjdBKCmugz2NnIDkr2PRedQ6ZUEBvbTUD1hl+Z657tu
kTQx8BEJ5cktliK81A7fqVK+SWzUyFRTn0a2U8sMGqyoKRfllA2/KvMvfMtrGSO/
0DjJql2orL+atCwITET/Ph10Q0gLdOFaonMVBCaOrJw8CFZSVK+nEKWoR0wJxfea
g1BIWm2Kll4m4x3g5dBOIi8BF5bPkVZlvejfZyqtKwbhTImJkjzL7W8hf7h8pQX5
fXFEGh0KjqNlkYhFnLb1MkcYjPjellRNk6HwYwD0U8MkB2I2dzrZz5I1Rw3P9eoq
iMM/LYS1DQIpyHhXSzC52y3kGN6aMuLkOabDoRrwlSwdRPwXH8RjWHBLc+tTc1gt
bfWz/4s6q20KKZLrsumWSIRzaHbUosNNwYDaLUpYR/qY3nbZXz/+40H6OfdxQUPD
1lVNR7ExHLKQpqVkhScbgGnitSNZdWTJJo3l68UJiugDB7ktPeq3CoU6GubFP+Ca
kB5jtzc2F6ir7kMjskHOa7YSrSrcopZyF439A6VXwj21a14aC2KdZtyrY0H+cQo0
WTmNlG+Fjsm8JzJfzVfdEAjI4xQ/F1p2nhYf0jfBco0JscYVgsMJV4VNsmYWFvv3
XpvWVqLKrqr4v/3FqELT/AYVkd/Icv1+TU6feI1fYrV+6gaAhD8QIlTk6Y8mpI8z
gxi+ghrOd24zbqLbI+eGe1CDbGMUnHuoFcQyGn+BlEUfat9qbNKA/NL/0GVXGT96
RsHOGa8DJWGAGolANJok5wSSNGq4/w5HvRJOkpiGSVH568urqP9HF9lQmslSsiRR
nYRJUNh/gqUiZe2bLRa/GsyP6qyHkfGC7bii8yMoHuIDygxVKpELR4JyWAw/IlIE
mYwvblYVoSE0R19AEbpfvxDciHoyIGoC7jZQotdDfvAyVwd5CHxI7c/zWbpwyq/E
IGuY5AtyGCca3BNQ9Y6hMlAw0PR2dOQ8PGo7i//a2Ic+L7Z4eQnbu2NGTfcHDRW3
32PpyNKurCfMHz72QHKpOelcA0BEQgFAF3mSMIpkSOY5MxZshOiI2llnbE4/XDIS
E9l9oT04XUTuyKnUu66sFKeAYt+WiL00sf2scgkBwCbqaj1yTff2IA6SVSMF6nbt
4kQ9Xo51u4lbwedyTriSqdSZX/Kq+zSJGaG8saord2IW1MiC/9zi1pd3+K9k99dp
SY/fiM/4Pk8FUY7Jx9mjKyiQ2q5WH76yGimgLxgqZtYKT+xtv26TUpJJ0IysBYTE
L1mX4ebVI1nNWrHZvGjzXvXL8UXxZA6aUOJgXbKntr8B5VGNPG7qBi1+FpKWoIkI
IBmV6OMvJoOnN54TB018Aep3jSRYK5Ksf4NKuWVvjAucMqxp8IIwPbpAQsG5ymjy
4KgGIxl8/jDNwZkiprijKpP64wQP1TaMTfDDsTzxHSrRCRcT8YI410oou4t8MH5S
9Y+N+9VzP9lTsXcOZM06xhVJh6RYzFwSKsB7MEbyPP8XO6lYS55YbJ7aKlH27unf
e+xXquUfF+HO9/3bUdgfJicqu8cw3G2Yx+rqE9gB5cSb3ZEmm2yjMvRU3rIQGURQ
VPwLm3GU6+6NvpJgpw900IzkHuYGKB48YnFw3r8wTGxN1YAtWYkGHhQypHfXZ+1g
Es0SFyX/41p6l2JPa436r/TPFlFZCFRnAXNur2e6Gsn7mnhr5pktn3fTpTKzpDpP
+2RuN/jMsT0Puqo3CTDJUTbqI9sl4InuQOEoOhD8pW78zIn209Nd499v1Zc/eQ97
/fbrrBuZZ7kURYQyW9UsjTZ5mXKfDrKhytgTf/pEpuWFR6LjFOT8IKfwGCDqLkVT
BgEpx+jx4W9vnHxukv2w06GFUGDoSRTLdEaBmG1CHDHcujTojxCgqEY1X7omcGaE
fbb+Vr/Ksnyvo2aaGohSBhPg31PYo+yvrsowNzSLPzilMaYA/7F9YDA3+c6Rcu0x
BXJUAdG3jyo+8GgyetPFcNH2gukQorID8uV7IQ1i3WcHmP/5sQk2cXrx7AVw0zQ7
yNFwl4qDcNVNKuYDmIMNhGERhQp53HINueaWeqZxUkIa0UKAa3T5NnkutYUGLYw0
z2sL5dm+NS9uCGLE4nQ8PS7tjaaWGBNbc6C1fX9GUa3to1rkzYCMt5LJpyKtaDZL
rSMgPddXzDboRXzNzwZ+Cd1Qemidr/osLrJaMeSFYEp32FwrX7KpzCwfK6/Guu0c
UqkdkpsNG6mIlzqFCVlgIid3Ajp6dsCpXTv9kurq3XWiOkt+tdGA+eYdx2NbJBBJ
e+uoqJhEwTxKaA+MQdl5vrjlQ/ufd060ZCJrKnVi1ChKt0pAi6kz3G4gCEpdmqvU
YfYUoV032//EJqKt8lnU6O7w+CaBqoMmDF3IOLdovo/1nLnlZaPmExVfDEaCoLvL
aXgdzflzsHGh1M3XTe2cLits9SZf9o5FZvPoSWqoQ19yvVJuNrtJdKJOPHxipa+K
lktHdaP1N03eKfGyk58Zsbew44XZx3X6BkOb4ZmWCvhkUJEFP6Yb0JXi5EDh6DDM
DyAk31l/YU5zjEzG1CUya5PuzPv7UdA7RqztRgK/b1p9K0IN/Y5IktK3Sp2TCFiD
mWb8yYm/IUEPjSlgz+/KCLtCLw86RVyIApSrwzLEU5b/nEIe+VpekAEsAOggooTG
1OmgpSYZsBIuz5lFQEh6/qOwg+tpnFftFuOFmjegUy3GqwyQVvQ4Dt6OIE3HvGHM
2FCuJQs26zkBRh4l+bhlG4w+vQV2+v4ML9gp+qQoebnf5HuD2gk67E1yChvchUya
Y74p4IjHjacqEmqkPvIFuQC71kjP1Y74yTjaQ3DTeQcoevkSszB6E+SdsofT2HX7
v5dkC9CjZQi/BqbNMQHtANKd0uzagSZrzpPmf5KHdKwO9Oa3tAkm6IJW9PPVGN7f
GhlytkOk74J7+xOvnQhrIs6zAnqaSYOaZC+lRIsV+FNMFK1stam4KWDNliBs6a30
58EAcO5oSU7C4/2J2tefCHOXI0k55aJBXcZN6Ppo7IDhb/thfToRAKjHSxOch0rC
LUmIstpdmlqliORoS895g8OzdSun6ZpKAy7DGeZtGghFe+l9fKVH9AJDXdjw48gu
sPcsvWQzfl9/ZENF+LufL4PqGM4dRArifQwYCY8+ogByTMk6czfy+p6Lcs08tdgf
K4cDvMecbpU7J5Z6siaEPRf0vIazI9tG/4+4k1pRAaMq7s4B+s6Jc/8KbNqghIBP
H+f51lWJ4hduz4fX+wSagrYUQZtKlyCrsKPEAfC+qW8v8SckUAZUtITjNzTY7SQe
P/k6GPHRQKlLDMyt6WHtQ1fUoAmMkTOyq0qRrVTnto5BT1mKw+sHKi8XQKJ3m9cW
ljwNQpWeCsppRI7ihv9jPCna+G6NGHuIrCKrrCzVKZ9kNhUQ+LGmGH7RbokZGDNv
XXvdHKeGx3mg5b9u3qUNwUs6em1dObzcLDukWF6P+Rr+2xQPUez5yUa68+91Ba1x
NS4qYq13lOHObOyuPQY7YcE/HgYmD+z70FdL7C52PTLCa6oMFiQGuZtet7hi/VNx
s0OLwNuGSIPb7Myevd05Bze9+6kU934JquSew90gLIE8bGvnhniVQcIoRHjCc4ES
yKJaCscTrCUjoei3C4BW99WlTWPizZBgke0CGYGptxa+Yy1A/ez1MnUHv0mnqjrn
9Ngok9enygWpeX7hphvMsSIdurB6N9CW6hrQQdcwt2NUZAkEAHzKZuNMQvF4femT
RGdg7r0B35Ou5Dz09y7Ihcx0RL/Z3M2mThaqzAuQS2+O9kiNUr3+OiAC9YIYZnat
5BM5krVH0yO0+ifMKlvG4QcKyq06oye6JF97gRae4Ekd0U3F7ZDZV0hi94aMq5jb
zSN81ZTu/F1qv2LohyjyjviZZcxjPWqJnyv5/AJMJvnh5iEs6sNHhvT0wHprwzhJ
qk8IyEi8ksaKvAKMHbzCuweCf4vVlCcWJ5O2bpHX//vG+SoyRsPIEKLYFPoLLk5c
DipN9APnBxdj+na4zLhOX4lakOSAhk/DZnWwrHKTmdpo/AEbby73ijQ2mDvEaMRM
AJJTrZptw/2HbHkVza2QlDjBtKxIxNMFCZNwkU8EcWJs5agL6njl6ZQ8URkzmZno
x/en2iLJi5qO8hPOqJD+YDmwRfXiMS1XA3imB+glLNQPhS+OhFLJbAqYGQEg4qll
WcgeRYBEHoqCJH4ZecBs4uYRMOL6QRcIXwSBuYXyyUl/qqXdTis0GmfG/E8+xrZQ
iOGZjwbO3ticgY3ztGag2aqZS2q1MIzWgDmmBfUWiX535lUQAKQQ+902AVlC7K3g
mzyDtZK4/WbgC4c6CjJvk42cw6DB1zOcUb/CBwTvpVizMQ4JFiLwY3c96NW1IsuQ
W1JTbUrlkEKC1E8LfbAFuDXTs0KJGNc7j1gkuMhLafpl4Vo3tV3kzEu/42w0bFf5
55odHBXS+W8xB9NRRHirnKTr2Dm2t2/3HXV487kg3WuKln/xb6Ij2uKCFVmg5BJ+
0o4altXCtfCeCFuo6dg44q058MZIWhBYukMCeh9/SHpKrQwYT6Pb8OKEeEX9ND9r
Ds2HArDoHXY1DCOep4BRGJRtcuMn0p6ZNNw2EcS6iP2YZW8o4wwND/+nni6WslKD
oOFpvvkixeCd5YVRmmxY1neBE/vP3UUnxZIA/u1KD8zlDIlLD2X9hhSSFmuOs5sx
DB83o86B7OzUKNnC5TWOICWOrHP/JsCN1YQjyKTK6/L5rf7it1UZF/nFO8a6MJA0
t8lwjkVHODOR6poJjtZwGVDusE66Vqk80b2AAJaXBR8HHabIQ8PDTZ/sgJvNEU7P
c+uS2KaOoStKA1EDTePfyfB3UtpW5FMNgTw+XRZRuyA5Pm065GiuvNBRat5qiOPH
X7Cwxq0IPTvVpCP+XAJG/eLqQLy3dzTs2+Pcq9BbfnfeMaRvvhsnM2D5jQ+w0EiK
ZflhdKR1QAiJtnHS2pcjq8pQH/yJcqXyRcDWOBIq3PJVa2RnnzQcnj8HY7eNj3Eu
+AeaFST3C9aJ96NfzGXv7BlAqwjZvDY7XZJQ2a2k3kI8lAahfKiDAz62g9gOpwAX
SUb90ig+UNyb2CJESNFAugjhDV3hEQziWK2ESbuupQbZejjF3fC9HV96YJ1rn+Bi
98laO9Wktj8zibYBGOw+q91CfQLLNQRlPq/deICt78uVXX3vz4uqB2BzzTXVdjtw
eHDEBz8sFtnhvbhw/H2JSNYlhAATTzuftbQuVFxRs0wKGQRoX0T7TFRLgMqmvS7b
4cQnQddTPh47kJUW1xnO7XflPV295qlgH67QNIyYcctKIPhEVg5QmLuBzi5nVMEX
UPmBof+HiZOWAVM0S1QfQM6HzyfjYnwxNShAkI9mk8zcqPZIFJyfsKlCBu1oO7PX
v+Ag8lKWOnNHX4qvKc8u/2q0twfiP9UYvBM2xbJZPlxyb8HKq5+D6us0tu6UWW9V
y+DjL0B/oddUTmeq/g1N9jRqLbIKoduVJmiY5Vlchb1LldJWYKcPD1rv4zhFgzrC
uPLJZ1bl19yr9/8v+NRzXXGmyscIFDaedzRLG2yBcNfi49K/gv3XyR0+owFXWpSW
Q5NlHL54wTJ7gZjxnoGdqZ9nTj/alzrMz2gJFjewOfC9yktOxb3SfGHq/SyjCpTl
1ZKgD/s4M+BMdTA1/a2QD/zf7LvoF416NHhQzAAjHWUpUFj1i/BLEbOj+Dyrqamk
oqvzZBDPLoX10T+lgvFQ9N3dIee9RIXh5fk4PNOYDvwFtPkXSJ+SRFACL6lekXbF
cqcN8sR4OZQkz3SZbwrzewKwwhKYHzibH3wfMa0sadRSiRqxA8dOuXKDgILzPwQr
bwSGFuSA5o0+M/oHqoMZhZUT1K0cuoxDa8F+kt4hPN63eWkAHx/MYyBL3wimLISz
sGarF2QnwCJ8rKgh9YaIHeQbPPn/rFnS1gmV4IXs6FSqHRquASc2kz94OFBOOKPO
YAgSAXkE/zxZb557VzfjCPL0uZydX6ZI0duVdCmsTK+UIOZLLxXu5Jjk96WuX6dF
A2s/ZV+AzO5v3+F8Rfx1BCZb8Ti3Dot1LztSnyGrQHhpsLahvSVBjh3Gvp8wu0fj
zfBSRd7HqAeFB1JE/qLh97DBiCrc+lY75LBHTDyqrF9HUyBqmIKlSxJQjhzlf6ss
fu5h8Sn2DCX2tKjiE0GTR2bHai6+E7VtGW3bgR1fRaQl6QtD5ekhdm11Fw6d+Vnb
c46+HKSFql72mrKupOX41GHSiqf8aDjxynbW8zA3Yv5W2A2fxKgri3YJrtV2LGoY
4N3R4VEm3cXo8BIuvx85OPulHz/VEhgDLmA5vuK2sfaN6+EroclSGW1zuFExmS1C
qQsx+GDUfLqSlTI7NFTXDcLMX9ry/dqvWaO/zkzx1dpYVPjmj/FqaftCEr03FYlg
HTv8uruK5AgCwaPvfFrSP10MZZGWMh59qw/Gqs9K9T/yvOCXj7iKEfSK03vFxc4o
cL4ASooVGVGerZCevsPlYZr9ITOxCJ1tcb8deGsrivUyQu9G5MJbzPaOZyvWzKDD
li39CC6wqlFfMTdhjmrWH1k/efo9xMpDXN7ebiXlxny/U/BnTeaIwS+rm3TUnBdG
dQIRlv0NqDZOY/mrFEtVAHq2+eyzJE1mDLxpYuGaET6Zyl50ebkCwsn0ezOfFLJD
kT0jOMdqJMW3NXJ55pGHSSDfPqYkI6ZI8DtplKMv/GIXRw2Kcvuk3rXb31e1D/S8
dq9H94FiP+OAv1jtYb2BYDLyEjpOt4cyDlfuWJLTXK9gdYBjFnVEiCaqmFfSafOa
WIi9x7+ti3XWpr19b3yBxsPXeMawFQ5q2x+lb6vzNKcp9J7uRJmUJ167ikzvD2Xi
ATHPIoSGQjIXeLw3xFOiCSgsWDytgtWHsZz8FrYOZvNoqGyI9Ifxi/KEhYz0KHjo
dbfK0YTCRt0nz1PnKgxoXA/JjnBP1/+5JV2vDn1IULfLCbvDR/pzXnXvswNxJ7T5
R5jsRUo899S17srQBObr+FQhrHyM6DHPc5J2Ab9ATeYN6gInJFxn7UZMFwD42V+k
Xsl95eUMPSVczaGb6ouMJkOD3lsjBaEahAFhCM5yPZgb9emtMCUFGq0rjxnxqy3n
7Bqoy5ReYazUrm0ku+GYVpLecR6lgsdtRO3zjyYMwROmwRPCF075qD3V/R1hSyY/
xEmJsTcKF1/ggcWO/mK4pZrDeC8VfxLxteM4blvqnrLjq9l1aULHjy7IV68NSCS6
1TtimLrlFox4dMEi6Q8Eb/5fAua9DVxVbd7+kJ19MEwPLVN2IRoyKFySgUKfn5vk
6tpKkblXgb8BRq8XcSA8ioOYgqUFS1gS2W8w4918pBqO31bscIlwpsWN3A4JWDA7
Z+y41M9+SK0VqOnOeRkLxlwc9fLHGVbWRJqNN9MaWNaWP1k16Sl8s+PABK+hqX87
nV6w4JtzDgC2CMPEuhU5iBa7uDnNOrFdTv6fsjncLpYpAz374mopzOF4pz3sMkY1
ce6yqrlSaCxlsVY52gjVpAHGBztNDZi1aPSsRkHIqE2YKPHnJG23TDPfF3OZRFJg
v3M4ZZKrkd6Du0Z3UrKX/+n83Y4FyzSdLXJUwWKo4HFIeFlpK0xJ7J3l8bYGn7Xa
pGOI28o+b/mtmD70wvH5j62tQCgqR8C49k26kjcgoaZ0KdVieQeqKPsm2c0u4riA
U1SE+ZWX8/UkEWOtvU/4T93xnkviUCLT23KrdjauMeUjgdS9pNG45OwKkIqTsDWt
H9atCdEfzyVkoraXoWxQUJCz8hhaI2c1muIyKSDBf4s3LwGfV8pnRcDF+BwaDv3n
q4ho6RikIa5JajprpdRyjR3H+pn+9CUnsDYKwGNzPK2UWIysm622TJyVouNBEyDZ
10wWjIl+SliID3uPvTjqqUm0xIG53xpv75Z/2dhkjSflfTX0YjWTGTZtmr3jkzek
DP0DN9QKuuiT2cH5OPEfkT7p1MrU/I7H0Aw5M5Deay8lt5zVbZf58WpvunMDXPDC
uOP7gEHA6tcac0+9Ypf4wgbdUkfou+4kgN/TKULWjIeFqCjoIc6BmDO0S1QVmWDa
3eQpFggmGggSvK8t70JIDrUY6K2kZKH9Usm41CkM9Zja1fOajxcYrVBbmqkA0WH4
ZMrCiojbp577cebsBkyJxpsQJwrR2xdjv605c85yc6RDvOQSX3evgs1AmCS88RgK
IsNRVYgFg28nZGwc81CcfMOu+9pcJ6ERyDv5bl3MImHRz1j8CZc33Qns+mUrnNrk
lSCP2xNGCBunhr/Mjyppkk9ON79fyzh2rSNn1y8THgziAPhcJaM0EjuaETLzbTtD
hv/HfMHHr7x1B6Haf8cPBbB9aOv4ykolxgjWJVT/1ce8QQXh1rRnOABQGoRwsiH0
CvnBI1yxkprDWQXI1+w51xvQYtZ3S2NG5EeVUDkiliWm11zfQDJ2Iz4i6TJZWCUg
sEYr54/GSNfYY+UDG7mYvWjE63t4QvvFZGxYg0oQ2Pqy5uAaE6m6Iao3AyNeibtJ
AfcqhFBYCn5zpEd07REYVl9reb9CoYpewDydf3klNzMUE1j+NF6S55ZVAr3cikeD
mVjwthPoXcqQMgR/t3cSDq8opg8fvVrssxyxof+LbtaHjayOdZAIV2dR/OL97GhU
EPUQpSfnI8NfTLN38SN3SLmlW/PK2kpFLQX08SowrWZ2v0ro0W1DuO/hNOXixqRi
rD9EwE7EdRSUtCMJpO3SguQa97Ay2hMD9DqcbNnoy+4NocFhkPEN0VaCN7++Iq/w
3mK4UN2ofDRxj4GwtjzJi68vgNcmh/S2567jHCCKb8/ah40dPyCdHwXX7pgZp12P
1PwRd3zsblu9zL9Zo7hHbb6NJ+vAuFScIiHbQN/EVW5D6fY5UBrI/EEPaaMS8FDG
pcFM8rOE5TIUbhoZwSjyEaxdWOaN/I7ZhWvSjigtgUFFgbOQClgeM8p96RwECTxH
4O9/SVKkT9JZDoKxicWJfuzcCdtnyzQ3BO/TNZhe4b4T4sIFZfeN983fzklVN+L2
RPqaIUS9K1PpX6v/LcShpJwLtv6QAZif9xzEYUBhkxXVePNI31W4P677w2wctG+0
sc/Xe+4xmyJJS8ZuiTqJeaIlYgs2U+0CIjOpJtYh5zTnF6MM0tBEAk/HcZLlBjtP
/ZC2SqFlcCWxvq2KrrXWw+KAjgJeIK8s83rbbYwB1kesREy0IWs6iTykTkyRLmZJ
dq3m3f4xqOSvRmvlsYifKB96EfBGbqfI5KmQc4k8O4Jbi3byc/orn6Ml2wpG7wPo
girYxNc5df/UTSnbL6tJXhX50pZl0oWwWb+Zsr+CzkPN8BlOEU2ENkxTs991fP1u
NPPnZJgMjMP//Z+7e0wYW/5wuaKv3x+IdA0kR+3h6iLYprCPf8ipDnKjr/B5HWkE
LJgBHFr39HVMs4OPrOGpe9KTpoFnKEQYwx4PMLXLSnfy9mb24PPnbzCJoVMT8s07
jpV6RpWVID8dM/dJLrkWE9spop6U5fCPDlMRu+Nm3xu2pYEaC/xaZO2lvRoVA2la
10K/41tqDZWXOI+nsm9ZgdtRFT9KF9I6LIdhElLPMCG8EwD+plxDEookt+xHwWeC
r1cEuNAMf8mYgUXjwms38zHSDVb/h09kvkTfoJbpnIWeNFzmN8kCVsXpNaPoygmx
/Jp/fV0MDSOAFh88XxUkyHTqu3oo9FK+262tl+XTSCf6HhjUX9Ir/GzllT1dcLlI
l3geSKDwlc66hSPmm4iwVWbT4JZlOYghF8YPEzDOXPOCIlYurHd2UrVxjz1HjMfC
14Hm/BC5mjqPtzr4OgdKLFKSlwmOEzlOxIOC4dshRDdboPmp1Unx8yrmVFxeFe9M
kcQiBM6LP/Yk0MFNOPITUy39jrXDNBloZnVIz9IRhe3xb6d2GMSWcKgoP4Ak5i2J
3OblOIVLaqwTP1JaS0CcynvaFKFBBoogKltetGsF/EwrkWPRgDFs3FgQzBEaMfXK
NCay4vIo9hJjSz0gP0EcbDlzPY1no6YXiw8OcuutIbSSUsIZP/hJBIK02XCibxbQ
vDto6QLuTbjD5LTZHRbYgeFYx7CeEq2tozCedb0QwtyIt0qJDsbSyjcy+tq7nQ+3
moGtyQ7ROAt/Mn8eN21624BcLPQDN7S6ASb0JZ6TjUoAgFbHYbsEF2hOom4Vlg0v
OJb8UVsGyPeqDm9gu5BbnLLVR7OJJHsXgc+vFDYQQ024aF5fdAwGHWAIdeldjdPm
I7ceHJQcE73sDyyh3VxOiBszexVKhVy8BAFfCSXkD+A=
`pragma protect end_protected
