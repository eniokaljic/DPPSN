// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:29 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gV6MgOp4Ba76sevnrd8ZGllrzqG44cFmvcVY4dxDimgyRlx/rvStP1cnKj8l09Rm
hO0V3i9th0YNscw13lurN2ESRqZ0y1BOBvbd1Serzb7b2glkLf0cc0yLS+XJN62p
C4ILNkkJ4ukKS2BYJ6pF7QJbkVmzliVknDJVanPe5Z0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35376)
R+eGDXnbsbHHOiLfGzwYhzFecYwPvetZ1dPv35I1esjSy24KW3BYlp+ryJcVQ3SL
9TMvfqjvPehvPlTemVAZPXhCob8NT8dpmS5//mv26m4YiP5hAinzguscm+XDz2Xa
nVNVJtUKKNdsxaXiwZQT/A5pl5Tx3RVUrVxWcS/YeWf+bpeH55RnxvAH5pD33Krv
ht2NTS14zaizeCmceRBt3A5b8R2k3DMNMDr7clPPjrZw7L4yv918SflLheAiryS7
KJXpGtH/lGhFXkbNdCiBJX9FPDNa+IROH3qGZkOzb83PPWfRqm52AGC3PcwMtKzS
tH4gadYMkgzVhOn5CA9+2iPFVrRz8yaVwz/XmIOckzZgWU1eQ3Qd4j9Ugwnne8OE
vUxpSvDYGXs0ltiqoSNGpKi5o9Ka1mCAjGF2Dt4g+URmr28/wZiAytlgnVU3zelj
wbQUiWtXgdu1jZgdqE7pTfAZYdaWd1/bb89Fgl0zNK3YuPLKV23IDk2hs57AvHSm
mf3TwUinNkZFyH332fsVFBs1BevFCfDsjFd1wC8tMhmeYc3fsDCPXROKFYrWApZz
Zle+dL4yI/Fg+OpF9vb9Wklmtl2TISI2nAtH1YlPCVyFenSpx0h1u+1UW4XK7622
ghYMxMgPP7bH8cIBhd18nM/gifgCjeMmY+/sL1DVwEdLZih3S0dDbQe5v8569Woi
7lEw5qVXHvlcKGoG3grW3jPFKkmaV9uWIzjv7hwX+nuekIgAT9Gg2GsQheeOtuZh
TZ8vkIeUBQoyqwS0N/QefQpcsNj9LnBrtB1Aj73m/eGvAYdNW0XRlFYil+NM3EGT
41pY6eyEvBodqJh8N8CWjWYdeLjHjAOduKvAarh2D7G1tI6NgiM5rXBzWV+0EsLE
Iw2haGgptv7DYPvWMmdreukUVO0qwjcEbjb5N9B9jajN4i3ag3lg48ewazcIFuD+
95baUZ+cToLVQO5tvety5PvCGjOvEZ0/1WMyaLb3qdeLjSw58TIBgEeOAOYRl+NT
3AZdt3tj2Y0E7Im0XjmVFg7Cd/zFgEwgO6tpKRmAVNbHmunmgXr4bdFPOqOO41Zp
kFpcsSFHy5+rBjwA2GeST8agEmm5ZPxYJ3Mp2sdAzn/9UIJ4ESNCPBnvPWZhSGiP
qhYeZ9eg07D/LMoNFA/43G9Bw6pm0++lN6p8vp/RsR8jWD3zxcAC4irEfSyGewN8
tW0owDXsNdhuEBndk49uh4C0ZfX4HLvJsqrTUPLFAN9g5ZlcWHxZaFZpA3JY1ELW
rg/zyzrlL8P4aD9hysL2E1NNkHr1pJ8o8ZzcEfawaaZRfKaITCBNrQWOJCIrSg1b
Pp2A57/FdpsLriInjtVZfznLhat3gMQqrUtPTv03Cy2WiV07qb/Hk2758Akbw2qk
KfqxSz5poLr9FRC2KsoJqwEEIzkfbQZCboHfzpQ/KF7eyL2g4shoE38+JL6sqiPO
l9gLih+amGV9d21EwbW/DFUMXYFHSlzL2mgpO+bT8A1HBtxOyXhI68QUYFafPx1e
mzm0QfrdI52iyGcyM4dc4OMkjX91M0n0S0B68I977at6TraWOoEoyLRXSfzeG70o
XZvgRBbQo9Td9TOHqJiuO7XHDHJtBlkJjw/Ps1nsiyW5KKhUerWQTxMeQT6qBzWR
xI4mKXX8/Pik4Yoh9zcYh0QzMWrgLfF1rqOmPtWfeUpsNfb4eJECI2uF5vyFZMM7
jjkb7+proeq2wO31wVcg5+j4Lz272+G4f27k8O0y5XjQ60O5JMz7PJWUWL/Oqoo6
rMjETwyE/04HKlvxs1TpVprf+u7vTzYuN5N6rOkspZn22D7FL43s1GnsWcksmlwc
NkvjxBBi9EdF7OFhXxPfjDfvFacXEi8MvSQtoKKl65040EgDEWDN5Ym0EbU3HSnv
XaTmu4Cyh9ApyHDKWVaGSMCOamvrpxN3HGMyP5iYY326kW5HzRbwi8HGjLXfIGjj
h/0sn9r0ligTa5sVMzJye+ZU+Wfa9TnKLxYTkBh4tsDkJ67Wn29IXilfEWR06yDH
1xC2zm8qN6WlqcDAPvmExvvc/EtFGYtr6DQ/Gv21ubcucKwhpKYN6CoqQ+C5UBWR
TFNR4XOTr45+TdX/TVTMLTArS6NdG1H2C+/+Oc4IXMBsCMtEkJ292pdyasuji1Kp
8Kcx/1xvysxptgtnrRUPXYAn+Btc4zNTOfZdqjjGesR2UQY3WqMOaFpERICQx2kV
2ljOIIaTkXiFLRv7dnwfI2FICpMZtuktdMwDKfqWD6jhKuT1329Fv9iyV4Zr1PN/
/13ZOBkjEHHIarl8/jo9JhpWfcrLn7tzlpybfgUQAXA+DkHO+Zidk0RpexOClizV
z0RDAepUhGEi1Qk8vEwNRo7FGbJpSDc9sVwXkVMYWopSWJ6vc8js4c2FPFH2HN3D
pAR9yIyUCQMokZtiYfw7ZqgXVpazK89coNeN0Jrx4ylGV4XJ+rHf1yXRnuqCkYYa
eP05RAJ14nq2kaUKnVhxze7+eW1priXAQNWlHBpTUy3rX2zinIXcHlG+Y6FrOCL5
iWZXcn+hodA7wZZUlNzm7k+IoaE4LmGZXrOXgJYjG9hzGGRWQ7/ki3jZhKgj1Njm
HCmjb/fJ5xAbXfLNVNLvLBiu8t61GMOy9hCkGeutKAJOWEE944SjsM8PL+3bB51/
Eju5/uFyWAwiWF/Jl6vWKqh0mFoS6Sdlum2GGkjLyw89O33OStozcpgQOGazL8o1
I/mBscfAbGNnGyrS3KSUyuYIX8IOWXjqsWlBuXerts2b0TmUd/hGWA+GjeUM9fDP
TSBXrxPW/er8xLusuAeWtFTkTam+8kPe9svtZTvDg7xDua7oJueuT2Yp1rHqRA9W
oQpEwiITNMjA4mKsDUy6v7Dabzy9qb9PSPMWZMpwP0lpI8MpP+pthFZgyuYDYRWC
3WIWXBYvZ36pd63ZumsO//1s4QUbdq/8QPaqN8weo8FDskkCmHc0n+DL3cMgul82
66mB6g5FZk5pwKUwVR1+752ghIDOeSArBYh6bVDBq8Npf0jrIH8MAQ93nInheX0A
UhzzNhqk1BWyvIEeTUkEyUvQ4yWjZlOUKxqIce0GNHNpjnyNyLTXfpU6fsNSWec8
9irGUIi72KqZEeeqTMy2wTqsMGFyKX4vIiuWdpn8F9Uk+TLsWbeXRLwy10A/HnAU
GEY5vImY/Syb+Us7hVIvhy38dBB7xmzzDg/k6GXj1A52c85k+3Ixj9Exm4pxWuHk
T0scSepFUptH8M1cZpJNyKcsa9nPTyL+6nLSdgJ0MhIWmnleVRXWAKdZ0eugJcYT
lorUypxjMzIX6LK0B7wgLkNOzub2u2easwKoSd5n82l91d0j1P/uQGDFBhjZXKWA
f5fbwFRM1E6coVM4KmH+jYWkItSrAX02e4XoVzuIcAnhllkuJeH8dXbWyE4VOafk
4O4Dxe/eSpxuN7ItuFh5ioCaLcpKrhoxJpjpAYBe5Sq2i/4Zbhsa5/VofXZlWOAB
M0KDbMPZPSAZwzuHyUPyyrfvV4Duqy61pZd5GBxELzNkBS+tk6jkAkvX8RSEMMMM
5PwVu++N9u17PPROf+IvT2OR/+NnXBZvDe6jNvsoMiJagpVw9kwFsaCCYzCtuCdW
cdlH0/YrCiYgAcz1OYAUGaWGBvXlZCndXdv/XR0u1YP3Mej155JNqjDmigM2dUsJ
oLC/dXiiR1Yn/D95lRM6bA/Amv/G1rnD/ggEg/K3j/dUgiCkS/UkL7kRKJ4KFWeQ
VjNqlHVaboMRg4Qxp5vGuYwHtZyX0i1I4aWteepycweeSUK7NWRmP5ZRx462E/Le
/9yy5bYC5XkXuzc1NktvtMQcTBSYCs+bi99tANQsyzNDONcwosKNXS8HxDKLbDO4
nnKHJJhAScoD0MbsfyTAKJaJU0Sn2MUC+6fIJzQa/ZPba93Qn+kEP4plBNLu3xQs
ofie+z7DkIAJfSCMD0/+tOgVhG7RuYHW9o5qJJXEdO7fsCsUunaERZmkv9VofxAZ
EwA9+z3PS18Gb5+WvWVo9tCC59fEte/iLXYhSWJCUl+/ITy6W96GiudfSO7AnZbn
MqveYUGXYZNElWFO+JEEZ6hOdDNlNAt1Kn+Fe0sNZC00vlnkTkUkK66+zWhj8uKg
8CfuXOGxikLtNT5fdKHlKFzTExISAqlnHM3F04mHtFW5YBmUMBmDGmFA6norlpwA
wNHGmPMyanIZC65rsHSo2j3yzqRvLW3bup2Q8qze73u6hMZPxcjC39MB0VoGOJlh
8z8wF5gslhU9Y4x5FMiu99f9x9K1DWChpijfbyZd5LenthH8bBp2VwTAX7oTm6hg
5agmfWx3BRk3iR+RfVWJ45UiJgLvY2TYik054AEdqyfu4BjzVPvukXiyW3QqCg0n
0CkoiyN7Umz9iDZBkYafDMPqCLWXv3ctsMwLEea/pKCtcVC3OTVbJflMqK7ClTlj
1B+Hzm0ylE7+4/6sWC1aPUv0zPBde3h5VlGk9p8hszdBDe5F4hYIckfD33JA+2bI
UUmb+gI+w1oL0fokRCg6Gcc6SCPHeDPYvbCfokwCb0o9eOhlEcF9iREXg42+/9R2
PeoXtZM1wvV0kUmjFzHB7MsKWxO0XVI0okO3xk1t77vK5ypVqrq0lj/jd7OkbGN4
J9D1JjCRbwETNYGWyDDpz44kasSNN0yKadmE4scXwwpSXUttLWZUcaEFg/XUhSN5
n9DGmf1bVyU49Bov4dtuzGONFI/l23miVST+f9blDaN5bcnShvPHLdICTBmTNnLU
3njSmJdS1UedMj2pdR12pLAtdpNBykcrQcS64lWEyT2iHeCCWhykbNDVpac9vWtf
Na1VampQxR0RetRdV4yIsvrtF9n9IUat/x80JckRfCMzekIfQKWeBKiYHRLJoWF6
IVm4ziEfKYQccf8LgLIjL/i1iU+6+PwjIpoytJsSamW+H2W25R8O2yX7YpqTRtm+
iTeAmNvbhNSB4Cj1h85gThofkHhAooYH+mRJkG1dl0AisC+7tvzhOTLj7rDlfvxa
pZ8w3vTGVoV+aViw7/1V86YZxqldnTH6hOqoAuKDuR3btmvGJJhDRZcNw1mAx9V4
fD7zVyXHLozQ/ryNmkVqP7C58AxgOOy6JPrwGz8HZgkNirkBRU6Ps975hlXTXAom
ui09oy7vMeiMUb9FHd1+u/21kd3f9iIZju+cibTShuvIgjksEP1hAJixvUQpUIYQ
s72iVaZJLmH6QmpHQyDfwCRVjL+G16/L/K9BsEfypvAUkArdYiFAE83bCjvep0V5
IEi5WcUVUZwmGQh9PnGHWM4cuWMtOgFGunPUr/tbNlFpkti/SiDAVndga00k7TLs
Ai1lSv0efJQXGzzit0TqvdBpiYCaQYwxL7jUqJczHSQx0r1WsgXlQdhH76jeoCWN
MyXaA2hWVm2qYKT2QVEwpAQNcMWNYkV/N9FRmDEIX+G6a2irHbCYe/+fABYRwV6E
qVtsPem0s8fKXxxYWTWOtohPxbF4F+LD1vwXNNco8cW125x8QVZ/DSGpuIySZG1/
77kTYdMyDUtqo1He4jsjVGBcMrk+goaDl83AOxG33VB7Mety92K/1Jqj14Vvhp2m
4uNPhu3QjnAk0aLzlb5ZTfoBUm8RZvkWaPPxlA+DjR/FZuyyL/o+gsfH0AHWjpwV
+mrpRUKWdquIbcEK98LZSFA1z3b9NAe/rKPmxSvpMZKCr+ceU/k6t6+NpplFiaor
8t+8JWLNWoe25wQ+eTpCKtwtV7xDPirNLerTDMKk1Qdfs/cVz1fxh4b9r2KnOzJQ
MBvvYxl+onqXhi2izIsX50Yol9ycXR2UeFetSHNPcvdHnBIYxI7BEu0OX/da5WNc
9RPqDzSLJtFAsNYZth4/Z5o9bcrGLM/+34WCnD5OW55kzjZ5h0ZKHxUGWRXZWN3u
1RUEGbLSogXuuN9VojJlnjoCWpmihGAVVoZUMjt8YAaosk8+4BlnYfw1HxoP4Fos
71CbXAsL5T+xd6vt2s3hXP2aTu+WArfMcQlN+UnOA5boZiPYMwPYe6QocH3/FgUJ
KI7utqftgEQ0AcH9zKtsZj3k+c02lCvmI8M7v5CCR8xkoG+3KO/KOX0ETrbL0xAz
MHJ9PV6VXhCC8AT1Sg1jebJ003ou8l9HvvrB9obmdatPKTjgbsteNoUSRH1FCl+b
wzcc68ZaxtwtotIjrchgJyZDux8Cf0v7fTtJAQzU9IPmbkMszeyHdXgHplNe3XPH
lqt3UAi7j8DEoYgCp8lwWGm5hdKOYdzG15nVwtc355ARt0p+sHQ/TjvIQD0jNgTW
aQEFcBKQQcv2hYxmm5kRs+VXssS7KuMc9sexwSiQwnoD0//G1OYwgX9zR/6jvQC2
Vk1XbH64qocF/7TGFeZ7IXqX5QSXd4dac49PMlTiFs/vLGCACGgKplY7DnMX8StJ
DTHN7XC2x705Jr0cu8Qb2ruqJHwBbMqq1TLOFItvr9/6GxwiP/mYwVxMhuO33/cc
yHXPoljvu3iLnKaCKqye0Z2tZPbvPyqYv3xF4Sp8bCVRtBU2MWEc9Vy9aedOi+sb
RvxCSCE+HVxzCzhb+DYZITKqAqZG0r68eczpBWeT9zmttPFi1s19gZPui9kY4s6C
3UF/qcinAUcNKTTBnxoEMEynzRfkgdwlsxS6nAIl5Nh8GWZNyHFYztIJKIubiW5j
nxCiR+W7r0EVK41bYnPLKkR13pj5K5/8iKUYa9Wuy6oakefWOpa8jaV7Swhgrzyl
ILMixEvdG/VsPeB1G7zF9X1zjwIOtz9bFbwrGFNegcOmN85/KauQJqFribcfvunY
SptkXC9Y8SxxBLzZZEYr7A1wnNnSKGC9k3T0TZhTBBJEiQI8FoMCIC03zANHbYbT
U9cnhN+ge+EIGvk/js8akoerVmjTcdTZH5r4KhjAYd56+Pm73Zhodl0Awc/Mp/4P
ooGpofBRL3fc5uCbjU774AO4RooxAyqYOAKrKv42n2gFI3N/YsDaecwXM1AuQxvC
+Kyk5wABIZqB02iQsjrxArgGxHB2V0Xb2g7vFNfD79VN4tBex8KH8wQY9qrSf2nz
o1to1H3vN5OXMyCJr0qgNhFHtfmZriaxqmtowiw0rfjQSoofNLnN/Q4mJKshfLEQ
RoJaYZNOwNKpvMPAjy/K1b/meZWg1raGjq1dEZ2r2kMMFqs3k5swevSbhX1QbtUr
tbzDrEAqzZbBkQg5Evh0s0aMs0GLgFjEdE0+a6ehAMg2oikdJ05XjMp9V5pWKDSD
qjH2bN4pNIGXjVNXUD8lTD89FQ5+EVjo/yNds6tVvJxyE2jfDEFK/7M6Z9rOrPts
DypCEuzmYWikLwDxzSlCLUqeKDLtqok/gxIV9VWWkc9ZK6PNucXZJ+N//kVdCVc9
373SgxyL01dgoD4R4v4XRuiIKjYT1ul7mPoIrV9T5KUgVNwn1adMiXFxS8Ad+8pG
d5TDzKHZgxWx+YTUdJB9XAJPMmWDjlI9Feb0pYnE/WBt8v1TOa2x1DPxVO4IM0nh
PQMQGSYfGi2q3ZSyoAqSm+C38l7y0IBjq0duFwSd8jAkcs1DnW+6LJqKdaa3WuL8
P/sbrZifki2+A0zA5S3x8Ns+pzhm0QU2QdWP/CQCBHIP662YimLrpt2r38V9yDkk
VQY5lmWPp1aVt01E+XCmPCeHnpJoNWkOnpaY//2mcP4YIbZA2KVp/NcEBDTQtIzm
zDxebuTWvSjLRFRJbR7ZJuRb8OzwLK4rfqqopqUC++wvRu1mxNrMUQQQTCfxxLqq
nTj4pkE80sn7Np1WV6F4ULAKszN4kXBOe9X3uHYF+EeTuv0mPbl5dNkEPwlNtAC6
7f8b7qTDSZ2c7Tpz46l7Et0K0TkO7BZijrX5jE/PtH7hs3j4LTV7Nnt8fDLe9quZ
OcMVQQulhK05TdI//SvRNs7vKxREmLvQaGZ3ToVcrX1lJ3cDyq6V4UX0UBhQcSEO
ewQJ1Svz8NFO95hbrX1xmCoDe5Pv3gjgtZE4PY8m9xTBSmxCoQIyqPBZQmrpKdgd
HU74+/cNaPNIm3Odm1fVZ1iKiJUKdYbNJ5CXycoSjNvAFJQXL+LfSviZkybBL7WV
9npeaSRDFpDhRurXAQXq68uqv6I8aj95hbjp1tt5wo5Qx88cho3ZTHptKkMoOdFM
0LLzSTtZeZPvdaGBSGvschtsAFVOMA+bBLpiaamMjodl81SxgPx/osU+r76NEn9Z
Lp2LemORIgREwPAMWdWNqw3j9tJmPPuD6QwyHPMWY57+xb83Htyy3aQSGxRUkHNX
BkUMd9IwtScj7DW/YQl4AozQVMt/fbOYKxYLbUXuDVbC38Fcfqr2PgTo72TKrVFH
JIUQRfz9YTTzMcy2Y8IxhjCzQvy+BpiNOChi5XdavIyScBDRcg3DtbcDXhYvlgQM
JxDJ/hdQ36y6lnsOhg99vI/SyAwtrXMsaw1rjisWSDpGI6pzlObMM2+KC30w2I/M
Qt3q34o4b0fIJP+9XexC4mgkY3fsFA9nihG2nvw0ZooK3kJlmxH+Yo5II9QJE2AA
HI9iFylV2ejFf85MUoAuhckM3EcBKCGMGtqGzTDdShrWHa9bixqgUXV1Hw+2R6mc
JemRzjDUg/qQj2jJz0+xWaxVpuF581iocoFY/3G6B8StywmniHBjqmNiZ3HgXlKV
yvqMFr96XfjF4EPxOXLO+y7+qYTLgt8w5oEsVLlQ7RdWlJ7ArM/G1ZjMZY53Ap4B
uEg/byNaRbtxQv/EYTsv42HzJRCpGsHdbXJXVHW0NDKh+39I1xJY1FtKjyEsG6rz
rdqYyzQU/WhccZf2M8bfjSKY7q6COGcNEIgXxOiAnw7W+p5UdgwYR60iGup9IBCx
lA8twDSmJZgooCm7XhGpPNmBaezShNPinO+9dY1xoU/GOWDYQvgLNQpmi2ZHRMgB
2iZ4Cdni75zsel2KYUYbgCOWhpsP4sJXzl2p9lAvFmYtoX/WHBUMkL6L8AOYovLu
MK6Ojq6CL+EF9vydFLt2RfMRxMNK1uJtqOb5DQAvll4yd7UWxarDF7lkTWM2w3E1
8QsOFTMrvAGc3kHxvQcgRrUidpZzzbSoYeyuv1vueG8022owM3NSJyGdNivkPvc7
D82VwPJEghOIzRFK6epS25MSMPrxGl+EJy5O1O6nX22dVJgCjSj+X41HNeaC4sQt
Ug0T5N2NmbtfAEmB2BMp7QsWlSy9L/o7h4wNY1rz1wNCneDGdplbLpDiuVZlTYgW
Y5x3gmj+gBpxyFkMiU06EHL4Rbc/MNVOs/NcQ8XTq0HOTNw1m+Ou4qfSfRPPiCxw
YSReeI2S6bbQ4RqSziIPbiRIOfDWVuCJjHOTHExXqR74jbTqmeTyasTBVVvjpDS1
+4/657dx6o/TU/uz0V11mODC/vpUGpAllCJdImQ8C8XAsl7tDEF9I75cB1j8P/qI
DTfuQyE1yPL+ANt3P5PGjyGdo0CwMClq3f9CRfOYvcYGwUR8kGex3NYqF5lXtR88
f3vEGPQjF10/p3zkGQd6vtV/AFOK7R5JOUjv21nys6moQ+R9BkNRLMoDEtFBina6
1rAA7xfuUW88WK8o6MOSpo0QerixpQrPCEA4yZpzkDs4xz4oZaeOynSPRwWl6k2v
1sYi3oV8NRy7QWTKC8Yd6uabZnH5vGgX2Ld33BeGvhzg8SDiomUscqPx77zPblyc
kP64VJVpaV7NahnT2LY3Bo/0Xtx3/Sss7K2EYi+zlcESaz3NJIveQTEqeXxUgIHK
wczEF33aNMQRBVnHH2TIXBoOMWwPWK5H9yXyGHmz7NyHEsQUu1iIAg5IOdTg+RBw
wEiPBvbqj/DntUYmOM478VyvSJoYI1FXleI4bUe47oBaBLxXJbMGMgtrUmZJKLwR
rtx0ma3kpLKOKLHuxTdTkCYpKI0RnMF72RFWI7Cyu2D/1Rw+l3Zpin7oxcRUsLj1
lKCgHb7513jdabP4alWfckjQshf4qD09kGb8y40CFl1SIV8SXwM6y1ksMIHH9+ct
QhFV1SrMuXbRuJdFhyC3XX2rpCISiP1wWoz9SR01EMBqUgFILExv2EBHAYfvzRwH
0QgrrTykcJS5CeRQ0F0G73FQrYY4KTt48eMmpktLc18TSZcRSAbkdMJICpU5O2oT
r9pgZ0ErTUVABESbOzuNc8eepUhehtjG96dyHyEKBrcocZR4j0SU/DlWy+N5hpS7
MMB+Uf3uLTvBYMcF1eB5CobiNgFXrPSrb2cATe/2oCG5kuixrh0VwVR4bZzDTz36
FPlkTbx401f+JDRngkIhgAhqScclD3T4UndWTk8jM5+MBvFxkRiDa12gDQaGPafc
VHic6iEja09vvQh4ap9ljziVOlJ/Cy9c+qY27iq/T+WrYABOyJzvs9QCsB++NVe7
agjVjKhbd0hbkJospD7slfcPmMqmrBfUpv3/4PR0JHi+LlgJPErfSx3hFYhSWM6W
qUQU6w344aN1CuzGXa00Gz1nglKMcJ6ShGMqQM1ivdQKaTQYuLUKMQrI26zZEDDA
fxxgp61cCZ32s0404ZUbZjnLhL2jQE+WWfo74buWnu3/+rpGqeMKuxoZx8BLS0Ui
VI6NpbGxNWRHX+c7kh9imzJPS8pZmkh1qqtF4DphSX8wkRGdR833jQAC9uXZOaez
OqgWQVt2lzyZgbRDN0aIXPrues7/iU/VD38xh2mn1CO6Ld4i/5CTq1r7twx4UNFH
BSrYRsX9Aj9bOaZ+mORdzXYuhldqRFLpBG+ZfzM6ldTohoLV4PrVrAgOjzrfTW+s
hAq6OdbooxmzLHE9R7CbfAkJSOIqOahnmCReffZ9lQlGx4tf1UAWM0DX17olE1H8
YImOVliA2ojzaIQ3WwYKspDNMFNRtKAqV0Z8i5xWZpqZoyyWzHJZDRT6bwn89ROa
Nf8IQoE1aAROLSp0kArddJkllzvXHVRX9Vt4wom96v8fvLG2AtQz4wSPKYrVUA2P
rtmcsk7d0QAq5tBbI2UtBIcje5wXUHlxjlfAoQqMp6RG4cRA9auw98Ea3IwnkKLH
KcBziiCBxtFRm54ylZYltCgYDc5Q4GUCBSiWHpbPmnuuc+KLS4SgKiFOLUWw1qZe
Tr/0EUtodLFTO9dG96N09tj6pGpmY+SSZ2nSnwvhhxylkQd//lmVssI5qNkSdgf8
Ctk2b8PUR+1bgNO/wWWjnc9C3Z2pL4Rsz370KCFBLM9j43ikWKAIwkwb3KVgB0eY
ikCHgyqlyIWGpMTL9GAzOqc1y4Cekx47utCT/HdQPQBj622+6L1QeUY+colJ5aYI
E6zZfASe+QhulwEDYCG0kx6E7fmSoA6dYb928exQcaAiI3Eji6BBnC+RFMXn7vAk
9+BVPGdczAHP9cPKefezfa2t30whHM1DUl+luf9JCO78nJeXH6xMKfDHoBgLy+jn
NmXp7Dgu3GjnqQE5dYjpF41Y4onOQqMCTckyqe55ZU67XT+SyzmgXpK3iyk9AYXH
YxzLO9ywmkU6Df2ixwRLG+xjEXG+69p/OEts13bS+c4WTXeJ+K7d74790NNFSYdz
hhX7DE1KEYRPc1/eYyIVJB9QEdW8MYVzFhYSJk8pSI10YUbnXKOSFqx8OsG/oJoG
57G/lD1baqsxx9gKghQzLoAth1DpJG2p14a3VPSvfz+4Y/BjHY4YwFwleMnUDUfx
g3OjIuMJFciPlwKisf4JRJs3mMVBnJgMkAoTqx97Oz/GAh/Yy4ulZn4x14ThzoBU
p8C1rPJ6icr9LIfWVw9cBP4Y+pdoNSOVIg2xY6YV8pEfkHXCheCjQebkG5nWyAXG
3XUol3/YsSQujqpc0sz2LuzSo5JPZHu6LFdeomdtRFFNOd07K+vRsgV3VXqi5Or/
JmpniXt/rE/IN1HUAQX8t1gp5U1GT0FFrPLrnx+5457cQhzErXalFCmc3xdQKTXd
bfmKuTSk73R03n10x68udcUOt+0HC0eBoYeRGLX39W9lUAtYzRf5d2P92bLoyj15
dE4HcTBi1aug+apYC5KFGiQGThNUiv93MsDOU63jC5a18w0aKjZ+tRoJ2qm9mS3R
o1Yyc7VG1m81l54XEYPHl4tO2tTi7lSaqKDCfvjgHwlLnE3x80CL+r8kWWUEApP4
PO7s9byhmZlcn3rNLWtm3yP7rHT7rURwYoNnt8ssdYS/UitLw7NC2ICt97R7Aj+B
k//gPvwXc0Ewby9utTJ2vT7u9I4XbbYMWOdr3j4KCP9ka03DfwZW8rPNxEVdLU8q
i5QDd8wLxjmMt/N8RRy3Hn/G/FWk7v+QmGZvagvCZumXSXZ5tevBlYJfgRabmK2e
EQ8pCIq6GkvslntXd20+D6yYEdFSfPo1vqPttDRhQb3kIeisvE3zPFRyvr8cqkKk
0sWYPFhtdpzG3AcDFhcYyu0v32CPbJLqcM+FCOLGU6o1Ym+dGCOlU8Ku4GrSywYH
YnaJkkmU1WQFAa9YRVOIfxqy6Ua5lxHDap/uYEhJi8ZlcL41ewFQSXl2fDCq3+Xq
KW0VFApb4Fy54DLJOjigHWuj0voUY86R19fm0lq773dz/xw6uWoeANYqrz1Gme9+
4nZIZERVkLmd7mwNd9Kf37JLL0eH3iiHc39yXcc8gkvs60DrNDQ+BJKy9RDGUpIU
ShjkhFpGDxZVFVug17AKwTVzqk9pyUs3aDQoPAZADgD+IpLnkcNqMZrzueUsJU3P
FhtELTuhAcYS3OWVTgfyoNSl/BrM0LsyMscJXOO1UTWCEYiv564bS4AoOLtkjDKM
t0IE01vIgR+h6X4WQWwtAwoOm/VjJ3Ju2ftJ3uD62Gi7yPXy6ThFA6N92/N/GILp
XXX/Epe3dg/itIRWQUoHI7dpc+DRZQKzZI0ddsbdqTziaGyzbnI5Xj5nLGlNiECD
B9wvWsWa+BzuD46xnZi/7KJkBLpnbOgNKY1yIdBdmIgJrk7juq2ICyROuwFQ4aOg
SaP8JFjp12fiet9UQAaR51NtStCYZ7RTNUFS8tGeaidT6WzgRQPZ6kcdj+2ZXVQh
hnMNgI/KR4UFlzK54TMkkdUrEtTFFz16OePx0viA/VK8ja6BWfKMWmnVQylH9jcC
PuN8V9Z74cfy09BBtoWWrz2Ejq//P6r7K2o2KbbFTE/1erC3mySICuBGWnmaQARc
y1cK10e9s84/nFP/o1ch0JXBWdnIDBtCh6euIzgT9KLW5dfl5/JuiTd5XOl125De
mPD2x7Ga4SZmeWO8FpSNr3GpifvYEV3DEV0kueH826ptTAtyUGKJM7DTxZkw0ZqX
DOC2e0kEsmZCBUzDBgpfoidsdaafw5VEv7g+djeSB6/a+kMRAIftYcoBGdUWAuUq
bL+phLmAj5MAGVa1CupIskGaK0iPVzx1y0E7ccMvE1/0PDswDFbSpKrBNx32Q8ic
7MxTJEMv0RX5ouJSUx3FDaFjnO4yG/tF8nxanAUex/lTD/rzqd4UlmmwYgJsliDi
X9xA1dL3pjUS0s13QXo4uTT/o58CVlTqsM9U5a4uxqo9jJv14rkxahE6LM+TQPQE
OPHYK2xscfrHd+5m1iO+oKrbiPaEmASO75NBsWn3zhFrq8YKMr4Q7es+k2N/6UR+
xeprmo+v3x0gNVX9mT5gL7IjKrusmwegX6X4cd2Aj3xAvAMjZ0XmHjUZSNCtUPet
cgTt06i0eUgRj0ubvcpQbMQczFhH3ZFHhpuO3CqR1kPUSDfpf1GuyMeSAsxIercb
29vvCppzApp/vYEcLwlOq10/GZNlOfW8HVEoC7oQMBrAG0AQwuteTosbBX0O+ipR
d6nMaqQ0zZQ0K9VIvflPZZVHgqBaRg0Ml1CWK8GXub5iU57a817mIC703W8VDz9M
Ts87XFoe6bHOan+Rsj1Xk7Ty6faf3xHrCUnrjhXFKe2nZwPkLFyeuG77XsMJUfcp
G688663RQ7VwCnME6XopuxgNWfi8Xb9ry/m+9eG4UqJd96eKKCvE1pfAjft9OAJh
pNTp7WhKU2MYJqHT2QFbLUsLYGzrSjmPSEHHC9aODQODWQEWMmxX/gO/nDa+48h1
zphzScxRQA4V2Ko3tNiPvNbyM96JVzkSoGQtrvwQOTzCi57JE3gRT8jlIZSTS9fu
QMo1iF3h85hIYcJBlj1okIk0ghAHB5xUX4tixmquvQl/by0nYQusuJzC3Qm8GP2o
N3qPhlTLVKD1mJtgEkvwMTcAibf2RDSQp2p1GOM1yVo6JUCGSR/R1Eo9IqfJwF6f
DwoYqSzfK0qKhoFn9llVsaKkPV2dLfuLimqg+cxlX6EFlJsmO+GAwz2mTiAfHHmX
yVu8o2Zn8Ll76krwD0yABIocModwX2FHejAZHJ07YSt8F7f6Dk6DjxNHGgpBrUEy
EvnSHHXiVnijHIDYfdywGFG2j4pYHrE45dAlVTbVkm3NRSLuz1zlpri0/hlzFLqa
aExhFkMwfTanUGpjUgBdurqcP4iZgS7Y+SzDQyQfIjD0VLgUi6vB4E3+6yqWJ822
m9Z22x3Ui9YJG/rY/zWas/j7o0k/0z88Guy3WSuq2nwsSYxFXxoTu4gjFDwLF3ao
ErsUwID9STOf7W1mLy/C5FrO/9hACBIikBROKZFJ4Sgdiz107ijNSquy7SGqIarr
sTbnTm7LpHfveeU17yUnTpXiNead3ucZl33yUX5KLf36vreyOQRKiPWqTpNVVxum
JmbFAYOzlya1pd8GpRfS+jTCra5IfTp0pt33KzgaeLup1aAaezecdZS6PV6TeDyk
LhsstH2LjimomydXJpr/LD1lYdHeQfESvajx6UUE79QwKCOAMqj3Sxs2HaxpFBk6
5uOGLeilalK7V6svEAPCDydvnCjlv/d+UX2QfTEjSFluw+Hzn1M9ZTYdRkAJdeXx
SczNiFLkx46Niz1rvQNkRmCLP+LgnEtnNemwbfeWZ6KmZC6GVl/DD6lqs89hDCPX
XL5VYr0X/xTlyNQu0lOReWSObAxnxk+BW9XRb/ba2pjXu7r0a3vOtfHO1nvGbNnW
OVyHD+onPERaAzE5RvakNY3hgyOMhU/k2eMSglK3Xgj9jGVstJlV/zpSEgBdwkAo
CO3lgf7wHtabHPNO22KRuCZtfX5LA8SmoJmcigIKUq4jSipvbIonjMmlBHPNnpqv
4Ruj8/HwqRqEYcbJf7bj/vCIPOgX3r+8tl73nJEDiNKMPRUfH/VS69nb979qL7CO
1XHxrcg8teT80EZWcynjh8Esemb7jq6aJ1DbxAQKJgUx7xH1L+NHK4D7iyOFeb5N
KxDfSONs+gnu0T9cWk2AFQdJsBTKxjZ75T1yxYOGPMVsOFPpNEzfF3X204jHG02N
icjsRlZ8PmjHiFGOXPOgGf7qXmfsG9IBZNDnak//4olI+X70JMTa9bzwRA583WZw
FgJC1anhgaaINWVjVHzaedIULONBa+boUh24PWFw35Zt3/TWhReOcDO6V5uDXp+V
wAatRq9O9e9wQi8GiHOjds+EjwjumgCUu98BuwpnnOfbz+W0MBdG4LN3w7eZxPcn
GMr/Bb6YXh9AkZ3y3OHsOKfU0nS77WKwK0nXYBRybv7U744MJmoDg8SjlZzl5jEe
PvKba1XHL1nQnVy4f5htwsR4Qbsu4soSeCxBjR84Pu/SRxN9A7WzoLHG5plpo51Y
AIA06IMsMMOMHGUeLqOPh6vSfPn2y4Ap1fKIERTLp0ZdkccW8mEzeanVVGQ8RwCD
SeTf0z+D3lKnQ5vsUKeM0mdt4rEltPP2bO0Uwb9IFcycTqOm++xIhlP5TiTvUiH5
0M9uE8+D0A8NKLeod062B1GDDMyMP+e29hBz3Bu+b48COth/yXPtJQlo9tAT8n/u
QBOFVouVsz38i/h3HubPJc/FI8/G6tknuMyNfhK7j44NI/eF4d79sfaezYkE993c
iM41RIDj1Fb9jNRFElAtCs5K0EcB3YPuF9U5j9BMQM9Qv06jLzEiG9Fp8xY3ARW9
3rSKpw5szK/MFVq9JfSAuijmMzq5lOGBcZuahSSPPtFMspvsDp1Uo4kUCcJiDcbH
Z/rKpyfSjf+9kjCyX0oPzbnEzwNibEy3KiQdZzGkpNt5fW8vSOs24Drr8ENTlxzk
yqjdw/pWrmmB1piRS/QJg+fXxaBdYGkyLoBIXWRDGVXuAImG5MVXxuadn9mviv3j
LQzINqWGaqIyuEoCR7oCoYKWWhQNnePVUhGLAFvT8Jbr/Qfc+fnrlPV3dhCRKq/d
31Si3DnA/i5QVoPXzdJxafN1VJ9ZdCC0sJ01eM6pmuro9l8wEW5WSDn7fQsBB2EJ
YDj6ogwsm9PrBU+hbPJ9r/QhhbbP12UxjmKDI7czO1cLEuImAWXrbd9N8oH64awG
N0TvclXiufrbXzTxEX8I1ntlOOpKh3myTc7Grc1G55Oaf9WErMKcR0hJyskX/Yp4
t5zcxk+fH2YWp/U96synloYuCJS6wF4kA38i6E2TD6yrKmafmqJuJDFh33rI1/cC
E/nx05QLWKQY79yGgWxfU+FVvN9HOTFOFMQP7UgKpqWAd5t6aQhg03WTWGnQR2cV
LtZXmn9VnXWHIv32G2z5W1oKiXrT0TsKwZatEdZAA74MLygIcaQIv+QpYCgkszWf
STbqdSTHfBh4o6vS1JArguDEpPFGpBI1VXWHIgc0bdhT/yGINXUksFhaxEX65xL9
CV3X3h5b77vcH+sH4+wm6ZPUggH5JZaUbZIp53H0WMrAfv+kbiwy2x+9f8pfE2Hz
TL/MXTqJhqSDqC4pmaw0Md/xqOydlQBiyI5QdWZaHIoh58KC/TKRVU1bsmdDS+HR
3xw+oso/6bvp48woU+SKKLm0m7Q3il2V1h2UYJV4kAB1fpg1Fy53wi0UMzkp9P20
viCclgelZSKCwY+TBj7kO8rA+TkMV0S5w1ps6NGdilJeP8NZVj4VSeS027e2V1Ih
15FVVXPK+jy0e13gOkGa2PuxHNS7gbvK7lVX+Y/WlJw8A4wOrtbsXBYhUaTQibRv
K3c25oueY/mZgS61UOg9vs9mTvEKm5p4PCaN5XPPyVBlzBgOXgqjvT+Sov1LE4jF
+q9yTDA3VEVlp4F+/AjL2Q/XayAkBNiR/7/Jxm3K1DBiBT8tG6SY+Ecu3JRYP0KQ
WDtDQFhL2ni86Biv5KjCUYtxXRHNmA7mQv8QfiAzecdF8qblaOIT5xP4BIRmsN0h
AU0qigknYH80bPEdGJJQm34LBKkukAgZcMXU+Z0NZDkJp5y5DuwnXPf16PE7OkUU
S710NL3fS87tfHYNNAlrZD3qfeyLE0ICm8j1CtYynDWGO2xKAtG6T06rQSmYY7hp
BoeycbBaVCT/08migmvQIX8id/WUR1GEfYhextLVRVOwVuo1CTyZMPS5rV6J8qge
V37x3DwSJaot3tduetAz6/cqpRL9ldoIVFm4z/R/LLVfhhQLq7GokXRzkEpMe3aP
h/POoX3AvswrNleebhtoL51LbRMp+O1UTVF0PSF/kg9GdEJatqEMzEsRXWOCsW3x
IVDCnlPTXa3LwC9zIx4FXEX/YRiAP5wUB6jww2ZjqOZBUUHhpfvK69f23LZ7RR2c
NFsmZSW5MM2hRmEIkKJtcEH/urodgfAPy4+9pUS3LvFlHsvKd4+BTqDS46mf07/p
qn2hyjtS55GtvQi3YNMI1g1FozwHBItnO61el82GUVNf7zmKaoSd2RNb+BXD0uJx
sfRb66kdECcF/uLQXZ+jqRrgiv4sgIzU48iIRREJ1wSCaTRjKHSDRQc3ni4LoRsm
u/+CpGn1b7cfcopvdJfbcrg9IFdABqPUP4DaU7Pq9QP78piRomex5BQgIiCLTbYM
5vEQhJ4j6Psz2QKc3qChThLFFAHiZHn2Vi+FRGfazgHde6J2TUcTfW8c3XLT1n/p
JEh9IRUcS+rGbMn1RVyB3ybHEhCtpPxL/lxvTHEpy4Dqr026u95pBXm8Jo+qTpQi
R2l7hZ1w2jbrigfQmWxaNJwNql0yaCwwq3BmZicP8V1AAz2DQBWeWEuyg0mTnpl1
qUDRgu+ZYv+uQcZVRYb02s7hT5fE7vu/lxoAIvIwuU88PuiXjTbVmJzachGZCWja
OnGPiBdST7mUBMZU83Zl6QfhiMGSfvGBhUnfF8TANJ2x6MDO217HhccbAoFXl8y3
Y4dqYs6+yPxcyIk9FNAmB3/Q+mLvimUR9FSq6hv9Ue2NA5VOM4XLCN4hlLWbQ4gf
VG0fL/ETWIeA+mxoUK4xG7OImHP5DbQZp/h3stAnpibklV1aoOUMD5X8BOPwWj0P
BASxIRnTs345/Nj6jWjBekH+dNA76vNMV2ra+gfJagHNjujUXcxFYrmXRn/TnF+J
fAtwSdTNY2lWgIg/ZoiqClrQ89hVPJoAKOLWUFlMjZlAN0cKmxCpYS3M7C77/UbT
9CVaJV2afxJKh8rmxrb4b9d0a8LI2HAtSLGoIut5XRLZ3GJAwvzbIlyBcOh2/w3/
ALHFRVU52QyX+ATt6FHBSeUmTZ9rM4E0PG8Ylo9YVd2DhdLKYGKg3aksTfB8ysOv
FVLThN+TciPWara492v5GtNdpaa936I8q19mrQg+jUfRBSWDOw8qqUVff7i6c09f
mms9WbzDFXNn/uu1C3+dZBCkuuaeTqZisRX5nVTOkIxHAOtL255g/45gV13mnRWh
4jTZ7lZZcopIH+20ZxesDxYv5Ycp9I/3is2dLg733ajXmlYaJwLmGvrbHm3OL67G
Aq09UvExstqDDimbYLDpr2uiclcMuIB1TVeiPgbuplec0NZnmJTUrU+n2DW0Osh4
n064lvlUNUVUxjmk/J2jUf5Zs9ugL+sk9R1/Gh/0qA+1qMIqKlLmVHSQhUSlLHON
P5hqrv4PQYTjOqBdFVaT0PuKyioP21c2Jh2lK3J0mPfahYNGyUwU4+M62TLwCC1r
l9EAzC8mFYJzat47+VtTtvJWZQSp3D4qrFsXGnmQeDahQadDRaTsNPzEGzIEEeFD
O7YLqBs3haWxM0cX7TAjFzkx+dn/yId6OtDswzGOSaWYuqf9SHHZOw0pBwqNg1XK
OwsKHi2Uy9RjrKr2bTrut26bX6nX5ji9c+gxfpi3ZKqZ4V46SyAM6P6ATnqlJHEI
6XGtVmRZhwrPcRu7FyRKzOldD5R7UXP73X58rMKosprndfW9+25ZY3oEnWtydUpk
t8XG4gibB76fcuirjroFBnGUEKFECrUXA88B/b5OgfgtoYfc60d82N5cag7d8fJD
2lO3e11n3KCb+s1ycSlJcXXRM97oBGM+z3uflJqHDV77J4c5Wdt24sKCfjlm3SmS
+cLvogW6NQhJk9X2llswCyitT00bbkRK5UMostKO+FkXut4RtXlk1wCvO8Z0rEga
ZKPQdDwKCkcrdZtCYFTL1f+hSypuQFmmrUED/CjnS6a6R8cM9uKGlxgEET9psm5r
ubdyQcKNeIPEXBq5Cv60gs8obAPjp7xxrS/orSdvnkh3+A4EE53iVRiq+SJungsi
R+lXQfdJpQEt5RwVKIHQr5nSaELbG09AVECG4FTL+DmGhfWa1iNvIKPu8rcl5OgC
yZyi31C16ICIPvwHO1ztv69FGjmtFFVnQHHVW+miFWyJnijiDgKB+bbaZAyoRIzC
30rB8Y1vaJKYb+phj4eGubK60rMGYkuz9A3SqtsHzGKNW42zUhgwlgG9ztYgXe82
+3gj1BEacY9JCDmV0ue1sxnEisGt7CAJDVMYpHPFoV/XKsI4Eqlr71DDgaDrx/GM
CikHmoh6/A8fxD9aA9cRavTGZofczMTRlWC/WddcupdTe1kzifltOLGbcFuBi55R
rLW75LPSqrli4L51BuWdlHQTJaEfQmVb1lmUpOulJBuMAFEswEwVpM48n7BJOHeG
hS4mKra0KQxS5RR0lh0qbRGU2Y2J9m+9nAwTAUhvygzy+tGNRZdGyLyDFMyK63G1
7pU2a/VkT0e661VAwo2NmVSjErduPNZ3HB2L4kMPUP5AExQNPRDyxyZJvXnycMxv
0EjbBN7tEsd53kDDD1CM3UVCOZgS+aKuMA3cTsMHjvhAdC8H+7yHQtx4WcBhTjyn
iinS2lWiZflDOycBug8rf4yeN2LZJRnnGYZivs5u7RMqU6wL4i2lvAXq/rXhU1xs
jJfFTHWFxXHtNS7sxpm+qdF6fW2MdTpuc7Gqidx7NtfvB428W7AtNJ6HFjo6l1a0
0ymFaYHm0syQ2l6RYgEssFdgycFKPlLVW3w+CCKJu86lea/VZPxm1m9eGzvXXr7L
C7b4opoPWr8s27er03ffCPrxzw9Z0jBhiEBy91YocHNEtMKiSlIkZRHzGZ2ORcLQ
Dh7KCRuL3lz9x1B0POpRZ0HmSFincjESg3DteH40lQ+vir/aOEw1cLAhqmpprrdl
tWT/uJ+DTWHZ2GOpxoQuh6YLeQG/836UII9viyoXvQrCjM8DfQBAYgcPFpGGg3vC
xRwwN3JHfWLX0YqeDy3weGiOHMh7skh5zo/ivbjh4sgyihW5t9pNApEMdgf8Xmg8
iaIjjZxPJAPWC3VDQu4Z1uBHuYgzrfeRCCIwHWWea2+0jmIcXfLhO4SRY9arPxus
++z403HZSn8tnShbJ2905P4eAAtmhixyXhBl1o3r3PMAxi2cdSQQJ4i7QeKwiKXm
49uYnQRTpbXSGUNcDkgz3PvBWzYGH+CM07B8Wtj9SJnHv1UEtfLpadz8LTq+qMZY
JXMUCVemFMSpOoOhnmOHqSSju47nrxCXOrogaufPyf0eurzMFShjFJtXItgPcxSw
QSn75wf6MTNvXqVWV8znW+qFddBINdLqNIMwfPI2u3kzclXlMfSCNgf06E5ICodT
cuIgbl47RJmEGQdC2UklewL8XcxkuXhC6U5yX4sLFtS4WD0QCA1AzN6wwsNbjLqU
5kraBlQPP7qkjxPxWFgYmPf8we9WjjbtuFaBYjVNVyfxKv1kEVGwwOVRKoUxbQwi
/2zTXDAqdzMk17Lckeq3+oQpu+5JjAuOh0iGMP9ufdombhLm8hW6TALROo5zgNb8
XPFrxUO+lFWg5os7cVJICy5EqXNYgXI3qKj6tvIFeYYt6ufvRAhZ3LYplPaHUIub
T7Nq/AuEua3j0g9PHg5eyC+snRYULURqUX+AXYxP3vJfJDYVjgsiR2XfQeIYry4/
zSRTS4edyeJVU3EPP7iIhNyw6Lx1soBx0E2lWuKP0gPnvTb/x8p5BkGH+Gl1sa6Q
yZvjtkNhr2Tv7JkrCPXf6K175HrWrY99b8M6U9z9SE/ye2wI98ikDI6H+eYkukFP
+eJEEdy5PaDJD6qtyJOt0meZxLvAIoEeNySQzwbQr/j+UfcaJEealvgbZEulazKo
Sr7pDpZc5/eLb8kmqW2pOjtYmfOnX3vZ6QrvJMitKHW38DMDqS7X7t1MeTQhrPVx
/SP49c17/eiNjRvJwZ6jAcSEPmAtAFMY0e3w2DLBF0tWN85/K7W9ROH0vizr66Lf
D8wsB/8H2YXv7B71yZS5SOwCanTtgFWbO184k25D07W/mXxJ/fBLyKgCmloFmQvp
DRm2RrQNL7bUVymOZjv3xz2Gzs5Mq2h1rMdvCB/tuFr90U0RycbHuqyauctKB9/z
gssJr8XW5aP6oaDhZ8XwmFPQtFoyP+V7rMXtwNbn4VpxU8/HxjwHnQ1OsG3eyLFr
dx4m/U86aM03/0qukKJKRr8VLH4OEHiwMBfOgO+fmgD3Io0jb1VbmcL0zrwmTw6R
RvTDpP+cbKtGZ7cO9QtJ129UqLwARpx46WL5iISAQDcxwKpA8wqaA9Uv3Zr2K3L3
ehEixgLixveiwZ8XpRHZIt/gfTUhNewZTf58SFQX8tM5g2TNQwB82CG2Xu0dBQAy
jUF7Lgbl9upd2BIVzLso2CMxsX51hopCTyJuv6b6vOmnk9gZ/qNcGLpRqFTUbMkC
27J29Pu4RGSf5bJ9KlJ8fEFG+61QomtUmh9pOyVSD2cZCEbkchALMrhWLOcnBEU5
mKOt9JkC8BMRUpeUGUhiSwYuqUQz4pPOAw41LZn3SB5C1Wkh78jfyf0rsbk60KWd
QnMqCYMF2vSlLohaI91mfEK+MN6FUVSoD7/Kc9m45y7IIFdxWAiIKO6LXGGQ3aJi
ybkPAdINOv/eNQ9FEU9VNFDrObehd/ua1l7rRwWqvgL1nfRO4OWbwogBrp+or7W2
n731xr+qbmgmAIFh6dNeVLM9SJHTQbzREd6FRwVbkHVcHKx/ZU+ZJwOHSPHOciTc
SNk0mnloy5lMcSgJncn1c5DIVJjY0E06SE8C+4aUwR1BrLbqJPwYcrbWU77aIMFe
alo5CZs+7purNiIyHgRK0i5K4o4zhgzdyxtXPuIYN+egMG+WUaYOsFz1bRvEB2Ao
RYXtjmdI0QzgXBn0wql9dbtkCOk1HptHbA6cHKIvKzj+YinOvUVj9CwYAwm15VHv
+Lr7kjte8/3vDNIkN8GeEMp3wcUa9pwjJHs7r4OYIo7nozwRf3EqjbDNzuB4MS3j
UUhj861F/HxzSAo3VeEaiMu+5X0lYXFP0x1bZGP7TOkc6biKyMjeKDzYdmFxww0G
O29sg9WaR7YRdtp6ckp34eM3YJ/Xk7jPe1GT5HT1x1jSwQyAllt6HGOJIOolvisp
Nqb9+OApJWWwc01e+YpnK/e8yEj/+xLQK2X4RPi6Ky64sgwr82lRMMoLIuagUMFy
+thzwatyVn8NBvWUZCeOhU1YUm82LmulsfEJRv4uYHRcapse722D6fDxbETJLwRs
HnmxBayunuYzuP2C2Cul7Bogkndd0GTbgZCORmyaSD7qz365FBO3RQ2Y2svAVBt/
R+2Zc4Bw1mqJS/MCH+lXFxBGzKFqeizowIPnj9E5UIxOJVm6dwxLC98ipgtgLRgg
XXYG8Z6fWu0DQx8yWrWhbtPdzzQyCN9ZWV8LZds3CYxRw1Ry+PHa2koVGWRSwMnF
SjrCBpzXJx3Stn1c1ixapm/B+o1hshIVrK13yUYwR5r4wBOTKxu9Qhdq3rbfr1X7
fJ7Sq13K8GNA/UPhYg16f0/88RiCQFyGv1Oo+lkcawFliqZso0LF32DBHDPtePZ+
+J8DtaYXUWi01CaVBDjxVrijZIgc/fzda2NmuExG06MVDTyebBBntK8or5dEpm0N
JttO7GhcFpSmdnogXwb5sMwIlyi4I1afD/T2k1pE+eqZy+dCYqI9DAEVqcllRika
LE2hG75SYIWieKrKTJrN5RQW9NOPSXXfXuam35EOGzDN7x61HI90ZKkm7Bw7pRx+
e347lLQx20uFdZAH5nPEjUhiyUOqa2Yus1S8Ytjcui++gySyv3AIu+wonxp8oHCu
oDZF5XvwchhDtH5EvxWkZKcAEQqXFkC74xMomJgBmNg15iOAkFFvzhqMI+Kyjp9D
aG6MdkU6u2hzo5H9RackXtw9c6f1g4QLgm0+Ux2wIamH4I1gMMwyTE0gymn3qvhS
gOK5Bpc4UjSrlCorzmAw5N+8tkPVuLOtxez9md/tr3rHDwjog01iHmYRxnROmfJS
vFGg0Nf2YmGSY5hOuf8X1JDmPd29wikA44xsQAEoyDHUgh8BdCiy3HR6LiwDMoV2
IWyqCbuHwPBPTQJCSVkYcJxl3KtryuwM3fmK2EyxNLfrZwC3azU9AZp2xMi2id3l
4touG2ejyW2bweddq4PUyFOQ3GqqXYYzMkzkLZ9yAu7WbNhFWClvKEqenuJPrUJO
9cj5y4fFuOwhFmJCbRUhglXO0XkaC4cWRr2I6/A3hgq+NEITIWNFmYtEeKrGQBs9
zyuOondyjHGh1DBwukhCUGM7JB2Xm3etaENzO9AH1IzQAZwrtjOSSYlZnACy8uny
Hg9aFzzVq6eKEXNMv3UdkiCin0BVzEvphC/Yy4DkmBJZgBpW6xKv9WIITJqUCr9t
zm+pvw4RvLbC2L7WcOM6NrmQEx6114eABahR0Fruq1/5dZ0JYZ3FW4z0PSpVMTls
npMYTeyIYvhiSVn3K6vWPa3Lrwh0X+j6OW9VAATNmv3ktOKfy+/yLGyRyLYcSyGO
23nPgGie468giCakfdaACtvQvM5ZgCCRkN6kVN4sqXXIWvT0c4E4msuFwcPd1/rZ
8HmS+tX3VCOQIElizsb6Bn+27nfBj6f+Xsx2xdso5LWqFBmrBh6rVzr1B1i/M/mL
CHExtLzGitAaV0p2AnG2g8PSa1DjIDQ+8WvidGgb3My7IRLnNvHjqPG7nbS57U0o
3JAHqkC/6ik4fqqAjOh3+0wPlQVZb92f9FdtasHt3FxRtTm+MxV7IDAhqtI+gXWc
QCNdKKtCL4nfiZ4HItPE36csxSnHdVbAtMnrUag+FwJm/T051bWFbhyfKDlWLEWy
WZjwz5FkziFb/TWNKU/3R2c3aqc0xSZfNjNyyHuu5J/QOJi/ycNtNaaF1GDpu/+I
BHaIqV98wN6pMxEweRp03vjAwMR0eEuFDjuS5R2wASsCq/zs2Tg2KUKXAvbvCPzc
D+eiyw8nwJOjOVYcl7Ncc/JIFdVqnJSV56cICZHZAtlnUMDA2bd0dyA8iBzXTU0B
uB2J6SvxCrqg9nVQLFfqp648YcTwOsqF3ZrkMM70VdiX915GHuUkTL7qLOtYr/Ii
LS2RxQfIzjeiK9GJevz2z1VhTToE/avclspeu2brrZrOdRLCU+gR46fgO7ugszmo
pXJqCNy2o/HJuRYnL6g5lXs+Pi7Cq1qAY2g8Svs0aMn6KX97AL48T6AH6/vks0cK
i2fUtjA0Ql/17I08vDlrMDvAIvo5Z0U8oU/0kHJe+eOYYH+tZWkc2bG/KH3/R/od
6BroGcNgmV76ncwuTASlSbyTty+QA53PvkNrPltBzAAOA6S2FEQQ7n/dRpcWoy4m
vCSrdW9N8zWRxkZCcrKoYJwZNu8trdOq/MdlJoCR2TSR1f+XNGb6LdGL3+I9BIkd
tuIvFzQ8s0Ttm0Eg91yc3Hem2CUzGAZWDoN086KYWG5C+AqNDxoWrV88Z3YX18G6
2EECOCincnweEfmm4udgKviWVU1yXDaahvC5nMvH7v3EVhVDcEAIdzQ59iOR6FpA
blSZgstW7lkNtBulA37Mjdzrsc6Dg+TQ1MZ6HDojh2j7KHGdD0eMQuFmVlDyWPer
5sHy16Md37srqLeIO2NrDBPP+iSolAlzpXjBC7e2msN8S1kiQopvSbVeBN5bSOTc
lFMfxKYtrQ3ZHxqdcaLNxwJwqDTBjxptp0zn8opE+wt2QjprjEFlte4tJXRY0csx
6juNkVhWLQLeIlxqZG4rxERmA0TitJo+VOtg0NmN/YY/kqFa4QzWCq2g5/xkps6/
4+bsaBc3Q8DGwb6nuE75LZ89N2DPA3QGB3BXEfQhys+KwUVF2MxxfqfJi1PwDqGm
AdvMG8ttoU35obbcO4q6BVyFw50DUnWU8K3Yx8lQsUuERQtK1w7+R857tiNZxuhN
Dpj6ATyqaUoUAuIhfrSMC7OF09SU8Q0kHgQ2cEMysUeBWtkpx5h7xZpTWBNGx2Iy
/sn4YdULrSRGT02vFKa+6UooGI3FWjgmUbcO1E6/WxSRdFcK/9MScWozHEyBxT8i
g2Lf6RhIIaxJj9d+BkI/rewbcBryYv9mlTTnlv493W0iLPASOEmEn1+Grv+M0jza
Nv+mGYFcZ4c3cs73oj1vISKXwshoJeoXCkgEn+DgdSQyDWjCIrw6kROv8nZVIQ/+
c7WK1AdZ8zqTDN3q1yk/LcsTPCN3+v6gulswQh4tQApUs9U7Got3K5fT5oIfHtRb
52XQx2iyi8fUnCHwfgzi0zPeORuqbYIhNf+iAhzDS/v9FQ9iXS6XRCb56cYwcdSG
U/gAkHmWQOcFHifn/AQqtSy/j85P1RL/LY/yvTIBM6nChZC45yHQ3itVTlae8BTr
SCVkfdZXcZNz0K61NIU8ec+DXZktYug5sugWVZxa3QhuF2zo3Tt8itbN/gSD8QMa
kbVBIlvG5zJ6dIaGHu/lakv7liqLzt1N/YonJyS4SIufewBT6lCtjbReGrN6t/jj
xfieHXCcG5JmHrssK0zUtd/zN14tnHz3ZERw+xiFkPTkpIExskehUlelPAUteRe0
TeHXstyo2aWMjPjD3UqIT8x/OVGhv2TdwJPm35sT99VzHdeWIplduX7qvGRmUp2d
DkwUakvnt2UUIhP8ub7ZuUqh9/nEwhKdAzMUc1BK5pBStf6Vn7cptMAOg1UiwwnV
Ygrnr0gk63GPSsqCmmwWxkK/vOakn/tSpVFyMy8sXI8IPftj75odxbJZWnVmmFbN
mBachipLMs7l+Q5F4XqPdapMxEHEgqUdA1VQ73MPhfGE03gVDouEJvL4V2RMMGuq
4y6aQTQKnPEaRieCPyIKw+eozoMfcMwVwA4e9TbrhoC1vbbJ3SxWWmKXYDY74tF4
s3KZ2D1QWj7BzvOmAMeKpyG0lB970cVke9D7VKcNq4N9lwk6pqT1/5PuNWHVB3nj
pfCl+8N2fBbjIyWTu8ztY6at6nZ7sr+XnpMK0catHH8EiK16I6oHZSq4eqieZsC7
AqDTV0LeDjfx1Cjgus5CWgMYYXIPN05xm74wrLM3JjgWigMMykCberktlws3T/Kh
JIjNRhB+y3zrl/Kij6iDU6H701BOvbhCCe0mCfk/FmeY04e1TQWYlq466ZTUvwh1
74/wBtQu4XIdd5MKGbHyBdunjbLqQ04wbwOqPseRa98v/AeLCb+/jML0FBLzzeSd
PPKnTUO8VZCPM5yHTYTO33fUanj3vjS2QTUje9/GlkAA5KQc9BGaoUxPIT2smBS8
Ie3z54cWUePXSD+XKNHPK3EAfsV8KiTT/wwfxfixp7ijL1gf+adJn+iO6VSS1r7j
TKr0yZA0uzlWk17rU/VyrEjN0EZYR0ZPGXq1iOkD4aqKyOmqtZOsQ46kSUJMddV5
WVbvKU8zRxs4bkYVwXXfcA96ISu0MEZpbhyhu62cabTSHiG7WQLnVQ4fwOAj9FCp
jhtybmYMnuBQUeGBofe5Z6YlcBKIZIslHC9GDRmn4f8niHVueyNJLp2mP1VvtS4S
PV5SFa6sXwzzAfq5t8GplRfs62U63DOT7C1yjYO7ip69E93KDzAKDPsYW0rN7YRi
/n0k/wNdVyJKqHx+S5ByT6/zDGE2dKp1f/R31h7Ggq1L8ckYE+7hBH3lN48TwFrX
ht/T2Jo6ThYB4hXDCkrHVA9mx3eP3eL3ztX2ObcQDw1LEhZxZTGUa8lr1o04JdkT
Vh8SABjHTNXwWT6yY/smB1IHysotdAOab/2zN2QUBlYlek7mumxIwxPJMG+Um8ho
r357CR8b3TqDprRCjx7X+2wDpuwrdFjfDr++CcrBMzjGWpf+fJuZg7+aBM6Wetbb
BNcYZ06YujrgqN+5ROlfFpKyWrY6Ukd2EWknPKg2ZEySP7qq8lSW9e0YtA38YIPo
5YvNYaynFAqWAnkSsCjrZuN5SMyp3bch20eqKwnNvyLWGh3sHMXkvg5HUEh9BEkT
RHWZ/g8Ae5r7C4yQSEHiftARTKvr8nYnDhi/x+Z3fCpMSwn7cLuROmqRT5Khhpji
ZZxySY8Gjdyp3htKThDgdA0b/J6XKDEvn2q9MMiOkct3gKdvz+umi/k5PJ6IbTcW
Hv6BU+eep9cUP1NZs7a2dg6v+w9AUl9A2sBuC34qs3UkClG4ZM+79e3PNQ4CxWW3
s2ff0u7LKLpmhx62ZYydy3qG5F3gdqqe3X8sq936MH7kTfa7/sqT7Hh7YJVJX0NR
3Pq76tlZg1kVPRDA+VWUbbEXuSS417FW8V3x339PdtDuWwIJGcs/KwT87lk35/Vf
iHSFaEcbjSQDU+dOQcH8JYb1A1E/a5zjpSbDv67FBIi+4q7xqUu+1xXIHoFl3UUI
BJw7bLxdl5gHsDhAzGyp7Bb2+CaTvd6M/tOh2yP6Jn7OBFQNe5Wpvkk4LjaJ3Lcp
gdaB20otH4YrLpdy9MclFOEat/xhuKf37VJTtc/Ong1bBq3I5be1NTM/GwAXauxw
C4tFPPdbdNNbArcSu9SmAWLZJuFv1rtJY5hvS75M0Ks2jwFJ5DLWxAUadCVTj5PQ
fRZguanQHNPuj984QInDCr9zJa6HFk94HnL6pa1fT3u17Mgyi/NXalNjWVkw+Sj/
9hJ0QdPC1GqHujnjgx1eUFdDcOlGcf8RnvEPBrPNxX8eRIzjqfawd2PtVYapp/d2
BCHLj1QHLgxAhlhdjw4x8w6eNqvKpvCve2ydnlMZJfeKo3o1+dRA8leBWn3J5n/k
4JuL1HDg/ICocXtQtF9xlofTd249iF5Ri0acW7Tx5PYoMc8MH5BV2k5FVxLX+4p8
xMnUCn3uj5RTytO84nhw5+i2rHLkBz5hdkpgyCNNUO138nO3yfC0E8S/jjUO9yWV
RzTIGcPB2EGLX+VSCUdQMJlt9R+Uebd8KKSpBEfkktLYbNS247ssH0AHurJbU6bi
U7QsjTnxhfMlznvaQmg+eROYTsRKx+Jpczwbh1C+5PpGmKkzmxbTAFvD0WSmRKM8
8NXied1fYVF/8qx49LYGIYUS4TXjzs4w80WPaFJxlFnjwFnKcwhDR2Xel5cvfK4d
kN+d1PLgyL9G6RDq9YSyF0arSaBM0HP34j0kY/0rUKfAge0Z+lOYPuSRJG/CL1jo
p5vuYMZ+pd8LORZLY9DQoCq84td00xQDyOko4p1Epwv8yI3uNxWd4iDrISe9zVZO
AlBJqI+QNNaYJ6SpcziNUu6sFpT3yKcSta9D4BFz7HD7VnMV7UGrlgPgOkgnpaso
1RUaDyI0gErHOj6RcwihnU7D1pMvew09MN4jG2XSZKalhWxb2/Z5aZ2RpBrifTx6
aIQsmt94fX+JRAbKVWksW7m4Sd6pvHOD5jiUjkRBx5HR1IOOVIq37nb/KAEaC62R
37yDmAaaNtEf4t13o2GhOtmP6ug49nJA+SxNJSUe2JKb7oR2H1N60ND1SREUbhkL
XjaipmHQPEER1gVPp+nSljIuiocypR9AbeHKYUT0rQwfPIMOpJcgkFu4JuInr2ur
vg0CjMpCMtDE+nAQPUhhps/su5u0RJoI8mQezZ3eYGEfL7/MzxTtKltv8M0dJd95
oQP92NSTcYd72+cGx4YWIOvXiJTQQg3F3wKlR0o72BfPsxSHKBvxF3HmHtwsqpfN
E+wN/rOfuwBxeLfbZm1EjjZMkKEZiKcg/4PYnQqDc+wdzMzXZS6wGZZjhfdS0bw+
nOMbXwcoC+xCgpyZ/1QxiWAJK8UysgqHQPzltSQzl0Js0MC1dliSuuXsnBxtl7oH
2XXp/Rub1wL8ctfr+hUUKvgWjDzobhzroOCMyoxEp37M5/GYNSJcWgeeXuAAHE9A
Mt+5OwOhH9cJIawWMd1EURBqugvKZEONvAiPSu99KtYWRE0gmpEaRR/Hwv5k5Ia4
yqPi3HN+WVfwbXpze89xN3tcwnA1JCkMqoIXPL2loeXeMfsp6sx2qqlC3xIr4qEz
aMVqqTSbFQnImNSXi0QS7qNBjWbdIl2Q2VH/6mpvKFIuLO/tIRKEuymdNi11uDsL
PvE8iXIeur5GBtmHoGCtHEuola6VIX0wZ9qvAWU20lDDqnzhQX4nDWbnDPg5sVhu
MUeJFTSuhZv/v4c27gOXkwJuZBnAyC9JQ5MOI6va9Ecii+WRGblEqzDXxgWw0KHV
nilxcsEpp9WMvgBC+9d2j+S53XpdepmXkpPsZkk1sdjypzihT3snhq+73buOcif1
uO71ecRvTrYA7B8powejPAJ8y41F3TyY3TL9jO8j7v/H6ugp8Ztcc/RBxYtIUBo1
6UjTwt4zViS5tHKlYswkCDNeTvOzGNDhLaBMvBYN5MLdGPZB97Zj3Nr7p6Fxk8Tp
267RWZLe6C6ydgFbQuHZvavHtDFS4Xl7KIYIoLoen2v09GQsRwDRFr086DsKO0gt
blyfalUowcGlvhveBSZZvp2LItTI4UH1wBRoSdzXyrzDCYCmSTmDCb5sga+U0SLD
1c9+UidvQnnrRiZE58Ttx0AXv3uSupdzfiugxiKNGmzqCqeNBg5kwPQ64mdpTEmZ
s1kO/6Z/ZOypM0R35CVGvWQWIsv7uhk3qadwR3lLjhndT+uv2vEJ1DVzwusyG7QB
d9p+2TPBCkpa5wQytMTfdQoJkywU1ZTFUS5BCYO18nsmpofS36PpC16/S9C1OXYs
vIc5RHEJGlxiiCpUk7EbsOhREr/rMNO/sD8ra5a1sgqo9KZbNygl81dhsiASRFCj
M1qcK/UMhcJ+YS5BB8nfEkiBIH2XnLLZs3NrGwmXxFZDeH9PYGOXezxVKWMtNMw3
FIfkBnpFdsj4ggQ9HHMC7xr87qHzaUjg+y/PybMHk806Tk4PLBirdDZ3wfDnykQ8
Go5c7F4sYCJjiB+wgAzbaqegSE5nFRCeTGGnTt6f2XgiCuYS3eNMu0W6VVqaQ24f
tBYmPPaOYtKXCtee91j8N9FmeZ3LDmho5bxEpSQiFIcNLGUsDYHOjq/pAnJa8LlI
K52223qgF7vmsYo61MQ4+QlGnulvndQGpc8kyAyeRehSCJAAXKmyf1u6S8TDa95I
2L/NBAw5Nujml8o/lDl9BBs+2vgFxl/hqExhFfTKReKiVQNYCjBC2NDR5LjvtCPT
JqrGop8o5lVgDcIxtaOrq4RJzmyJHbio8L+a/0d66SucMjsR+iY1pdcTw6FdpTnr
hs0MRypsHlGVvcpranjaNApkMqsj3E2wJuo/+DN16qBjjyk5T46E1H+rqrVNMx+8
CQX4J0aN9vqTa+S9ltRRdny5UGEaKKwmdKdBTX8vyNCIAbYSDqz9vbrAvWHZWlc9
7WNbhQOMRmGIe7IeQCFg1LzHKMTjraAUR4NBAYnYi/ZOKFWpI5dxuZeY1Uu8keyT
T2bcf4WnrNyWNCX4NM2seT2Z0UxFmP8EXmQXT6A5np169NIYTqgXRSacR9HjqUzC
TGvaIsKrPOk1I0sa0+RNvhHgwcAEw0p/7jI4dFq4tsS5kJjNgDIFwc+2/i1m0azz
JC+xOUuc5wsfoLoDXOn7K0B1tGxBqz6NAzS9fuRMlt7+7qfqEri5BpbntOXljX8E
FbkxecDxggrO8laNzIduZ0+ek/KfPDffcI77rGJA6Pa4dQ6qVSxA0TkLt+nmQ7c4
Q6MVI9P+uKEt7AZ2Qjn2BFjhxndtFAITC0vrcg/P4H0X/janjLI8ZlxTHa4KstSN
QsJx69RLh26Nx+O1IzRy3+LFs737h4MAorwh+LpEemp5xHEOE/cXKRjJdVSypYY2
HjDDsv7zTYB+HpVAkUBF2pcGVGk5Bs/6QGlueP7FGASXTFS2+/cTycTvL2RfZiXL
gHee1Fpd1TLd8T/3aLziKcKHUa0Qmj9e3YNnoZTUI564BHFHZXrq0f2YDdYdNxLi
o7QO9XcNvQqK3aaelwEr9NyGiuYovvUUM+76zywNEv3uv6R41gcjtaBSiKLK66Cc
TZQ07v5Z4czdr7nowsGoHDIyJQZQaMeDAXKlZlgz/+njAIzaWGcUtG8ebKKPOUze
rqEIwtmavTCiFLeI7bB0KvcFKf7SSomgIOj+8Ue1eNbMBYPooo/43GS5ErtS5VlN
5NbRc73q24ubiFIBtelaRMHl8QbhrzwQDwItMdnEjp1qNhd578A6872GaP+sjn9l
WI8hgJxXQm8UwwsP3VeraGRrtZxyLMzA8h0qzUGy8WHHDW+vrx32RRDoYpsmnS4N
7B9HdmuTuFiYB7JoR2QRXWSAhTiBSD6hhBfNkHaWrnUzDpzU1XZ+/0MxCo93NoGj
C7X0+U4TfxLWaLqYgvcrEdk/3WVT72Mb1+2UbOgq7f6vpHhliLSpL9yL2YuL+kVz
me47eG9ziCSgPCrg6U9IP9mz/BKst6y6Ri7rNCQAiBJWYq6s4PQTBv550OqCEFGk
8XDbaStLrN9ACaJDJri+HCrJvPIVM3sWrhotPY1DpKEDdGqyxHFs/MAbl6CCxuCq
sU/LnLx3Mb7HpZaDKpBYhpGFOItaQOdpxtMAoWNl8VwAG4Iat3UkMTUKm9Vgoo3r
cLSzNbmp1IFPlba+DIFX7IQNmz3AHXOpeapdGjwO2tMYhTpmX97daPyEEnfIlHg4
Z72hR8Qj8YwvGd9N3gp8umlx2zMGwIU2LoesYahcf1e0QW+tbEYq1iVOEqqRWa9s
F4NzaTL+7n0bTJsb2nHNJRew65MYfUau8DJ6sQd/6lf+yNh2wc4awTDB6nYpUhXt
ym8/6yXfyvfRmKn/at1cgqPYrp92SwTrpW+xrU1vtQEwtiB564M9u4qZi0/YvzKh
gjP21Y4Pmweeax44P//90nw99t+KbfLr79ZPY75oMmjpwDkyza8Orr1hINqVwUgE
zALdoF1LGv4SgC8RQ0sa10iIo9JEDjOYvcxnWCfeTwj3UjBwbkrrVJTlFrsyzrsj
QqYDwO95kxsJaFEcWB1H9sW2nIC0Xaz9FS4UfPuSd8qORcifljyc9AtpYqne7CQC
cWasCIylCOe7HvAQDdtVTeHR97s+OdS89yVa/ZYvAYcQu5QIiUjJ2brQRP0/denK
Q2BbgEVEY13DdrxZ02EsI+C8U3dBP8F8jb01TeTrg5Lu0KX+ZTHdKMu5opX257dH
0qfcS18uhDr+VdIObyZ2kZZBJPg8fp1Xk+3CU4kvd9b9rPRG4yX0nW3kNRrKVj0E
ul/8Dd8GFbE5jzfgR7DynYLhP3hC5NF52PlgTLIN9eBDjzZ6LqwSjWHGasPSRksP
BQZSVcgZWWAGpQn5C8n9DZuPzm0BowTmfLkK/qlX4tfUwOaQ5348cEZ4jtBGZTaQ
CHVY6K3HQQLe08TSkIlZsAzuZuJp8+/2RslqK6q1742Jg4gKkswsgLC8f3LGDeve
YBk3iFnFOTjNEOcIik+fBkOvrwqQH7Pvo0OCDj/VXkocBviL9A8kdJJ/5qLLGFiD
EWskxm1cN64CguoOQa4qwoG6FVGFsZwFgY2fxLOjJeKMln3z4Hn2p7kl4NZXaokO
pv/dN+Gh87rSENWbv/eA0J3VdFGkcjpoDoHvNH/LUwIHZrrep2cRx9O3AfkX0tTv
dv90/KdB0wK89ucBzRiqmVhI4Z6dHapHktONQfBec7HUAVhuKNlb3aSfgCjsL9ee
u96tKgIjwf5c7YdvOdYFquAeB/uQx+a4lXFvo4nJ8pdvMkiNqqpk3EAefQgt5fJ4
mnGf2G2kbYD6eAtgerO750OPhFkMJqLr+bP8wYZo7aUvvSABOh7XzBnuFyEdZOsP
qLZ5guL4BPaIj8nAYTkueAHXddPjMgCV3rrTtE0V7Cm2LHjbMYhaV5DzmfHNepXA
JaUekWevTigzmbiB4JxyxBEUlLQE8T89qUJplwWDMXbsdufLxlHmuLXCD6sDwtWR
2Sw6VQ4/tKxCDy4eIdcsy7j6olEsl0v6U2cEOFXQ6HN+2HGcU8/S3eEyC9/oGaFK
Ml6qryCalizervl6FK1Ch+BGBSQpWjzeR739FTuP3rXexuigk7hMVdaxDrhzgQxj
C4gm9NsA47XclVvo2eRk58mAErAOeyA+Ah6iEdES3bCCB4zMZlJOdO+T7FLR74Z7
goZI4ogrP2B79oS2b3ySC1EVqJ9LETzR+FryFFcakUq9HRZg0t5KdIKU2tO+EgOT
bU3g0DjiqE3qUMbx5Tfuo2zX0+3p0zZ0omiiCnRbH+9nbnDyAo/CIGN9YriqgqYF
7e0ilak3A9nOMfprQfWBCAJrdIR7Nxl9M2rzA9EjNLSZjqVloeAZVM0CFVR5EkvA
hTmzujghO54XxfmUaXaOQPm9w6PMxyH1ySbT62XVZgLlhOUgJkQZYfObGdmAlB+S
l+sNz4U3WHr7XdBq5xep3elYR2RWcmMvE+IWFmObv6d7cFNoMdx8peZxM+gbmi85
umv/kJGb9NDgMdBoOObFMhVCOTvftGX8UbQPL+KamjyGOYkFTNixpvKpf8zIGvme
xSjRdIg2TkjByaASphynq/OU6NAmBmIe23BvWVb9buYnmrbvY2B/GKk9IDp2X+Wx
S2vpcA6ScPS2MpKwCXzShUq9V3aWfddGs7AwisBuxT3E0/a+1hcYxWYXpNjCuhBJ
Ht/VPYjpI8qdCh13qISHaRpPPFrWE7zLvZSlwN+6r5M8FICoCYUSziI+/hYbGQxZ
n5F+30+Sm4u9PCpodHWXCkN09sUG6MF+qNzoMAGNprj8a0GpIeHMl9+hSStWbdNI
x7vNvdo6cCFhhAcJ+1M3J6WqG7n8Z9zMB0SomJGB7JO8FHhnBDApCtcmSZBtvxTz
oiYOcaEvq4CRCI6KCkLZsWoXGaz2uRnA0+ZGQHLR63fXeP6+qVFppRMcQRotA+dT
4sfuZK4asNYeYxFLAAhNLWmwPCZXUsowizD95JYN0eWh3xVoLgHlW29ljc0VvoTB
bTiu7GU+dzk59Yzb0h9696gvQAuNRqbEM/6mQy/6okeh1lamGXrUcg3DPYXSymdz
tlxVqaz/fyUk8drf2g8qD/1gDm1BC9A+Y74sAnEgpHxCZiv2kMgdWoL1R04QlzGV
yb2Sagz60abIaOlzXU9pgV5N6YXu/ZWjC1xUKclDYPlt7YaGT6tM2DA/R3ZN9572
d0Ub4hR3/XgtznJTUAcGRXwkp1Aol7lrCB0yhm9LjW6ITEP5I0lES0K79lbKGC+P
fVwJtTsuM2Fj2jrjJ+zIWSQXO/HgMapiDAlHd1we1QDVqX2ljuKFsodvXCE1zKD2
cCXXOaI5TkTDV0GBEsXFU84KPzQ0zlrK3L2nI+Q5pJzww2czOZk1DbWw39r2jajE
Y7etadKgWeAYT291wpNR4vY6Wk+tUFJzNU6EVdJY2NPMpUbAIlcdTZy7pdSSQi4B
L0u9O1p7HHiw/LFXqPpVa9MgkwODofNDWn76RrZMgLKm2vK8RVb7s14A2ms1ygvt
OKBR1PP7tzpLKn3/Mu9dDPavC9T6Ij6ct0RXhBmkupn4A4fOLiMvwmJaJP+7MOiY
gIVmzCzh9SINaLzZYzU9s01IC7o12VGXkrcivPhaTLeIVzqD6AD9PIEGi8N8+4DT
GEThhXWVpnOHqaXiw+A60mBUpF2/UxHRGHbtw4MOsvX6yEv1ut//HyGQ5ToxMmZi
IxrtKm0JBxTMVrgDYYR+NdkkbJU2o0VqquXEBbTsexQ9C/dVfe+vTcHLV9x9BqcN
0uZ4Z+azFgn/6S5k9YK94ixMDeco+xpc7vpS6HxsKskI6GxsjrlqFPNcKe77dnhE
SgF4ohFtwoELwBHP/BrevopTt6DBgc5541MnSRaEmQegQFW174bqTYqlAszFKibd
lLZDDAq3EauD/Nnyx+vchRf+pQEnXLYLoi60VmD1iDXLHxoGWVelDxVc6aExItxc
A8e8PtBPjcNS3ZpPlXSSF6oBYQiDZdPwKi03UJGTGaJX24HJnzZQlLTVlWZwVVH8
BwpR4c7FpDr4rEeGYfWTbDzimLbPe8StQ8ltg5HOALrGgdtmyPv9jXLpGRT7ktZu
dbkZNaQT+ic8uw4s5U9VEyc0Ma9Gsa5Ee6dC/HP+JB9J9Edzkv/SodtOEzeQ3Xps
/+qF0Ku5vLKcjXMHsIQYxtxOHMNKidh2KUNW9hGwFsG8geO61Pq3uIdA4jMG8U6V
gA71CIvKLiitftcuUdVHm5NjH0wCnJ2IVUVea8BtNZwYUupj0cscBhNvvr3L5bs3
M2ggmIO23q86dJ+MiHnA3zrtBJ8iMl1CaGtrXovD6UtHpqAyTklMUXN/gc4XlFro
rfSa0Js1ws3KyY+mt1cLL2bhcYDKJK+TxipZwWQ4ujZeBl1KeC4RhhR0FS13kG6b
owGDQyRLA9sWj1hjmabqqNaJSddFhtm1ugQ04o6zLA6agDV6m9ItgSl5ylzLipf0
leByCk80RL1bcDQKBLLzT7+TsEqGdDkzKjiOfsMN5M6tuEYovbEew8hfjU2hXm7e
gUoj6kunuNa82SkavjHEwJfH2ypYZnGFtXI6cNWkNCmBYYfPH5yX9Qat3xlSQprJ
KHkbJaWKxKS30smqYcqIT4fPFzTQWRefTSRKRtn+29swA1riOBDBqfFchfsz/k7w
JYhQoQmxtKoisOD6gLsa/pCfuEkZnXNwy6wbtbhBqx1hgryH7xDNGLjAI5Sog8QH
td2ceCV/jg+F4y1daVD1aPc8htTsSqICMubndHiqy49kj8rgf0DlrlUrnLp6Pc2G
AUkFvfE2ImoPJXmJCs+byfhPSYSGaLBqnG8heVedszChgI6hgsuhwRxkIdAh/LYz
JL7BQKSa9ZfwNo11RjMNbXk/2l5TEQ/wTSSEZ78oK6tMfppJDqQzDBDC0lTEwA9I
el/lovZjkY3VpNf6BhY85s1JmTZECIdRuhvOwlU6Kspyii+ejQw3E7+1GmMv5SU7
sIcamsG43cr62mhBmAvG0k7i7SbiiBX+tSzrHwO4PMnUv8nvmLmvLG3SQl5d7t0q
nkHRFUxx3oRwCWWrYZmUSZ/fSw83URX+XW23gtprT0iei61a6MKa5DKvtndNHDjs
08G+rzY6l3hYCGS4tx9bzCPeQ2c1soSqa2VqZhKYHkl6hdAjiyivBuxAJe4YFdxX
c1m8g2Q/VbUUUGSipXY3d/8vCL1Rq0lWESfd1gvz4KL6JW0ly/A0rQ+c6gD5N8Fr
cLi06If+HJ3/g55BRJoQ38hmjK9CaoqKNT4h327SojEQrccRWhRujd98zp2tPXgY
dXc97HYluuiOFcghV6VbP/PcfmhaLPAcOJxVjzXtU+RR54JikLTtQ1gS5SjeV6cy
Y91fXzXoKPkBS5Yp8W6lAXqlTSov8uq0TUCjiLP9yu/MW9ZurWYLtZ27hrsmijyH
wenYNdYY/r8EWP5Rn92+49142h/5tOSACmpo0M74zM0h/k1UazHMdQ9DIprqRt41
/YYVLf1xkEiAguxB0GloFb4eJWcwxj/pB7Bbo6Y4dpk8LijcW8rFaAoh7HpzUE2A
KpYtorUVqsOcQV1o82SFPJGdexGNkSBs49QxkI0DanJKY4XFDSjr2E/XxrK4SJIf
TWBSZK6fTCRO6/b/ALNlCREfS8ak3K5OEy5tXRDeeN7yN+f3bPciMlew8p/t1NVS
3dGuyv35KEXqshjgxFAT2PEYvhbLnVO1VoHw4Cf+GFT01qB8ZL2q5fsbJEAMO0bf
aqfSwXWwKOfeeZub35aYfL1zRse3tSb6dXsUBt+3g5DMZkiEG0K6iZzD/LPuwR4P
KQjpdFpGbkrp/vPTm+GZesQ0cKx7uQ0Kt1Wb/qF8ox9VFIXiqRfd2lqVF9UtP7b/
5JBjKbNpCxUubwYUUuQJUdfUpRS6XfQWgFfUrSNdKfbh5Hz1JC85ba+hqEt6Mh88
sf9rFwzdBxMidEcurGBItZkGzeQRx70ge1h4XXOSBqn6TSL4Xr80UZ2BH+czDgmx
saPilqWZrX1SsiJIQl2P6aQeHKb8AbCGqjsoghEy1gm68qg5vJp1SF4FrQK79xkU
QB+naW6OJby2I87oQd6mRYviLBly1cfHXvz7Ig2/NMGjv7Uhq04C7OKo/rl/Tb4n
6mpyMVM5ZYha3LJB/nTMWeEgQfdXJoUtzTJnmirh+DCDRMyzXmbl9JhIrQ3Yj9qY
8pZP15W/l8OtMQ9bGucrhNCYaIPXXWJF7JBqD+Zo8iMQA/GkWqJ/x3mIyFZzlQbD
8vgWp6hscZFB/YBEo91faE01P9XrZeGeip5xALHUDWgc+7CqnKi0Aa4JpANXzsew
3hHAPFrOG64nhDLlWM3VUEcV2Cqg3cHulzWs/ik2vpponWvRGxkaH3JFnGMoSPiN
MiEd7CCien6vV78kH7phOIzG/nRQIlK8baBQxo4HEX9XSIaW5XlfRkrsgGpG3zMu
qGrJ+opaBBYqF/idini7zwAVU7T9QFUV+Nlm4tgkOjlkDMVGZCY2TxAK3vTbQwJF
DDHlVpEyAkUju+jtg0cT8SFpznBzL5E5LtHHNk3lFXV+izoxz3mEQlLQ9hRxzSbB
MlmIsdQp2qLvuYpeb85e+EbwwaDsfcxp/qqKD1EectC3Ci5j/rThKc/x3kiTWDLi
mG7AyVnhaESitTA95KLZjV4EFC/4AyxONcsofcTxl2zkfgat82RjM9PGZvZrGI/Z
PKgddfzy5Jgh7P9R4L3D3MMRA08/uDkIHuN+xA40hptXcjfI+7IjyxjxrDTNbJhP
5TMWr9pwl3yldrnNQ3xFI2r0HQUud/P/ME9bLVPQBK8FsTjl++UdRjlPXWRlxpri
W60BLv41CDW+c5G+ueXkSfW0fVvXkpppoY4Atw/gZh3h/Vd73u9HHBg5XLOlSUI0
Q0+1TM+9kG683+Cs2nMynW4jGbO6GlPcDhO+aYX/3DHuoAxoDSpp00b93djOh8yY
eWFOKxOGrUqksDVk0pezpQwIhrtugyRR5qoBCPXqGpovC/dUMGuhd371qJyclgEk
E3uMfHequCU+PrYBwtCn610cTnyF8wKJA1/Q87wFM1n+LQfbKUMf/71R4isDn8pm
4GEVLwsLx2tiK1ZyazLmSLAHLLuvxjXWNPnBbPBejbkRP3O46ygdstbHcCfhhzfK
hvV6zhPIGxJj71El1mYeLeTQf4qEYrChgBAFUePjDHFxXdVRRHlws5boDIm8Ct0e
kG4X1p7kFfMZ/e+Bi26QIWgWMDlLZlb7DtHS3wDSqQnb/oTsvure0SZXddNdJ3JC
FiTlrwSlx2dh0g5mQFvxTfdQdKllPf1+nfqxWb5n2dnifua7HP1RiA9pynfmOOWA
5SOuVvBFo6bj8ndXI/eb9YjfHcx0pIYysKCyaJkbOl7ryE0jGxtxHGFWp/WJDbO9
vEYdOLGhvszDTIq+0LiwA9MyNkPOdaLzu7ZPUeMHFvCYqRiR2oIZakS648NAMkVi
1PuQSCbcCqWnUxuigf7EVoReunAkNn6K6Y89CeSFn7nc7VCe5k+jFXKM29nsq8U7
mCQzrz9wYcn/cZsfGK9B1ApDDxvLbxw/PeoN73/AtIjPaVj/8YwX6CA/obu3s06C
Sw0/F4ibJYU1dR0Ri0Si7/9wO+B7gB7xpkbAxfhOUp1xeBFoTtQ15NdH7YEyd6zo
sz5GVkwoNPdtw6BzrSEa+xDU/OogN8CY1cORhrO0iutFe7k/LAZqNz+dXw1VLNXH
DdT2n+lt0z28+a7miQhhn50WanfnOEiJDwUs3g4LBUlTOwL9B2U/OjCu6TmEbBov
npCUI49RN1FrKUYF/Z9N2CPGIG7Qp1ztjhzofETn62DROXT713c4XQOXtfanGpkv
c0NqjZ/kXBEXMhNtAuZWUd7PSYju3p7nx/ejW2eS6Y0QMBIme7hNL6ldP/P1GfGv
uuKkzf0Q9d0TS7DqhHywmhYEc61r0ra9QIKJAj3fDmHZCTSihbgLr4gVMhUiMRWy
TdE1mzbyOR9eTo5hMhdKo06zDSUd18d4DxJs9GMuy7uvOYex68FIdJellmxAysmD
8eEkEdMQSXa/i6aPQJ2EYyl9hm/3i4ppADkQ8EyLXpyvVR4G6SIQQWQJG4+/Fv2y
p/EwZgITjx6mhPLegTG+jOWRjEvZuZWIj+bmnrod/0hsIV/s8zMpLBAl0EMUTeOh
74RGFGco7Jk5457mkXFwn6bgUV+de+JNtDo3vDUxFZyLj6PNf86JxryzT3Jk5OMP
hALHW7AwJLFtoneuGq+I/MSvrCHrW5cSBgzeov+6ixM5/XpAbHLKbObsurdN8JJN
ycmhRYIKWRTSCXICFZeykbJW6EDpPu8b1HNWtSqGa4ManEI/ZLTYzr/FDMgGink8
/Y/KpMDts7m1YMao2H7TKaEGgKLwk31rfGMNKgx9Eur0QOkaZE7klsf9Ru3Wf4Rm
az0yBZt+vzPb3NRQuRy6/XulazDuuJWOf6dRB7FgCJcZbWlGmCguNQTNZE2yJLtb
gKbBt3Tu2WBku3XNhCo0p0IMq+j8Yziy1qReNJtlr5O7oGLG9hoBcmgyrMmly923
amiMBX/Vt7RBy6S9KMJ3WTgWMbkVUBmOi9nmtMkK56Codiixmj1R9Qe65LRLsF8X
LCLVDMjounEXJMupzDSNpgLl87ZcPsXs/wJkBDW+r0VHLGeThWHUyqZBS+VtzWH2
LvB6vnWNCtqqVyoA+1PUsP6iYamFUQ2kOXkOKqOvJIxQd+dKsVQvsE8ISzlwqEh6
9gY/qqFS+m3LMca6HlvjKOiV/xzxSz9xpnycj7Zja8gxz2C4WsSlArHAnBWpAzu+
WfHG5lSbu1Kqsho1qcAreWoLblr2Zpvt81g+hBxJvpOOm/0gaSCFCOvLHho7mRRq
RSROvDomYrqG0cp6um1SZaTO7waSEjIA1dEt/LtRl9bRnKKH66yL6euqk5huvNCQ
GOD3tyJbKgZTdtLGT4AjGdaFxT9tcDpgREr3uFOJNjlY3qoNLMQ1PniOJz1TXXcG
B0SZteHlKETMi/1bryev88npcQXtW7yI+l8+ervdgOTn6LzT6E/TpGmxHoKJIu6A
ry6zBFT0FOyeJDxiw8pMUMlmPVtAOtkNpzSzLR6I00jza1bvMENzb5AhZcAQ7yQ6
Gj/nx6a7Q8y3XaTG2DGCzp/lN+Y/pWX+c+rhZ+RAO7lWOZ2M67mKnBODmwWcYotU
TYd9Nxe0uu/WYPyEintyEu3vLGuEYAktZwoIJQBWB8kO7JrgPv4K6CB3VU3zwEMS
VVz4qYEgUfxGUXjQcQATE0P1by18HUbT4lPlT3QFgb9S4X1I/LzS0068EeRd7gZf
kSFb/ZsBCqfkmxuoixDpdrB7og0QxMmkdeMh+HKy8HAX88VDa29cG0LYXJ/bVyuv
ppHBTss4QmGTD/vHr3vJhRjzUdnE1lFe3QINkVJjgTsQXAuyuPP7fw3gmHZSY8p6
duhT6e78uw9GdECo+VPElLSsGKuTdM1mJypmkD2wWnu40eCeKm/YBgA86YPK24cS
0UHFHLDzT8loArS84ezO8tp/OV1gLW8YTACI4C4W++xlsAwDoJpUS323esTlBVUA
2JqMHUtVDgCZAgl2MaZlgOOQrhphySR9I/Tgp1ACZcyFLX83zEJVqCnBUC1cpoCR
B8MMX+w5JwralMscmNOmcINX6DnzoCXhldKXpo3e2z5IWuK34XwpPx38rKFs/sLK
SpSUxHV/DoLjG023AWORKcRe5aEpo4cxBqmHYp5sl4XzCj7xhYqBBwzlzyQIMlcY
yP2990+yiuqXZeqIeUapBLvRcz2/VW35O2SPUOUFRUcKs8aRyCGZwOhn2t6Zrl0Q
ZE6j6/8jV7NMjCA5ittY0ePgWGWaXaLLXSgNWpCYoUCO4yfCNKv4TkQldyD+bZzO
ed74ZeyVYnSgeMgFrUaPitqkGzEtACD2ie/MNm1yVZnZnj+kSe3jT9x52xqXKa7u
U0+p+3TttsrxsNNeW1ezz4ht4Am/uD/9t7dMQJlFSpOLT0oMONWw1bGUcxrgWugK
CRIDnMMun8Pm4q6oO7DXag3q8y1r1Nsp6eYhsLdIgkHdw6c+51QCm/w/NESNltjS
WLheIpX8litge8KOOFirSWXnFJ3QIwyBb9y0YwW1aAeeabSn7WllIc5YNZr0coUC
aeUSF2vx1ST0qTk16AWYzPUf/uwhUVone3AWTsmeYqYkbTCNW8lpvHjl6BjJApX4
o+dDKY5awgtXGRS3ybh9oOBPECi/PKy/4dmOMjZX7b7GdZtKwSjWMwTIVLk6W5J1
oWTj8af9DWQpQPH0AO5J4UnKDWLGfXAKztbPxgmueQvlbzjltcGoTy7AtpAZI9aW
n8bgBhY5Hbwx04vIL5yxIAOIekPo6RN25vQqDoqeFGiQAyWX6kwZy0JRuZwvoAWy
cH6IQAn4a+jSddtxZk37AyiNg9oE6pDEbIOX6SSRFM5U6zOE8EcJPArTkawt0N0C
dQmk2SVa993zk7QpJOPczb2CbUK4ehnH1xTN7Er4tP0oeeRMKROKZwnjSWTvfV5x
8fhQkYdItnunESjKeEsgVnEUeh5UZLAulPpwa7bLY/+nYtkowBASc45hqlkWn4oI
0YNCtnGxqdVkS7psZwBEhLCNcAlKX4HDzcdtO9yqVKtrRef+IcRVMdZL0sD+dA7i
gfKum13kbw5k7LcP7dbPRPTEacPmS3MRihy12C85xGrZtryLldTx3Gi3o3ukLOxi
jHwV53JhCTywRS1UfcXjpcn53miZGNzOGU91KSIOrjZh3vnH6dyqMHms4yckMxj2
Mi11wywPhjyvaSY8Dw3w7Op0KOEFGg4ToFLbhMwKsYvXoLrZZy/ZhHXDQb2F1HrC
PSwZcx5KeZbTgZvHKmxwbeuY2hSDvnzolI5UIPVZshJdBE/KG60Judfa4GSN0y/3
TrkH/o5rzOkdFoyRRYL2K88luK19i1bLtKj4hGbwODn73bsUlfq7RY6XcQF+bcBT
BvE72mx3uNco0CZ1NNhuT/HT6pNVKu4/7LZQ9VERgdoksBtZdOj0Pv5KSkGTfG9O
Pn/ZcbQdQ7niNmSPzaPadm6MEfY/VYT2KrEXa38EFErvCqoGBoyUgiDEt6CukO5h
QY/UkrCxa60oz3hngZRrcjQiK9YcqgGX+rgKYGjtEEVbVHTEzol+ZMH50QCDKBnG
R1LJd8XqIlJvxNA16uT5mK3Wk3S3VaxQjrZ/VvenamHFsn53ePmq/FCY0mJklwf3
MYiVeiJ8fnxCWiVfjce9qzNfh0O9f5vxm+2EyhZdSwQIfS8seuxeT/ZTOIzXt+pM
tIph2gV6LhJxtTuGo/MQevT/GEncJqo/JVfBuT5s/Q+VEIixxqABPPA0moeoaDiT
DtutuJoir8r1pdncMjO1znJ1MwRiIvSt99Kn4RfGnHUEpoaAuL+RcclUKodjKVjF
ICu9clxDS0Pz7uvni5frtLFwOJep2Ct1PvG7w7xcHCTJvCGLM1TyXwR1GPtJvlMR
9pNp+IuIdc0JAxRmbGcC254otWLJd6N3RilbJ2DIK5JTOEoIrlZzjSYrr8Cym9YJ
UTQwvaxP/zoJV07xY+Egty28Rli2xJWMp3m5Kzln9bmSiD1vWlWbP+J4igNBrLVK
kT7dqRXGRcviSU60F/niXn0VUk9LJQtx24ohmuSUH5a2nwXsh555Hj8VR4MrZGc4
Fa8koPVKReixCWXo7g0aapBtkYZJTXTCgigFBg4UnbhwLADmBfcxLO6w8Uo+tYMA
cKXIn4h8M02nLuOPtNiswOaREdJbc3qB2QBl9nmIDNg7O/kjZobuV4t6qgYAMIRH
noexeRrNCaQYVJtRU4noYhTYqqWljSTumkOOsibOsCCmEkKvA4C8JAzd0SJjgd6l
L+hWDqMQ0siTLoce2SxnH/dgs8BAy0vBcLUj/ubG9OjZRbAX9vHULASOdv/t/HZJ
BH/TGshB/TagzERlbyub/veJxBKypgFHR7ALekfnslSb+IyqflgBoKEgvmEyr6Yc
khDWyt9N5mzHCHNCrCdUcHExH1y16G8OY3kbvnxcTOHP1SEOuUhnm5cYu5B8FvdJ
5GwgvdA03Dl8n5zZuq23PB1DSguryhwiWN+43TIC5t4rh3pcetsrrioz4O45dcsx
CPSjRwf4GRENk9Eu2cpzu0a9B0DZWwxOjBa9shCA/Gy7lqeT752xuMOE+OVO5dve
X5rKFVdKIJ/PKXS9hJwU0wlHHTi5kDwI+pYHOceRgJ+QZ2XAbri4Ypw0mFNyRxdr
07iG6Gmnp375m9PTTUUf1M+I95L3/eBs5k5F5SqYOEmq+sthSV00rRCsX47GXCUV
eiv9j4CkdoK3g9VU+XX/9BWwXRXFVomubuGlfLGEfsiVEQJrFGv/cLd+4c5dtZVh
tMbOeNdNzgzWeYgPuMuUEMQ98b5/641IEK9k9rczE4bJgNKt6JK89NHFSf9Vw2qb
VrauiEzqv+mx7ta0mllOY02d7fa75TGLslxs3RsNKJ0WWNjqUc7MKoR2jpdBUFqI
51AwB1wTyxjost7Itx/nh7C4QyLpqlMtyYxGo13BTWn09ctO4QUItce4QMtTG6jX
5jCP4ROTrwQHy80bfw4SBSrKASqvqVf4I7O+B3Dr/jbdbb+7TKJGQMk9iVNQSrj8
M9D/NIsietJvPHgq1iM3jEB/jUPgPbeRLwZeXjmWIltDBLEoqFgKhE1cWzRlO+iq
48BnOcGsoJ4Iwtj8E1nHfrH7CltJRdruognULiXlPJNjiyTy7PDXT4ROMEgQz9F7
PiFJGOpnaM5a1AEw7W0MuvpqpSuZ9kZDgAznu/fb+ExgqFTieY5hcIrd5JdwCxLs
qgpnj0WwkQjOaPB8OJGOt4Ml3VN3xYs6RVqwKUTlWArKx/PTHSnsD72KnVgObPBB
ip/iUxhYGlyF+bIFHIVTvgbNXhzgEcVj9jU86plO5tZNw4+jZmXtxVfufaVij/rm
BDO+6XlDRltRCn3Z9FgfnJBl8gzKR2PmNp0PCIrTv3xE7JlaFo+oi14j7s08z/DB
ApAssH617pXLOeY7VSD97alOBeF+3Z2Of/EMT5YYnnvl+3fyJNIbVbpHZ1/nXm6v
iEWLjcGOgVcaXhtt3KO8nEmd7ff/M1CYVf4oxXSHEKnglXQesarNlnzW7PUOIaOj
ETFUBGg1lGMi0HOLig7UttET8I73Uid40EFfwF6x1Wacm9pc6/rZTyKK/0ZwF3K7
f6EZJhpbnHvbqcfQPTA7qPLAAcK6+SIqgZ+YNpr+HG0H5HWwRIoNIST3W7FiPpd6
q3F2a8pEzRpNV1JgaMEJbYy3JVgG4AA88U1a3VNtGKkdUZHerJrypp09KFlzuHel
d7C9+ScgZXCjUjcv7moAUi0mnKsfjTKGpdtdRch3wLgaXnTRcGIDOaSEANf8zjnK
i3X4JwXXvlDsOrMGwTo/O0SvWQCXJa1d7w8Twd3KICi4at0sp6o1rlDhrKzTNiHJ
OloPjS9VfDcdQRnmrnd1bX2tsfhzVTxs22i9Ut/BZOppF2XBK/Pvj7Gj+7uLviPP
wE6hgQAyhgbIyDQAilw6ehGAsz7/NB4alAPyEwwLNf3747r85FQBJ1wwwu0cDo+L
ef8s17C5Eqy0gK20r8so/QIDNXQv+IENTkeq+7UNMm5s+wU36bmj3TsynU0i+L/m
MP6mHgxPKavka1+y0gw+R4XMo1h6tiA+QihqrxNvmulhPvhsbK/xtQmmHPWC5UlN
WzrsL4GQA3zsF86l7Jik+p1H7w8BxvtQFw5PdBnNlBRdnvUwhe+QsTkPzHHPRSmO
oqaJyVd2hO8cNpmoSQYDb6RbWxhdYCN3oiRKoNyFF4/YEdHa5US/eAWvqRECOMa3
qwS+puQ75BYZOiJ5injfvk3sey4f/hTyY/bGlnAFvL/YOdb0qDCssUb7PZV2Idst
zWk8Tl46ZKbJSrrVAFydW5xuRTSQk9QRfzKBxWo9CnxlpGsdJqV22k7jr8s1K7z7
5OXPWYvkNNKoC/Osoth8RixjYsIFgNzrnYcaR+c2vPX9URZadYJ3Cf35KwL0WfoQ
s7cYPdFnuBl80OA/IL+aY1UN9mxrM+pmEicQH2bnrm5Cq7fXyDgcyHicLVmBKPaE
dK+TKJxOrwfjl9SfcE8pAQ+h8MQIXtwBnCQ9lLJ/ZlaT5infWIGe5YMl3W5t7f4d
RNGgD9hpugpTD1iIifCWaTDjKjYzJPYyBXIMg90VGhWYjXcATT3wazJo6sGnrC4X
2Uzg527qRUf0F3ZFLYUFfgmsuj2Ltlk+MwlaUMldJrNqz5RkDhmwZF3R16GNkTKT
QASLHhHtNePbbz5P8Gd53eGBJnRXjNLQxbwV+sID4owKkN/wFAgHf5e51HtvIEnc
Z3H86YYVE0m0FKT27F51rPP9zMReGyPMLUUsR+Ok5HhH3Dd+JYEdxPb8evO/zVXw
Gpj3SZqXwj8b4KcJ6AAone1q8jspEKTPH+v996VHAjlyPnqQjtyxVqC6D3S7e+j1
WI0d/QhzndVVZwRZCX+pFIXT7Efvw9AojhzG76h5JNzDG0oJ+0aiqUu02eTVD/Hu
QWRIaQtHjEWKKrUlmlmuVom6Kdqg/6SZKgn4gcXKshh0rrorgzN2dgGsPvG1B2nX
ymo8uJoTTqYLAK663KIfAa8RbmqyIf6Ye+7RvsBr4Jum2H1T3riqlo4Xidi8uIRk
CgGIf1HnLW8OGgpjKa8FIFiR1+xS+mwPUG7Y7IjHHiHWtMiFV2FfgRsWTZn9dj7L
+IE1+3RY7JcrP6ZrWfnpdvXeDmk30dLZ/Fukk514LlnQdh/JbctxEr5xhNaY1HD4
sZGP4Z0P2pc/lILE0tLhstRTExyLli4ZRtDjs2scV+6lhUArwDZ/eTlhKcMOof62
P/53eUdpy2imJez0xgJnWPmmo6lpd7iPWK8otJMUxakVYAL2SqZKPMHGELFfLOac
KKzSORlsWGq5Fyf1i1Zk8iGghMsxnOjgHfGA4DsRRd2LHlxnNIIeVNwKtd9QjuxF
tQmDpw9cf8TbHZhHF0jfLT2B3gv0OG8NxqIobGWs+A8jT+UD3TPavTbp3rzRnFG+
WyOJGZwXqXk3eq6KntwPt1O8y60smVon/QHaifyKNGoBsZZw69AE/YVN8pZwItmJ
Li91gGv2F+WYaE188IJLOAJrZghoTg7VGTUPrvYagQ2CD0k8SFXlyZw+HebWSat+
QEUZZm/lfo2y4L8SFk7gPDqMLFz8JfpJakV9SPXxERcvXAIAs5o901GuFaorPBWR
oGwaxcw1AsoQBOuiEmjeEsh7CyZqw3/BbVQ1CUpctcO6ssrLOqsNQIUDWa5XgpVb
j2Og+DBI11r998F/B7MxkAnvllj0miArO3s9Bb76S1AUKW7gJLJ06JY9FuZnryWD
zbwVwrCfD5BZjH9NpFFvdqqP0QP1e5+MdbozW5Yp+2Hd4Gu6L0LZoePmjSA2Tt2G
W7NqLfX0eZ6D32/QJrKcxNMcTs8CJfRw37uI3Y0AOCF+/jx+NnjGGKM2B1OmqKX8
ZnS8FmXpE9/+2yWpQvsYKLxxDKhpkJT/NaKi+1K4dwb+KwGAWlKE/ZWSpDq/W/3M
NjijdZxofkaYVne62rGQpmPG9CG4u+5JzlTPSkZYk3lAEv4A0t16W4h6KfHSkqHN
RSzkZzaSzvgCr4FYDyNR2opo0Pn1+uzHV3vIQW7nI0Kw5lTUONQoL3abPvsOeV1x
`pragma protect end_protected
