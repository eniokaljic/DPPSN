// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:33 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XX0ns6tNi5vFL/NQ76TBtDHCHbEslH30C8kM3IpSlLhMRgwNDttzCZ9Dzea069Xi
PSw2XLk/leylKo8IxIs38tNd9rssWczthJwyViPD3sS8I4kAfFyNBusxkXb7cRj1
12OSPVf6h/M6m/rBlNz/Uc8yPd+YR76cEFxEpl+BPKk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4208)
CwlO+l44xeqQPPwBSKCHcCbKpMEvM+JvOjthFxa95r3LlWsonZ8aA6O4iyavXbYP
AzGvczYlA/mmrkWrgjvRo35ZHi8FGTPhP/SseNWxr1iGw2hxaI1Z/hUuQql0W9JG
EtvZIcvoGyZ70mn7qVK7kD/tn6feUVdlzfYLTxBbJejqB0A/MizZuxT3zCY6L91g
vdpBN6tUOiDP/0h4PKe7JHhXdakxj9rdKu2CvAySzTVoZI4z/ZU8L3zhv+8/nDXA
FNp71+F+eusXxsuXMgs1tJJhr/OxHGIgeOcPRKri+37NXBT+nuQqWvwVb+v97fTA
5IpyUyUO6hFbLctfM6vtE6xr7n9RusOLlZKouVAcnE7jkXW6P9Q4IKu3TzYntiSP
pO+APZqsAnTll0gf9xx8uqMzIIUeOQrq9JlTRlJZcXWGy0s3N3B8cqnWUJyYowWw
T48xBOE6o4IvUJnvvd1NdK1jGaP2Yp+H0Gc/R2ZFugARSnh+V+cB0dX7+5e6BBG3
xF6u/GA7c59vyOSd+/SI7Nz3Mr0nie+mC+8hvOnv01/Gle8mCxlcQ2iCF9oCraU+
1mIxtGZhU6YvthsKlV1nuDHh2CNQIXleGIxo3goaHmFowjBo74lCppTLYN4Kyd/c
mqK48DTGIRtx6VUz8LErwvf92M2z51jJi+TeFWhHSm0Hh/mo3mOvA7qeuDFOfUS1
e/PWkMueZby98wu+EbkaeDwZ30BdL9DUkNFA4YfoTK0p6/Yw2zJZEVjAV72dlaP1
goVVsOjlW+pVsPTqV4IQsOVO+QReZY+x4kLUfYH1otcdTdRQuZfrGS5QPeRlFIrq
l2b1a6xfp+ZedkULRJffrrxNG+yH7elhPdAwnHnp8+pBGuoZ9DXeB3F7YYCkY0TQ
psKV6Tyi+d3QN49KmgeGsdxdKpSyl3tPGwvTf0F+ZGAT14eJCTHlqOzyhjwHE+ZA
E0/EhrbqZqEgtu1B80kLmBxUAKdheQMzSwdsEI2849iuqFa9VryQsXj3vNvc2jdS
NM7ArV9ZE7J2gUx0G/30yH3I/PfwDgurRusmge5NokSEJik8Ex1g9SsEXN1o2Agx
o2dvOC5UHBx5xfD4hdasfBY1/AOM/ijhl13lSeGQwaLTHIGOnCgPYhbmtbUkiG9H
3oUVti4rQd7kCl8v2W1a44w0kfVmHIcW5NiJH+cZ4DfA78XtpzqhdNjcvU7qSmjd
b+ONinwfY8lT/DhjI2AxI9sx8mnie1Uo0n0Lyzlta7cOsEqX7NRqi0eE1kSDCPlT
H9NZ/znexU3zbsDon5EjEJ/i7lqFKi2b5A3nitIQVYLhGPYFdy4HlhGa2bfCOL1p
6zOO+gOzTnuIU80rPZ1KzvHi3Y3hvLOrnmOljpVxgabctdPIIcdIT6BPD7KKhNSX
rvo6l7UH5zPt+Cq30N+WfWRVhxGQeQL9XAaBuDbGWYeMqY1Z4I9S+5bxaOhw3zcy
dRIlsmhJ1YLmghPcpJ0GGuFiajNIBRDCAP7ko0/bbZjkrk2z3T2pW8jXiQGzclk7
nMWYPIwmXIteHqmoh4bgrp7OsWJ0Mns77Mn31wFnc4AZ+Tnz8PlEcCJVw+zNBVg0
9FVkdaIa2E/904MXoL0lJHSM2lRNUHu+qVG1vSwvHPRm6sn89v26IpYuR2yxeNfW
I8lFwA0vzh0aCsFy2vEmSSGDYPagKTqAj8IezZkbdZ9Bco/wJFnjBdCQwak/oKC/
KLfCiVHwrbev6lyRociLb5PI+kfwKbvgBqGQIyCZHRAJlhqZojjm2eui4iQlRf69
6lrTi5ZvKFBl8thMPEDr37Tzk5gexsOcHbGLXRbpIxZ112uwod17kd8VWSKGLFeR
5NzuQT/dpFb+2bkCcsOyDdo894dSqhmneL8VOb9o0DS6YIfNKwpgTkfZArx2/HqB
MUKa1P+hMJs/Itmz4nYMsFQM7KQ4nICMO8zz8Xif3avgN0J1TcMfAS1Io4W2GzPx
ZiNsr6xWfxM7s1gBlQOk1N0BlZZhGQpyhGNwx9CYzmyLjn/VpodyhtWpNfo9JSjU
b/CdeZxP4WRWc5Bf6kVavvOTKEjKgXAjuhTxMIdgLnryTY1rFdlpTdj8ZtxvVAgO
afYbuvITkJsF66eorK9c5mJQUVRRdDvJ2dlQtFMNZHQs/C3ImKwc8xseTnz8Dm8u
wrS2CT8tKDK0CKYdYBegbin6Be8ptKlYG/K15z4eHKkhH/GHap49KcAb7cuD4TeA
3WWxgdPjgazMQEuab+geZC9P/ljUowwsmqM90GI1A1+bgl2JsM/zWRQpQUXa/WHB
+n1PBQWLXwWkO9kZ6V3XdJLZzp9BZ5eKYDQ4c7lHu6uL7g7prL/pq+pxmyZE9l5f
IUzOAKz/gEgQEtOp4P01D/63ntFA5WcorRp+WKVnhUvbPaSDpE7IWqb9dLs6LauR
19W6Gj9ELWPTDRaCKBS5q3EsBecvKF24VUjreOgpaxU7tpl78NSUPscdALtSdXPx
1Y/cBR7rB2hM3tg3elWw9Qu1WvCZnLs/uW6y8PbDTvp36uhko3K5j7qFGjY7tmwf
CtzcN3qAKZ5bKetFzIV1U0RnTMl14fNiLei0KisYSGC4HUtWtZMUy2yDOgSzHwbn
8lJ59mIeXf6zgF0uTT34OBfKFFH7GNUg+sXzcYh9b4nj6i/vCg/Sict9xx+Ak4Gf
wVHTEmojktXrTXrIWDF75WRiTkmBKGXy5ACIfKi3+MCKMcoriZD7KvDkRa0w3B3M
jj1MDGqp0aLAdW+1cs34mrBp4cZji4GlMJEsUwWAFoBy1s2dnfTrjZbFstbkoVki
2pncJa8Pf8dd4CIQZawmqch2HhMErCAzoqLPspU9rscvTvre4Zh16/v4/iRipgyz
bKvWVNtOty4art9QuRwh5CZOb962Rr58uFHsCU/ZW9W7Si6NgsqDPmDEQfpnQmAp
i1ccvk1LAyrJXmIaVXVbTD55nV4KR+g8p6NLRJ5CR+QvOODT9dQoqxiwN/H9FovU
kI1PB+KkUVXcmU5Vm0uVodFwZPZ0ISuE8A1upEB416vmzIXzij/G3eYjUgIbd5h0
fu5+vw3DI3EDqFVx0mv8s7ScL2hvYPOEF1DsGAQ1oAWiwHvzsH7RSLVv7k1KwxtS
16GvLjLbTCWYsSxRhziKSX3K/x801PfoaBDNPIzESCAKdhNgCuyHTPeuUHkc+S4E
RiNIUDgZKz6piITpdZpPopDC9Qz1RjrmCupMAV5XA5ShbyW7eWeo5On6xXDPQQ7w
1lyvwf+3LkOfBAfBJr18KYvWTXDGwWXT1LaF1OKvS8RYm7zh7J03vbbbC0znjAuF
BIu5ITuQGMpNDLC5CzHCGlFpW9kQDf51rXsAk8pXg5pgKV6n9PhmAnJVQPQasN5w
KtM7DsWe+Qu/yofwT2Klj/JD/hhhEu5KuywFaJA8P+p0q/wM5VLc6T7NfZSN0NkS
OZV9uFiLeY7B8NEkpkJpWHoQiMw7/LfOwmqP4bigRblHgUuXwJl8Y8WTL/pwoSAH
8ckL+xxaGJq8wYTFszMFnccqqnUgmXzQVXVk5U84wYx/0BlInEyHMI0bOuDAqP2r
OdT8YV2Vs0a0QWgJKn3OlkZmh8uWabWtxvyFnMyWSaxNLd7u/LbXhziP65x4GvwO
a19ledgbfty4jh7pA7/PJ6DLzJ3ketpSNLhh8IQLqRxjuL0zX8FyJI861WzzXOs6
/q+9DKs8g+40X1P0D+q+eswlwQMj+ZDPCkMUknt1e1mhI7lmGF2d4EiMkCJwsafK
iXA3HXwWwpF+EQIRwvirWjObiLUtaieHHFt6QIwD16z6QMnLDktNYpezog1uhpaD
eLeeBO/0rom6nFQcr9tMp6P74uysoXuHl1ekiFd5SF9SmosiVGNmSzIAJUNUvsG9
NEDyGTcygA3TYEG9bxyri9ASSc6YlZmo0xM+wWPJOwDJWfdobmoMXEaDD5yy1rNV
1cHow/2XX2SEZEnKhzlcFshgw28JgnZBG5k5yTlorVYMtofWpY+6CiXKUThP45DL
w9KZxFZVzMJ2m0LkvGftnc0I2RWhE4Y7e9sEuidJKwlr9/SD/44Cg2zCGVMfl+kY
5q1YMbfenSeGk8tCyWe95Q3ZwLeoHYcE674FCIkZX19vBtmkEwHENTy51S0AYU4I
fbO72nZFWkvJowbfOK3htQW/jT0I/5DbT8QDrpXk2MTwcUwJCTH6y3kSxLMthRss
SfzqxxAaVYqGqniOQaAeyz5UOngYaBDLd/ULLVK0t8KvbH8LDWxbXS+z5T5QYCZY
rUJzsUA6K1Sw0Nl8mIph3MjlQeXQaBcg2zVt8BwfvtMFhly/EjO1m/ERc0sYkXCO
MlkSn9LILRccT/Os9eV83bzBB6oicQovEKG/yO5JnlohtJZl+6xeDy3fKODDydW5
jnhjgsnPW+72GpWMgn/ZJTv1BKf0DGG0hy83KIQ3uFozDrYy0q7nIs/36A2+squa
ZweakO0v07ZZkk6+BRQoP7UzhRAZAO/hv8OKZvc2D3Ixib2zN9Tfs4Pci6IBYGqW
wRwuustpN7q5h2/Z16fRLZ8FUR8dcK/uMkP2Bcn8WSZeAyKLQ0PVyCfbwlgIu347
4WfHkrQPhUHNLiPh9hbvdSNXi4JW2+GIzM+ds6o4Lo4EE/iNeZFpH4SnUs4A4IOS
ZCruCFtYbxsslUUXjDcsJv4uiJAQsBNDwKiagh5a6N7rKJkXbm8d/nAalpGf9EGZ
18vakfGddlTXHtNvDIwz0y9yChUnIFEhBvSOVGv2r2mPgoGh/lDTJFh8ihoEcWQ+
1t7+OxmAfztTzqRpMpDqwCQ43toPTbyQqFVdLybzwAQ9tp/HXtx9r7OLpnhBophT
WnID5dGxZN7fy7dUtfmIWVpcddg/V/GDnmXzFAn+F+l9E6bIsmzr7QFdgk6yya9j
4O2L8ZSLf3+wQT/z5uQdhaIRLqDhGpFDewWan4fprj9Xnq+7eg6e6AIC61MrB3aH
3tBkLnVDWtN0jcx84XPRETJazCo1dPusJdID8NHkw/07EgW30JQn+p1w70TC0kZP
iW3ufvSysuTiPgq8UyJTwwffWpysg7eRi/7KsEET3P5GPciYaIaVQO6SV/QRreKk
rzq/NQFHhf0KmszQ40wh+2zqlnzKs6hAnW0QnlwQcxkh0SYb1nHEShvVLbdwK/Ba
KWb+ZuAZcdTn9CkkpPyPXB4TzYxe4L6czLIiIp1OKifazZSaE81LXkdJ3W4Huih5
L3WaeyUKcF+z0ugw6JNNJti8XarcVHQbZoxBnr9B/maVKYZ2Ycqc5q6HMF7xPkV4
XoMvo3eWx3Ya3V4jCr+3Sui5cCdRmc8p0VEEOyK2UcjXlGIXIkwQ3TyiCq9PPVHG
r5V6acuSP9ZMhizr7Xpz7nyNF67GMZrbuFyKfznYE562E+2lsvMixnM6P00Y8e6D
lvVshLwkKCH/j2OTolWRbx9JXGLVjU3OxUaof4Sk8KLpQL/qHLHjDi2+x2rG44r/
Lmdr3bVv3R5ox2EcRtanCElN16g0XkXrSM1+6DMaIy/1GJEMrHSZpGCuGnQmHkTT
uAK4WEFrD6Trf+QGTzT/E5YUnB/Veus99NeZv/cUIio=
`pragma protect end_protected
