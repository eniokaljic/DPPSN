// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qvROqc7f7km/sW4lQM8fPsWCqftWigPrVabHlC9OBlu90TvRS1clfySbcl/DuhwW
gstKFMvWnowKM+KNJXeST0AqoD7osE7BqZt8mrMJ/G48nNy2iYTC+Do/T77JHISV
r58oarGB1X3KYnUnj0PWkencEZFc6AKyhOSSeoTkXjg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
YMtBXtA/CrZ8R0ZQb8CdjcLr9IjmSXdmNd643MvFNa+ie0YrV8IIMdkodcBWenoR
yO2LoB25tyGr695xvq5pV9W9Uz4je5XkSWlIw24z+LusgQnKPnDoiHgBWAFI48hm
CZ3x6ci4F1UvW20gOBhFLesfKHTwhotuitcwwEgmtVzkrOrHJaU28IEVmvwc9dqU
fPcjuTvnuBOxPqYpVxHPv1jS9WGhkX0KoJApAbI4Qj7Hndgjb2JQrPgmZdFeRZ+r
oY8cyyadn6tX5S9cFFEkfabrtyDLCVru9U5sye9Db08vcdVKQAzUI+uaMicLUKzc
+FORDBm5Ert93OB865/Wlv75nvrnsiqe/euNbna2+uRAZf7YSEQwN5b6vr1xt4ZM
43qVhER49+Ey5liC3m/cY2Tl+zoTY9e4DIL9NjdJs6vEx8+3BAMCQgjwu3W2xpwv
0O9yKod3Xghne9e2RdrmzNzqzgUgf1eEOhr5nz4zZjaKwG/kCVvFx46FX2fA+CgD
2lr9+D+S0OIcXZ0pyf6OCEzrmh1jJNn/LAi6tJoDI3m+ebXkb+RNPFo9jM4y+7kP
8RabZWy/odMkJlFy/2gTyWDiDyyydIzaj07vd1ckvZEY+ZrAfjAee7MWDRdiXNhr
3up3vlHMllyTg5Xbu+NO7c+WcMFhsRTE4fFbWEdosYEJRFRsXKK+8x8zqBbaJZ8p
U0gAYDAlTaIY82PLekKxex0rlf2kpcZ+UsE0MjdCRck50nNrNJkHbYgKEggMuPAF
1jk8OEkW9AFbDrpGmJZZf9k/aptt1v/xy8zxIhdY8zrovqEVvKfZwEexj9Ov3wCr
fpdB2gdRGM++HjSzx7/av4mUptU288aNeT9UOh6fT6xyfw6xKuayGVTPpDKyebm7
1GICof6MwKoMkDlee395CKkIoAcVri4avgM0pRIMUuzmWzZB1grr2PzmQXXee0to
Z7PloQY6ENQYISf2VakFUsL0vKGSbWOhQiqzzI+NnuPYqa2Cf7QIwt080zFtx1QD
lcYqONkVWVdh6f8x6TNa8eUCkGeZwt6z3kvBbioD3R3NGirZtKG3UapCKpzqbGaC
j2d52KeyCBloIC75crsgtGou50DreALMVh73ilO1zCMQbgtWXDn3Tbv6kTn6vDxf
F1gVWMXx6hedC5qfDbqfO/JaaKvN1/YdHLiTfKytmAlOnDeUaa6asIwNsDaUATiX
Ypr9k6E/FXYoIpO1U7KDylYh3z9vRDXcWbQYkgq6fAhZO1Pmv9VxmS7VHjEnmw3K
tDHGEbtHFDgSgi4BE/0Oy+TAG94kG+SDixBW+pKsh2O9KD/lYA4yx8ICLg/QunZD
d/g63jA3j9HasSOU7YO4bR8fQJkFXZzTui9/bGrH9odqpSLEarPVbPzT1LDj5tfT
OqRKd7hvYKw2QwvN04uPHXGAU5Nc+pjcVTVYSTHAL0C14mPO8jrwR/OEFdfZ1+c+
4PTWb7nbvptWXnjTb8TLQhsjlpVQ5/UrOUVb08Y9hQQT15RoLjUpetFaSenYVKOa
3U9wzbRp3JL4FhlphPzAeTfbkUCfJrqDn+4X4R9sb63oMs2Qp1Kk9WNoPVsQCgV7
0kGmpsm68GuRtfCeD9iGPIkqJKR4RTt1hdikcozJnwerv+1ZSMzd+iFxrypZXUpT
V7f9QLeaHkKLeS6g0zGeTvEiJWQGdLTP06nWhQ7SmeeQKLYeHpj/MbqvJcfR4VCR
XNmGMJcCcUmJoQGscoGje2koGovBiIDWLU7OROaxFNOCOReN7EyBeThSGpJ7M9za
4fph6nDy5Zvhc+iovSma0VJXSflnxXPoohR2xByWgSuZfJbMBvArb1z3nBO7mV9K
RaURtZHJUypFw9ijJuAYD80VqB2VVDEcEn7w3mr1DinUjZo0Bsu8LtLogDj+P6vD
5Izk+QaniZVxSoJA9DyIDth+YjyeJul6U9hgrgnKEAYPgeij7ee1AVnsRj7GqlbW
SPWsTNjBhnBQF2iZZF9mvwyGOnmSeFZaArb06pk5WOGPWyAdlLn4JC4GCay9O52c
c9/1p6fb7IKLSiPnpaKxfpS68OyDoVeiRgrBxhzt7xFzmBXW8AKkUoeTyNCaa9D+
P5TLDHwHhcnfiMqm1xC7pELDQaZVb5PuTVSH7g+Usa0bRR8uErz45eEVAeY9lEiq
6bQ54kJgUL8exRj1GEHA1Qr1eGzQEJ70QCQswfkXOAMdUje66exAEnw+xGN8n3wS
bOHHe4kjPiRsYDzLTu0YPpU5xw6qC85HWbVY3AiC0+Suz+Me3ZQCXTBfvWfhe58K
mxbegApjv865aSWoY5A8XQQjSxgvIHpuw0CcEiUsWbcr5b4mI92eSjmgK5LRA7fm
jW5VnNMlDR8XfS5ZtI7zN0kpz4L+08L99O0PcSDvTDtKOeok05uAm3iU0qpBtSe2
aVivi+Q87Dnq0tMuN3Re9OfBaQ2GGHTb01siq4MIRYKQMu6tNLaU9cqj5DlPnPhp
k5tCeqXI7zbgy4iDgOvnyFM0OKKc2kTfga+/fTQvHKfLEkYxWnR2a7uwcfkad5x8
preniecxBPcMVuL1JuozidFRblWfltqskFWuI3AIBqiuZJnSSmwaUwG87CG2vRl6
oKU7ZtFkZIjJ315fpcJdAS2vINBBXoVlZcIVU4DZGnDU5IbvmofEMIfLO3MkKVu+
fuVNODmUA/MnvkVx7jJaBK1NOxCJvBj3Jj4k/FISiLlSgHcpnrm4BbIirwBSR/l0
7h6Q6AuESpxdXWXUdGKXk2u40rro7WJp4PzXjV9fWDCPNrMpIC/6gtHE9QGhc0wN
uNe6QL4dHhJj7iQBs5fT8dRgCWRee1Msqoul5JwjAfO/IIazAjNQcTXC7oV/Tow4
noXc+UuuxtNcTbIiVJBnLQhE8e6Uy5fR0halWYFKhLkwRptc3jHqINaFljvK+Ahx
7698O7u5FRpmTSBXKpVphqm1q4KeCvqDc//IScLwEYqH+PEhP5Ce+rnP6PqX+a3a
7Wg6Lz2k5IWmA4GgCtuaRE318EFaLwjNXx7o/t/6gtSy0FBo50eYW8V8FpSD8U5a
r3IE7t1wcWcaXs2qvD3GTUvT5swGkKYYomiOAqOpnQPHAZHbB2WgG/4CqZJqE6qV
x5H9Z6HyHcUTER5PGT3ktBrZUo1ovEmmMQtn8qk3qEMuIQIs9bOQE88utpuItUlV
3K0t03hlTmZQ5kgfTPVXeFBck9nYc+p5XUxytCBndmXbcp4Z75zwK3flDJXXUMI1
/vvJ57VeJNAP9g4qZ4E28dmcL1lPb5hh8owzzvOAxim9AfoyVsyU0tHWBOejdB6P
7RWKXYH3Psb86HjvSxEixsEsAO2K0a8zGUc307lLpFnBouUpTDedSFtjADPyfURk
ZyZeq4ZD/I+M0ZDzQ6XSls1ye69lUzn0SV/dLMp16FKSk6t6e9sc0QYuwYUgE0LF
FseOuQvshvmcZV83Yz4dogrjXaDhdipBjDtK83Ms6wdG7qy+xA+4l8sHr3r7uFXL
xhxHl9zE+RCWdrlabUsNYxhrYOgja1beuDk7RSCm4i9GodDnxwm4hj8lzy2COaa/
P74Qt2wJqTSqq/LtKme31u3xeFXsbPmla81yWKmpp4ikwUwlh63m9s2RI516QaYL
qIcB/LtcacPmAPtJqmq3+aIj18+y5ClKGUic9XUuir1y5LS0cJViLBuXcr4A9hx9
PEzJqohBU65ImAGlERKKOGkl8PvePXBE4380O3IM8j4erQMcxlgs9PqTLyMiuBZP
Gotj8LJLZFOASqlZcm68+EB2u7RrDjLokI8SZmkAR1Ont4A4FyyP5R45u6GwRS+C
mTSu6YETh93cJdQx+26HUmjDqK0qKsdKfRhOMYud9P2QJcJK4yCmf7955FWK/YMw
Us+1afUXiFXGplyLlV0n2qOw/GtJfzmtfI3Oy2c+PDzKXISIkpsnH4gDX8NiN9EN
ad2rJbp1WhyZzEh6nI63ALZAXLXkO52ID8GdjP9n+9mr1lsTjvl0tjipbOXoPDhK
Dz2+XV/H3jVPIFxQuE9i2w==
`pragma protect end_protected
