// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Gn2d7ilxL3jYsrikl3NhZCvsvAikbS9MC9lGhUXkw47eLkegapL5nIBzBvQvCzCv
IREXU8f9YESykTunXhDCEOs8u6ppxnFQGwtUemUWLbBywCChQs3qd9MbtD1+7K9v
jhsFnQqpcY/ZK5KOVRyZifnE4YW3i4upqA93QU1BMWM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31024)
O7vPIIyQ3M/cQJ9qw9QM2C0wDdex6C4WnN+g/RDJCuo5x3uoYZk6GU/YTKarHSki
d19xvI7TjpwFZlIsZqnOt4edyua9M0wwnAkSYyoRbey91ZpZWoqwawjOYhU60X3B
njMcffC2ubdBchkKIlb8IMBxBG1v5tM3AY42JYWmbByPXTRKUZV1VVyRsQaWN0co
Sg0UWII0N+zp76FYWPa8zsyGO6+0L69VTl/n0stPI+KBKjuca4YcSvz5939VL0AH
GwiRkodANmBxA+YJY+6sWqDyBMOzkrz7+5VMM5748KQw2JG7GlGPjPEndmwhCHWC
oEV/UJKsTe8qDhJ74UzrqkogYLN3Eao8qtQTSphqy63WRC37sFfgv4sM7ORHeoif
xea2QCMWq2Vpya8CRs7bD25s4ttj/2zROrpnJ3jp/TJlqrz9UpoCdNKgAlWKbCab
drDx8gzrTGoVpw8Y0QYeo7z8EavIMrP5K71JT0pfdTAnvffkNKjblxyGv8oHVEZO
TkQxsC1fuQpX4yQEi+3n91PeUB9SX8sQm61raHq+DbD45ThyHMQccZBt3FpjskeE
jsi0FU3IuqvPclbt+uojk0tYb3Wy2wDS5shXfCQ64Ki+XcH+o0Rc2n9l/1jWLGAj
mc3v5L6iNxFVF+crZWvAeBDrzJdHUALG0hgGTRf74XduGDO+Cj7LluxSfbCKllqO
HtiySYUnLAct8tJ0pkAbRNcgYUDNZIEevT/4e/Tr0jUWuNQkAZBuLqAh3DxLJj9/
GjErL/aQtfuveCrA6SjnUAEkq09ShUDBkwk76E8i6Lf10PQPoIK/OsxK2w6sub1d
qTVIBkNMc1bHtuyXa+RuHiMPWnb8kVwPTEnoytMT49pI/rgdfMwkrVrs/qklJZ0D
QZ9ziNa0175PCDFJMCf56hMwDbsZPWXn+8QJcS3l0xnStsm8i/UjoXwswOh39Vbs
JpIPoDH19QnyAIYMjoiTUfu69dE2//Rx4Xtcb5WFmRazEv1C4y7kR6Dy/gHYUq7O
4YdNKtKfQv5l1UczXAXY+lAtPBscCttlUk4YNdbo4WluqentnYyesnQgIQhwK7aH
1C0/+6d3tk9x9PCkRy8SY+aZqIkRzB22XbrRmXRnxVAVfB/ENtrGjOL9twDJAkMh
KtUd/A735nX2xoa8jlnDMsad4naSY5yhoKyaBXKJp9b8F6dYLWbTIVY3O7tlK+CT
f3L+v8WO70RHZCn9jP1bgtL2mDhdw9EX85yoeEkgKGQ1yhUtzpfIjWlHmpCdwhvg
n5S0vHn0DpqANzLoJ4nHdxI6n7WsaagFRnzogah6RQ/SRXq5esmHK+kE0yuNmUzk
fHTGpT0FI9PiVfQq9oX6ZZrMp7iAHCVipa2buva5JJ8qQzlATmzqN84SEU01Zhis
IiuhJ1s8wEi+j14m9yYVIXzbfvvqGv2u0yEl1NSkoB+xl6yq3/5QAc+WWzUkcVW1
rTWOxUMDbXp49eqfPWpKetTPGF6WyDeX1Tl+nBeGzTogEQQ6r4xlrSJRYqNwqx7d
e5+445fkRkPQTo8xRBEJm/O5XKt/0yXDwK8ATphCNBC2IzRK3KH7g4Of8KwR3y1b
T0HLaL4iLnqhyfBGEKm3kP4/4RHuB61OdrGuN2I/4HMtRwj8QDrCzPCuSebDSQfE
Uo4Ewhs9YNCk2hjZw/lfNsllQo49kDWBoayaJHTCAb7aYk16E0wyMK2AO2cKR4Zn
+GVz2zEAGzLug5X5oFIxbSpfZgueM9hrCy8E1A3q+3Zb4AdUfqEmDHzfUibKireZ
T7mT/cupLV/qt/WoJknEFTzXVv3rsuiJ/+XniG3aVxYh1xYGAaeWZ4b0E9jT3N6Y
hOXvcdvQOcWsAmieI/V1uj9zEN0iPkAjg0OmGC3tE7XhbXP01TMx9XSUeMpU6V4L
Rhw9utPL4dShl+GU/iTsfv+8Kq5/j5sUwbckdr2t/lVV2Pyt8KSL5++daiszv0Pi
HQ9ZH/nsPmkGobg8X7P+ttkhjD7Dtw2bjQvj6nSo7X8hyI3+/owo6wtIdP2Hs4lz
BmFfMWxz/BQ6yfku+o9QbqhEIBX+nG/bflMz771fEd/4IKw8i9NSyPwlJHdv0YyO
d53gbFur3tlYHxhW0/EbIAkSjsPrFddyYCr4vCd8U0UCgS78r3A/1qjz12+4+qXs
UXifCPVrdP61Xg2UZQDfYQgjV/O2UqemT7xeM/ZNzE9PEXSt4P09hAQuquAYtPSs
ZoHGUSUN6S+WucIhCQGPwiUsrnaV9Pd0cQzGcesnf03nyip+2iAescmgkiaewgP4
ZQhIyP1m3ki7sA25l7tPurwi6on+fIW/9c44vFsJQnaJkPa7OGABecpQq3QNyNIq
5o8Qmg2A3tOHQZ4niMNUUioV5lZtUFrFuMo3MXheJIn5flDFDBQQtIoMhMKK+Iou
FDEkKjwkz1pBMuvZIFqCEAb8SRVUvVEZ44FMpZAcz+HsuyNbk5pUdx0GJoucMGoo
tUPZBhiHlPMpdVYhbwwuk1bFIXb2O9/WVITDoUIX03z/qnricbiGfq0dn0YDpmFo
lLG6Pv+WfI+2hKI97LKDJs9bcJa0hFkEArpuWAOR2KtYi3T1IuM6ajuD6M+IMcNB
Rl63vWAYeAwwzku5gqjqjiU8NZudjMA/rAEektuZbp4k1vyV/XCcGCmwp/JZgA++
rqWTUXr77OQ3oaHl5BHsGY3+ppwMIHozo1ZWlTDaYuUQukWdlhrBZtn6MwoN9a7x
XM5eJxmZwiaqIwCzNtmVzlxYDqAsghgwUdR5CSrXN2WPvDdc3PoEfWcx0lac0iTT
IuBurSIggPG9AivCkyy0OhSRkE/sj13f0/hMUdPSHeuXRZv1U/ZghQK9KcpVB8w9
0a4XqbP/n0SPb1PFnczWsYuJNikTgRCbQZlwDZWmcIotHBIZV4QM3xlr8TknKjDV
FVI6M79QrB9mEVYSWp5yATeThGUQthVMo1G4zsF48xl2436J/pDCVfpVU9RIdUsR
1XX+YG0FsHtTksETibB84CNYA+OgaeJVEDnnLUnbk1XKgLwsswFECptvdsPmSqF1
jbAPBTjZsXodQHuhN4af7IMVu4SnlD7Y6B3x5rtOwBeYR/YBtzLCPej8UCF7tnsk
CaROi28nq6ZQAZsmPINqp512+1o4X6gDY+dddGkOW/FSumFi8MTwN1hpXeoArIIL
uRQEYJEVqP2SREqILFvj0VqrQNYm+md/slUk4vTpnGu4eBryMCmLWU9OJmeczlLb
Odc2BgJEB3t/JqgqAwRIbX25dXodCoxio6aMXau2jO3ae1udofziWAKVCZh+8EwC
jxVzfQ0E4WgcRakP8ytAvQDMBjI7XkoO6+c5AHDd9yHunGHjkH64ZPOhE/a6971Y
Po7QT7hP/XWyX06UocyM5EJY7tDQN375hXHlUEFFTyCanDZPOzjXkBqTDEk5K3rF
h/dtFHu996HqUD1JCPsql3TmAs+cmkw+D4ZliN+Hp0x798FZxyShKG+gwijN5b81
LtdFU3qhQr50s2NOq0CaNlKOPKsupnjEZV8hWhtayzVdJPaD1nroT1ZKrfxGtleD
ZwKff9K9Yv92Np1enG1kTk531OO45pMeecEpxNnpQ4+D615u+Dk3YlifDwXBjT6P
quPtkTdop6nzHhXe769V5HLPxz1uHu6v/kYDFtcYdA57kIiGpaHGE9m/S/5VmN33
2U/z0d8Wp7Jr5Qcjdoz8g1LkrCKfi5HGmAYF25kAO0cqSLQQllZ4FKPu86PAMTMr
tfw1HPdGjvOa75q4nBskhGz6Dkx40IdhT1gMhxasnMbj3N2otQ73EWexTUhve6Gt
RXmIkjePRw2xQrehbKtU7fsA0RiJUNvi2prcnetw4nZdNOJScyjmKBxwIc8vqkCX
IIJM7cW+CW9KIte//FDiSq+6q2uuEbeqiF9aPmglNNWxtLxLmY5r9DX2C9qobfZx
pTaixaf+TcpfvrAgR6FUB1ngtIWZdXTm+0tKPoqnU9b90SlOtSXNMQK9n5WgNC80
JZbHkpiuqdPb0xPoyiv7PXhNhSUU29vtFagSV5V6iQxjMtps2TGrc+Rxbs8FqTkW
QsRGa549rWtPAzeFlil+3T8wICtKI6gp5uEyO7I6aggDGGLKg1WzTB28IrpQ4a29
ll63VJtJpSNDzJmrPg+pxBTgTLH3Drjve3GqZzh/enoBR/iRFvumI1J6Kqh1S9gO
HIeg9YTgUKZ9U4Zy/jOeMK8b/TvWsxeWuetA34Fo3ki4JFGUX3zIIrg926lesoDP
ejVPptyn3+lIlXnL6FlLltGYchTGZ7wrwUT8nhXKLE5MOzkqI9NnplnoOFHv/Yua
PU19AHbDkB/QprZOqiQcNYbmPnnfIDs+C8dKXMLmD55NaIQ12pPPZaddpAFaQr7A
BrDEuDorJ8EyrOdjC5XKwoQXw7l+NJtmzeVhpZGdy83YZ0DD0AjWkA9iZxovoewQ
Bt0xOIULtcRA/gMbwY8nFdLsvTzxM3PH5bVL8YhnHaMwtKUfzR7k3tii946arffx
QxbZxNmzHh9xCEPRk1lqLezET7lSyTbnEW0AQCD5pj1chMlY4BeyhIUCC2j8djRM
apsefhZWCfn3+2HaQe1qJ8bPtxz3/L+tqz6HRmmJMlK6X8iIEq+yUngKWg8y3d8g
1XQbudej0Y60P3x5Zukh+s2I6cckhq25vtjFGzmn9GlPddoxvDyw/03NKVlPS3e5
jBGr6QVjdoIYA4OV6Mi0MuFHsygZp8vWafiA3TV7+TvjkIsgsPJlWGbtYh8UfdHd
l+iwc5tsV+nyLzbaBO8AGZ1jS7TBa0lGs9e/JVwKG8oJxrEFTJjJHSQhg6cG0VOE
cPH2Ybd7NxvDL9iPjRooB+w0yYiM3bd0zQACqXP4YU7LlxLdf4J/O/dU7wEQzHdO
C4F6gbrwCuZqWEHHCY6m0RtX/9Sglg+q2gYXqve2Gfa2pcg1vArpy1uky5w5S1pY
1G+DJQBqPPkF85CWCy1De+CawpP04aOHfd8Qqf6lAwszyr97wq493PgtBoFAaOD5
uZxsOe8Hr8lDfTulgcI59pUnHq/41ziM6eH6LQVlFzPwvJhawfHsmm701Tfe0LDa
WZqHM8ZSJ3HYS/v97GmDlIaG58q9yISjZPLG4XU6DFxrvWa6ZvU/uXF5Pfzi8YYO
pS5uKtHEmvZzAY9Z0DX/f/0k5V5wZgfEm6yYNCY2LYmfKDJRgcDoe1VKIVONlcHb
jkp84mM0H4VELE5Qtq3omTPsEcD3/H0xhGgk0UciCSGFKHV3TCp7N1lQHLkCV+Co
ucKiu73becRrh0P3zd+HstN2Aa2beIEzDyWkOvfmDOumE6MGACUPOqCjby6LOx0I
049rQPmJe1lCCAcpvJGbJ+16fwI7cTWSe+FdqVsp9AM4IrnnFFr33XQubZUcPiaC
Z4BuxGhNCBJwvHhs8wyEi/ML/v4DR5s1e4YQlqULFNBKQ8t/BQPQn5LBToX106cX
yEBmvOIaoQerZ5CsABmg9CwBKW1IxU3saaEaZxSCa82u2tUNi9wCIuBlH/IQzFHE
JpCvT1JqWFrHen9dE1eO0+uzbjXSsQxSzqsEvTO4ZqCtJ6aE+L/Aq9WFUsbfftDj
Q0IPUGRxR09Uy9uyokuBLfgS9YKB+0olwpaInbaep0sHDdk/GyeNPutT8Zuk2oTd
MrZkWwXYwB+WHzTQRxSKfeXe5GD6xQ26mGp3pA0gnQ61VvUZItR5SdZnCOEZHid1
ZqjnT05X6q7kfcAG0jVtcTE8ET1dGeHft0hhvc2wLD9OHVaymW9tv342HaV7pedA
vxMOLK1P+7EW/GyZz/EN+arG4u2+21N2BcSDk06ZTWJbfV7aa+z6ufeyMI6HZx2/
pvsWJcMV/AtqRbEkGh2de+bYOxuZRKo1KenBdr7xPQFOCQD6TvNL1VIl95m/GyKN
us4keXJIcFXRpSbKKYlSHf0Zt+Ub+nBfs8sA+TK87rSdVUYtbOS3lpmgq/6TkYLn
yqUgpz2C6NRsKB7Jh73YLHH3Z9qyTUgR82Uvl+aRhG4xYuIvjGLx4YZ4XDEoyJIO
oZ9M7VrIB906fFKvBQ3shmEWuSjRocbwE1igyPlPePer4JkEHmLN9WOPS1/w0RMW
2m3VJBFnS9RvkOn6ERuuS+n8ijOQvYpr02wrLC3HeSh20WJWTHNNlTpePBYRgcH4
9FxSNr04Mk63VaQilZjzR0Q0XGH9LqrGgunTnWsaIVFcerjCeXs3s6Uh36OM6wgA
Q05H1uhF09gyxiG9CtSvuvgrpsh6MkWHy61SfQq9QoqLIFXt7lsphC1WpRz0sPis
2CvDwsctr7/Qr6MjuKtA0/PsPMWbB8Eyc5bfXmkALykKpD1YW+a8uPR8+wjJjDjK
6T7fB7pzbndp4SQmMSGZ3R+2jZPgiPELpBHo3xWnovRKSUdqzqxtMmY+WESUglcc
pNNMrcpIP2eWu2bMD872w3+kmXmySrrTJnJVBpGB7bKGSVAyAfrTd+MgD69wgFfB
Z0pWjHyrrBKJ9cUaSu3dU3LSyRnFy5TRICHuoGHKQR61O2gaJqfAQAWNZ2X6SBeC
hsB7JpAnJAyJBpiK+3MsfuJZu72LfoetFWDMmYOb060WDme3SNt+UO3vehzj1pzS
FCfknXHM6i7zgs+Gqqa7RtHBesSTrLyHbfuj8H+8ELHJRcrDtVEJE8V94ErBF+Hg
OJDtXbX7fzskfCagnxgBbKOQ0EQQXFHOb1/yEIF2CnnAmb1RVnZ9W9n/w/qbyecC
t4jbwFqJC2LNeI8GW5kDJ+Jv84wwjfH5GShcge9IL2wvcK/q0J5gjnnSbmhvuzUY
5fH1VOgVWx8c0H8hamru83Kyb5I0nvgMMyTuPIzhwRwN980+nX5Q28PRCWaRun6W
bbrudhSpeaPClXwuKgXQKTXsWEpIM+/qANbMII3Uf+276FKcfNXqUSN9Jjz+CpUK
hdNmxbEriKssvL8l7fnJ33Xu9ShKRTH8lAD2UJCGeYICyLjFLfs8/X7DORGu+RZ0
wbVWeXaElD8rndxqcy/0mnWvkA8VnFq9L/B8QCRlVObzEDsn5pq0mEin0U1LpCDF
qohOFjIamNwQ0j+S0V2dOJuk67gpqj30bm2oHTj0Wa6J2a7FPTZcLwVeXaMLpEmt
jlZ7BatXh5CVCD37VnTvkN48IZw2pZ47D1yjb+1Nb+GaLxQ6bG8hT9/gmSq8JK+j
S9sZK7tY6JLQ1caFmuS43OCp8q5Um3fcbl/2YyPmWMwiES6XFxosWv2S6Q9n2K2Y
Ucrs7UGilvb0C85J+x18eI7pB1Z4NEw3VsSLGLle+K5dVrfoejKXBl0A8lQZJcIz
BshzJHK9GDPybTc0uyPfoYlG6xxoWHMCRR+sARD5lpNdYr6zwK9wyO9gt5KfSLGP
fGNAWiXSdLHdwkeQy+WypjaORD9FjiYGi4dmQzN39H1M1TSk+1IJQBRbmdjxrRmm
dWxEEbioyl75LDHnCSRQurQhfB5H/MwK/5erdQUNb9NWbttNVJpJYjv+gBdESGJV
borReBZxswcscD9OHPi4OhMnfacHQjxRiP0sHyQhErF+zxXWLOjDR8U2RpcD9uM8
xk/WbbPbzU3vwodocarWtd0Uene3Hs+TjOwVGVxa5oPZidFyeED76pz8zMSG6csN
A6siqS5Z9KGbZSHuY2JJZ/5e6thG+4xsDiL6tiGPJBqy57dXJHUM+EV21xwAIsuR
shHO86KVYXo15c2dR8ngnGDmLTS9L7SgmCOtw72NGX+lQBrw6IXwNBzA25nrP+aj
ZYU0eBv028TJJ4o0P7eoSxejr9r6bYwHT+YgehqXgzlGLQmObL490Ra23NW80ZYs
1P9MPqSnvc3/FEWx5MYX7hp/7Zf595upCVA2B31EZoOPst7L7lur5OI8EQtuX6dJ
O8GkLjDuxtQbZcb2ZWYSdoD0Bcxxrg/9rnJnquwRIlneAL8U1ksPizw6J9EgYWCZ
U7e9SQ4t+l0zlKsHtvTFUro9npAjV9WW3fY87seYBHh6beErVdZqubF01qP7EXm6
x7kXXUZzE/BPQnLsY/4QGk1wQiPlALQh8Ik7gjvPlxjhHUYwgx55+91X2SvfdByt
khAZRvc0d0Hg02BzJT0bTshU08mknMMCLLPhWoGVExNuIMXCJOBNNeCpziCHEs2M
cv0Abd/u281p2Z2BA7rhC9yRlFw5+s1qr3B+jaWq+Js5rwaOtcl/1v7OGEGZ13TK
7zrb8lnUaInFCuxhx01kojIwwu0/idJWS2bikAT8ZvDHF5nTh0U+0HIV/dkHhofD
p8Nrki86zNy6MCqZyWUPJzwWVSWulmXldrWcPdnrxC5VhSMJaPFC8CB/dTqJMlMP
ACOheKR2iiWFC05ev1bUx9/wbNB4/NlnZ4iSMNr2DOWT+RMrMYwpRz892fGOuwcj
x3OlnW0RrLPZKTbdeGZFDphy7bgx5SBriIUHPjJ72yoNMiPWYBR+YtUkt9nE9Api
jZsJQIjbNYmGJFgfgauaTUpqY4fv78Jv6l3WaoKXQGQyyi7tNO834pamViLYaHCb
mcGmnSFGhgNImEdZOCKRB+AZkOdNt3QzBITG7knlfJxXa6FYorpTGZbItggxlVnh
oPVzOgWCG5nzgIrMRXW+35vYxjNbm5zXclfANilDAERK0ODP4XW66P2wL8sLpX+8
m9eppSL/0mEWVuL26EJ+43WzKqPwbKZfKq+MabNWAkYIZP14cWRgjVmMcHn99wKp
efleul5jeugIg+IvDrkMg5YWAlc1u4N2o5VIs9tQ5uQEZToZpRc8n89vdbXiekHc
kxj5TLQbXz5vReNaQnpDTQ4joSSNl/Z6DHv70crK6bvthX+nwbhOY0axjLwS03bY
u49CbKZTNCLKS1DvkkCVjVmwFfvMCUT09jbRXqWqqUiD3aoY1kXSk4BhTkL4Wwmr
xI6PYKZDHxDq4U8xi0/l5dSFG+wx9/Eli0s8/j7aM16DFyMB4VgN2YMqK20t4QS7
f8MmYgo9b0r0/OlXJQmhDkCqq/Y/pzvVrKVAl1musNfnVSJyTWqUXuae73eYwrs/
7/EpomEAT5s6xJsoN4ZH8VDWosBc3XcLjvEA0GQMnuDSqQy39ZOraI0xFnqs02m1
SZggZhAaFsxPxzaHDFO5QJWYi/LYnueKsvJAuItWYadj0+K2PliRYyml11HyUBrJ
C/EGcYBTqcou8ptiLcHmPtoXUCOxxEK2vJ7FKKv19O/W+G9wfU2/WCn8sMu0ALrI
1l6+E+NiR7unbPYgFpRTVkGigse3JiKvJhEecktWyYRm/okGCk2l3kWk9+I+9yYO
JIR2YGFhs0TgZec4LEKRxkeJbBD1aL6F63dM6LuFsWjhrJFqj7FGd68aYlf3omys
pJibcEnQKjuno/PMvFnYdNW8O5FTGW6OVih4u5wZWs/TKCSVdVAeWOw4wTCjEroB
Ut4U9pdElBLgeoP06nKEox2aL3YFwRhOVPw47lqH8eiFCRU5c6u6RwuO1f3viwAK
kfko96HhdFo/OnAI6GIiRtrhJzZNe3zAf62zzG3JDdDK8g7K5WhVNLFf80cuSdO0
H60a3nrveZde9nYYJr/bEafjxVFJNnEb6pl+EqcoDxQt47uJ5+yBBaXsD6+bfkK3
iDjfrnPlHROJAhphW+h3gwVTuxta2uzL+8CbWXnsMqe39TcZJFefMQOfOOoi2IRF
KrowQRA8/Ugb6+2cYwGw8Mf+jEQBZtLcQzZA+MXbKRh/ijSzWA887YyIN2fEVkQe
p9v0i9Op3E5pSoVy9yx01Wtr/IyVzcli5m0oZf4HAKgAAv6COEtxeCjGocNg2jCw
wt2ZhnOq/HMIRLWQW2ZdzrD8T4YeCjNgL5W6Rw576uIy+R1pmiEzrM7TjqfJYiR7
GEHlvj4lHpvtz1AqDMXC6Xo62DUq/oyu2PminS2QXSe89aP9v6SaXGMoqzXK/dBy
XwWfBKErSFaKJNIh8D//jRusalZZ4/NPm9pf0InLPf3JExNKkI/tvPX3qX155qcL
por7kKqpsMMEu9iw2IrZzeJnByVjLtnMUONlvHlv+RzUw5cgPE/O6Bus8pZepfsX
n3bxU0dTt8Yr3h0YvTVwSBgXITKnkq8tTyt+hrAuW+XM5+vK3wrLUALMkHiGS1zy
C2m/0D7aET+lfBq4/e1JLkYJ6amhvmihacLbd5iCVgHwaOjHsn3ZVv6EX3rwtQNu
lKuPsDgM97uwM7dXYC8Q3UeEC3kpq5YpCdYqY6hc7/0YssRrqzZM76e++p4fPWy4
4U+3+9U9TtQ99vUhebPQ4+2S4HSV6ZA4laKN0wFhVMSCDg+JsuYpeuPIdNISTz/L
f+ey8jGFzzUgR6ofpW03+V0ADr8OGx9AF68QNDCotyT0bUNiIzMd8qlspdpedpUC
r0LR3G2l/c5IRCYtA8S9zSf8uzCCFa4qyet1t9c2pNielpsSv32aBXJJEeIUbJcg
J1ZHDF14gxbiBHwD/q+NX/2NG0Q4jxqN9EhwkqAW4j2xJAEnHPRP28GAGrqb/J37
t/MJySPrYkLhh0inwrgn38Vdhj48rHDtKvSHp2vOSBUK2ZorImoQDC5HWmR0sfnR
e6SIPGwUcH9HNcYHjWw0vhlZe5EQH2PFlCK3RWvBgt74FkQYsfvDMEs5EvNLLxhk
k8aIlgqd6HXEatJlDQBuehT3+nWx/d7fGWIpmZhcTbhq5u7uKX6H7U7+Z0NKC3kw
qOHY1F2JWSjSNi7Q+pRLzmojlmgAaL0Vb/I/7W7BuNU+wZwf7Tuhd38zN/ojzIP6
ldHJ+tdWBy7+US6xpSfh1mk6a7Nfdgwp45ZvRvtS8ALLISjg/DWWcPn4CvL8u6Ru
hV+znxSHtPtXVd6OUqOx4jfQW7Gmm34Zg+QJ0U2pIRWKraj4WqeHdmi85EbkLcOO
Le8oNlPyUXek+hOelB9MS6HaHLy369r28zZDx5vKymAZ/ivDcMCsJ48hzz68MV5X
jwuXcqzueNQv7yiIAFd0XfSSHLu3tpJPB7Ys2akPMPHvMtBs7fFm+C9UyXhqS0JC
mIe2/q0Q5+ahDW+tvW4Z+gpVVmu5bqplRaQwYF8kocaxQBmgDqyIzTh0/0/qnYHD
hAMIv2b4QYFNKC7Ch7eskHqBFuiCeBfj/eLHMtSz4VONXL/hja8kMIMwfmIDkfd9
fQoc6eI8rV53N8NEzQYrng/WW7NEKuix4V5xcyZWHhsaRWzg6xX6hhhIoXbITE35
5DtLIOuhbVrdBGQBaJXODT7NAYb2BTD8F1wBbkSUTQ8N1oJA5A2ddFW/YCUgVH21
z39n1yUzWzkZ3nwuP+oVdOcD6Bd/cVr/URiain9ON9jjVLEC2HRnEH557PtBsB/B
0celW1Kq332u2IqtBE1MS1Q2045sWryU72WoRwPflt091nWvqjU0eSfYRhMyW7+3
ywY0127Os92DzPDQRKWthwDWmmB6nnnplNEjKPHcof4Bijjrb4wYHOaA2uZtb9AI
llHMK8HiHd/s9IDUH6JSNlxp7AI2/z98j+DbGtk3W4xDqgdvuzdTW5xxckj7eD6w
vB6PcTQrKQKmmlKzCnWmC5likqdPuyWGzAgwTP09nWA3nWQkGzMCQVTpRNxW9rW+
yTIp1Ma5d+Y66Tc4N0SVd9kDe1oLWA7DBxcXp13Jus4sMZTIs3eA0cjF+jarhszK
nUO/R0iSGJ6SfPK+x4rQXXyXAo/qCGOxJpU3H600ZUO6dYm3qhx33EIfhnO02Aca
VYQhusxEKysGBs5Lq2JOH0xBpjxEeb+XVmODO77hWYPY6y8HeW6N599bRg254hNz
k6pzwCgodVTtVakNTmZ6CMHWOclsY/8I6Mptly9fk6xydpTf1n4FY+lczelwwGRw
3TiIboJVBftMltpo0zmqFMkH7DYdRPpN4QK3n04HygSFqZY6jFPK+lFHJOkM4suR
nuPeD8bas8h7iX3nPylPUK0ZldfE9FN51mUMpAnjinE/cmBagpDMkdvOZwdmcUW5
F8+aP24Ti7xqH2wLi/pPwLdf9B5K6TxIVxE66S6svXdJ/lirVP6gu51h0Lvi6lIC
OscPO6Aw0GEAPeVhBD/ZlNbuUX4gGitOG68b0ZCjlv2F+8wFIYYKlfKdGaNDJ6AH
/giteRV0wCUeJ1FzUUyKHUasr94LKrIMJK6yf8BxlNZNGCKDUCUnTT3LFG2d7KbM
ZFqwX+4zN64jm3+p0OfzAQ1OlxF3Mm8QsoWVS4Sn1eTDtvJhiTMrg5ULMl0IGF1R
zNbbk94BIA+OzwFCQ12JFnTxADqGtCULixC/1fLAe7i5qs/3D+kC+G3QYfQQ8028
GktqTv639z1LoQa+4A3e2b1wBNnce525vDZQGxraou0qO6ajIOL+xudckgJn29oH
uVndBJgfnrSjvaJCO4jWOCYCCCi1tBi22cr0E+zEYPe0JT60dXIo2CqpycoobHXZ
kH1EAOMScVBkg9c1LvMyKg4n2xS8EEEh5JwizveKL0QWVYviFh8RCwmqOiEy+zSV
MocPtBilu8kjLSLye70agIMXrQbuZCvpNoij5Kt6RfUqEN1ypfV/mL37SWXF7CvN
Oe3f4lDNp8CLXQAwfa1C9TR05csiIcKj+/Sm/p1660duUpD3SXOVwQlYg3BxU3Hw
cV9vSqerUr8XMJp8lnwH1qkze4G8qVHL0Fi2IHahaPPetiUqWNUS3CkbRdUkklN7
qpSbhV+DWYr+NbMpA7u3A0gouGiLdk0un0YU6K6hGP/MazjDzwshaj1cmrs7zSw9
rwbuJKhH/ZwSPe/uLvUpuK/v/8Wquveb5Rvvq8dZE9SFeWbqDMvJkI7d9JUtdH2u
QpjeviGMl0mtfgvkIz/eerkZ3jcrsjDNV/8ddIT6v9zxNHdI1RbHtKRecXlZryFj
lNCgQK8EtzepEtpuc45Oi2NfDVPbdI+z6oCwMOsEmjplzby83DmgCLB2yRpDi9jF
Kdu5nvqRhwxTcTAF2v9cf8xO8a7Q6UG71UYRTAnELgzlXCe3Is9jLljG9adZNi97
JtoVrqCOk17MdFLiyjFhgK7Wbqfl2lmbss4jTzJwqLQUTox942hTSDenbPineCcK
KGKHVFCOxQEP0sbRXqxzgpWm93vGWW0XwRxdLauQ0DKiAunIUPHeJSYK7hilg3On
glkKqUZwUY3XVck7tfFBzPzjICn4XyySWmLfhJDG/YEojHUMaUjiCOYNgVO3UD2T
w9+ras9PkG30Lj1wWAJ62mxiKLyUnex8tUY8KDyYP7+4BGP4Zy42OBWqrUyshLlK
qnSshAvOSEQGqx5s35BMBmmBX9ut3XZz14JkrAJHBIAvfxRQBWzYMrrlzJaY0jCX
/8nmMOFDSAAMNhvc7j8lj5Tnll6YOQY6Osvky3F17YJw8JDEfmjw590yBN6Ko0YA
CVxqnkkaNtkTZzc9r1RpBgstWE3tZSbl4gd76gii8I1kmrE8gMUS6lJfDoN5RGRy
99fdt/5c8+IFydgoRyiL3Uuc7kQeSR4hQ929OrP0/HGunGg2031BJThnjmxSeeEB
Cxss+5tldsS8wYUBks7lqVQ4yL3F4Ra/LVQtbBDb9Fwiu9Oz8lsMyL9AUvWADsyg
V/5iF/jWDDnVRq+Zjm3ppBbQMa9lsz7jUnbSOtoDbRrtNu9jwetykLkv5XhMqXF9
YtsvEBkk4yHZE1yhNPuoyDYTQpR7YXkQZDBOUvQIzCHSCKCJPP0gzv6qW5ZdkN27
UF5lFyVTG0Hug+bUO2qhQmzRouvcZoUrwShEuPlhXwGb4QqLN2j3ORrEyQcAg1nJ
+pAjOeyA49tMrWztiGxtzN3bipYPdEXbYoE8UfmoJ/UH0jCLmploqqnC0kUm2kow
LKmLVnMJFunsDJ4A7ZcVr4rAU2hSYh77wP3gRia9LbA4tL6vzNt6xuLzvVglE+DW
hRL5SaYrrjqo7yGBHO76jCP+wRnMvpVEe+gmiukDrG0HcKfKF7OjIHuev3QyST59
hUTqCsvm2kYudLYpPqaT3yWizoAYillPzDMwJdteDuaQ8QMaSmvLyQQs3/ojxfRb
mhDBxcqCQppZ9FrSzFY5yPX06vpIMeEF+JPYwbc+UvNyU6Yvz62p2Sh0rr0Q/vev
ug5kPbGQGoUm+Prkgqg+0xJLkbRZL/ZwNA1ejdkNUu126hhiBW8/nLfQSRnrOhV6
ROHHMoXpigdNhxxLLseD+PdRF0YaZFYrGKc0SA5fs3dWi9Hx4T9HnmlvBAI33rjs
ToTGJfoBRybJCDl5ajJ/vCMN9Q2FJGRzvrGbCeoncEKxD8alRa6hDlzisTzgS6IM
8KRb20XEJjazVU8WX9pTXRyNCRFhbb8ITjbn/oWv6iFOSVUnrTDAeNz7QT8jvLrN
kmZ/Vp5tzzS2jQwBBL5Ty+h3COr0k9nNHpynGrz5gfD3SVl8/217qzMBZLUv+Xmv
TsU9rReJ9XUVQhWjt2DwaHEyI/2zJXwG5r1vXiLT3/NCejhoY5d4pD7GBhGOotDa
8qCi1wLZWTldTRjscERi8y7Veo14OAal3eoU0feml3PYMSL1K/SfTcFSXYm7BgIY
NnIC15oKTwOKrYWc1R6viorvPRC7ycXT5+8vYdKTfM8GNArgoJe3TsG6k+1r9yVj
gjujUK1Q57eg9M6kE1iwAOoZkxNg8phaeN2T4C3r5nCinTndTbRuT6oXwZ8pdnv0
eE7Ni7VljfyWT8cWI2xXHRxi9LIv893VRPikbeMqHsDfY6WEY/TUaM5fh3++F4cS
6u69CAs5dtwwe0YgD+0EZDUUN6cDt1BM/Uu10FYN0196CcaF7qkbJjHAu82lbJa0
4XH1sMqsh0mYZ3xM63vBLE7LoWHiYAXwuDjsEEu7s7NqTZbpWMNLfqC+zzj/Brsr
Gca6M4GNv5G67xOEGDqq91Yt20MX9tnf/dIfys/78uaQaNoSFg7PfcNAfwdt4Ue3
1R/LfHNJWyrTWfdfvbs2FAyUtYhI/PQRd/dMzn3oY1vU81mZ5P+sR9ZRZTZkgDKd
PvAVeMiBA/xzxO+66Iym5dcoQDzgfkmAmX4+bUfvdxBcnE6H/9jqrQ/xrFgdziDx
eYIkr+qbbd5houQD4nAr2TH/OT13Sf+ecloAayCfKsc0An4p3XRA1wpsXG7Mtuvs
HQdO9PRqBAcDKKbxo1ZQthyN0B/LIXp5q5LjV/dzy9Udd106yOMjpbe/n3J5CVMx
yQfSVIoZfXAm4M47Uowuo9oTl0aT2I54JfqBA+Zb6bIomA7Ntdoe/57xqqvFBx/r
++uHIb6z/FSAqPOIsA9TQvy4A5psrIC5wjtNGRdYriIhOnSdWtrgQSlZq51hBBjK
bdbGdw9UQKxE6j/nA9CHO0ch8t6/r+3eqNVPJ2Pww3tEdxaCY1cYA2dyP0Kfmwp/
CYZYqiewLBdBtpa1qmRSMohwMmS42oJO/RHrk89mO+ofiiXPvEqDt9MAUZIU02Gr
1fk6N2W9VdqqxykYspQcXWsnmPuXAsjHhPfpowiVSawsL9hlen5kUxfej8Y0009I
gL5cSjreSf9vV2GlgHVjrCFvkjP7n4iML1yMO/2ELwO7W9wzKqt4kvr+X9Bn3R45
YMHOlm35WHHtFycwH1nZ5RNmoE3tYWwsoY7DUFXhyGPzf0H0J/M28x9UMX8Ph2tv
rB7o+gNUH62zJctoS/YzPBNU/r/bBSjBEpcwTH/NR1QQEdA4H5cj9djbDNz0UvrV
tWipzveN77Yo6SU4bN5x6lof0wh+wKWaJHeZaz4VSKTSWlj6m6jea556uNSVWxWo
+vHo64RfifjLJ+Uo2N7K3rjSUweC47ggh3l82EQZu0UvQrzqgT+zUco/OzbnLhDG
cm022VskHM2fSl4Zw75IUugARm5n7R6Abxej8WK5Tl7waxT6kr+vBiXkPijs2jjL
fJb8UPgaaDgug9Baoazpw3Fjzpr53EBqG2hOBgltQCptcZlXRdbnye8tcy9prSn8
8IO9gzTB6DfeQUSQI5YnBSV1DJBD3C9mMTHSeHlV35H5t7PTkIFA9uv38NJckf+y
Cqs7BYWTIIsI4b5suz/VdDRt6Eml5fR4xF9aiCZs9dmpSwu+1l9u2QjHz5QtlfLH
m6iOcSNZZw8uOF1PXNe3DMTpKN369ETDLlxE2VLOv3Eue51vqe2GEVJSjdiK4qbq
fEsL00QbsJozTA09dXZv/W4lyp2ElfW4Q/WC/Zi15g6WuN+a9vM9T/WnlBB6bJhg
FiHRfwOGyhO3Kgrr9t5NSotied+pzqBZyI7VT4/XjlotvIbRfVmLkgElnZaYt7qU
NyJEgKBqLAyBperrm011K9Lf9VDMQ55N/y05mvRBY2nsQlcMsjV6dFnmMk4USm1/
vamHNvrKIAPj9xne93FhtueNZz1TbRb2oucyQgFrU/FUFLENneeHj9Lhl8xpQAFo
8YMYxrMHrSS8SR7PtzlN9X4TXnvibuxuUCrcMf7wVGsMpmDbRVpPQX47y/IM0ro4
Y/Yg1aWP4UUbP2AUNqyDUpb4f6aZ2QZfbEANAOfBjfX963nbaQy4ybXDvHYkL8hf
M2d5RW216yU8ryC3aW9qKRZW/7R1u9mCf79Ha1OmMTvGB8EdL2gU5qORbBJ/PH45
P7x/NCMm7uXtOeWyyfDzMbN9IX2FEs/+fz3oMxK1H0kckq3fJgXEut3JkYZXhIw/
2qpnwbWQaHpKor3mtHBLfH9+SRKWco6JFrw4NDyjsLHG2uOomIjrwADbq6x74uWX
GNct40zx0vLqN9V4AoM99Up1017w+2Bp4PokeKsmw7aD1KOtWleXX9ecmhlviBgE
yfOOBRZFhA81f8xHjocNS5NYzYO4/1ahBVyCywGHu/n/LlrSqNeazUhK/osD0ugH
ZZIc5h6SLzurlU8LWmYN0QS/LOA6Q1smFO3qj8BP2zaGod8dOK5Ew2Vubn4JdUrS
7Ni1AnKOSo2IGyOffl2Q/My7OidGifhjLIHrwf1yueLtcmKUwjqBYIwJ/uXUujxi
u/TQ43ouAXA6ujaSgCLB5seYmsAuEPimrKZiLSkp3M7ipuL3fYCWXFfc09T8g+Bn
ZskPVHwe+wdzgeVL7iqUgM5T538HbUxUeMQweyTlTsbOwJXk/bDONkKwyntFYf82
AID6q9YaXJGTnRwidp/G+86kFin3JOXE4awEgdsvCZ2KDi8EarACqJHlX1iQgIHT
cSxdbyZT2xsz/iXQ3D7pTX6RFZZVF5kBKi6zCXBNdrclvSmbOuOQymlf7mW//NRu
gicVDN7t24LJHrAKSj0jfWX5M2k9pW8ozRe5WuWWzmtFp7fJckNuQAfULj0B8Jqh
8qRsFJyfbKXRfuSNWPnUr22/qGz72DQRSSaVDgbHiwu4Q9WfE+Day6etiCpcSciR
EgEmX9AGkWL0MeYSjOet6CBkCT5kAcg1iDWa2zw8E/uHNK9iyEEkXNaxzOqwH/Ed
FRbfawfhqyP3lEzDPZpO5oZeIV2VdsXun01wOX6wLLRmFkaGcPnD5ZL4MQLAv1gX
KaRqy7y3VRKZbNmDGc7huZYDuwtS1fLm5f/hKIN//TcsLMslDgDwA3aQlwDh3p/w
EMkMiFI0VGXkLqVzwzG1eGRwrC7us+Kc2fizCED7IzyGseVAvc7yQDsP/19VNSP9
tSLZ0CRr+41o6lGfQ8oPutwt6VmwiAqxB8+mlvgDXJCGutp81zWc6Y29kEos7+ZE
CKSSjW+O5Shhom8z2k9DyYH8IYE8BikBr8LKW+J315ypCi77toTHgM+GooTSnQ6w
lkZCAjmFy5dgE2lmzne+7r5iTPdANfGRjrv0plulqJRp6OrM1KSkPAB5OGR3BUlK
fv9TjNbLZdGHAIE3KoJ2iHmGRKYOMJ6Yn22tPX+XvCvySSqkcgYTnWwekMgs8OqS
dcd/hT2dX5XrFCoi143p+cPlMStwtldag6m3f8ds2zxxg5QRRIRVmelrMZugviP8
tb/MojJx3woeXPaJQsHKfa833FU5ldU5wEv9IQqWmtM4TIniJ3yyEU7Sj6LMZ+3z
Si5g0337KbtZijVOXEBvKlwSeccemb0WSTZcezg9hLmoop5wF1hciQnvhh1ZSXf3
/+hmKw+Aocuh9QCE3jxldw/2tYGslTbzzikV9uVkzYTnR7RRsoh5dAELPAvQDqrs
F6thZw6S5tY0EvT3D8CUAIROUAecd3TltjKBQa1rHO3MN48NrLVyIZcajX/IruNd
l9IQwMJNb8sGG8AHjcYi2sNZ+EcFY38xf18URGYZIi1oHsTrn/VzO4GRrhMxHWzY
uplVG++5JjQ0Oi7LehzhNmekoIrhlkfxElwn8ndIb96rcfVTtAKAmDRi3Oh8Kye7
h1W7f8fquecyT0HoVxamqFvB5sFojY1/os5ScPpidId4ERHxeE/maFp12m4nH6cn
HcbzrZ5xlEy9XnlRx0NQYZPdITxKh3j5N2ZHwxaeiT0vax/hfT+QADXFso+WZnS3
OxdvOJ7eLCpAgyXBKr7JEh0JSwYEIHl0f9MfixseEAJ+hvKzdIYIdqlfdzXOuTH6
Yj3Oj5qUMkdie2egFxAbBAQBvaZ5mPkVKXmz2jkmCaL/ae+ExHYcHkWEV8Xm7Myy
+0uBE5AkzHiQ7wz3Z+Q4EWHRjp4udcarhNuz2p74+OCLup274m23A6MflE5PsgmK
4H6u0xUp7msXS3MxJpq7T8r4Zgvzz1Vlt/0yOBM1P0L8YG9riryf4aGR2tCGb0Ki
KYocMBKqTO64zYlSIttWHqE5i1V6UqK/OCV4D+6Z/sYx+XZRYxuFUrzt9XmRBZ99
3/vQpBQB6yRHaPjVb06LMsaTVq01kPev2rJ/rWGNneA6P8AZ3uSdEPSJD/zNHtG0
2H5reoY8aZfJMWeKopG4RJL32kx9ysuddZeQd0OjGEZg3VJcv92hunIvWIySJ771
R7EQjWgmOz+WQxNsIMulIyArXZU0nc6r7Q4eA2Dm/fULz+vHIg/+qDNg+EtDPRlB
iM9r+DhrfbAwgJL07T1p2Icp/TnXgCbzNdn6kSomROgdt7B3xVy6wp/en8o8r6i9
yVxOuE4TCdWFb2zB7Mg/Ez4wijsNiRjp7vOrWu5dxSMIvRJ1QS3OsUViWqiozNfq
2mlQyki6rCk4XY+61lJx9cOrQBoppzm6isA6JZRUJeO5m9VBQLqTdbwHqs/tndwW
gWSswe6+2jSuhmD6l4AF3QBjcooZ6CTxkX6ZiK+TgzSYAgliw6fDAOg2ZdwoYwN4
FDaq0lusBdQeqpqQ4GS5m7WjRverv2KSL3OkjEoEGjYxw+FRjjqVes7nI/o0ufez
EhrWITo+ESX2nylLq45kbKpX6wOBGyVl7/vC3PBR684zjHEjmWG346HHN8rb+AS8
3B5prUE1g8D1poMkl9ZpKpemcmCxps51ndIa0J4yI4hgGupVhhtxPQS0Sjy3GsoB
6BhHcBzlOrSq4+Sw12iUEmDh2Ja+O/RKknG3jeSWT9wgYAiP2bi3ds1LfFtLjSZT
uu33oyxGuus51S3toE7A76s6Punj4sH8aLUo+Fwl8qHWkVQO5BwjlWlUiHo3W1KN
Gm2Edqc3YQNsdtJ0PC8HNbK+JrxtskcaJ5pnSF5U8WQlVX9uPfOqVttF6TuZxRu4
9XrUhWE07UrCGdi5CdpcEYPrFiT3mZnEkcjpYdAtRCN5pv4mf/e+uUHe4ct+SMeK
Wh2rNQNUcuNDE4hjLrGv5butTzd0ohttDFU+G8he1pTBKh2q/bKLQAFK2JckO5iV
UF1TTHNxr4etWjmldgdzCb2EbcXuy8Szd6DfVpM7lc/I/L5R1Fe1NXarL5kqYwx0
T7SdnBSj1Oe97vjHv8y2z6QqP5q8Qn7ZwL/Q0DYM/ZldXWcdTn6RIr/otqVDkLuX
tYglnxrQ0wrIfY2ple1DVLM6zNi1XL51pdrVQrIK9YF23+vEnpdvfP5drlBsjFxl
M9eBl20I3gl+76rQNikQw7FkKLuAWW+G+FvzkhhJApXQsj6XlKtZJCIRm4ZkH2rf
zqhazPaoIbtId7/5ZRqpE13iCjp7iQ7FUxel2aWxgSFTJkxoM2K7D9Kl2D2kh7/k
JVpeGnb+eCqj5l4ZR2+6R0qVk+VUT1hG1s1Rr19vDpCJ7k+k5P4BWBOWdAx0JEqh
W8IX8x+5Xjp2MrIvzLondveXssoIGufqyCp59jvXU06ei/Zrhxu8jDjGipdqth24
x9vDkeRMBSdqI6v9i+AlaD31I1UW3B3jdRF3queyblnNboUdwhzAf/b696b44AZF
zgo99yr/K3NjeGyDPjapn+jKU3kpp99n6jMEJE428X79AEN4doq2yQlHIf8+IbO2
Bx0iCr+CjXNNE4KzdrCPTitMlDbIiBbCUqs+/XdaPtor1DX+k2HWkGa9ZOvJbImD
2G3FceoMfMLp5hJvTPdYmwz78QFs3bzy515FY7UiSza9/Ut7X+6CMe2fhAG2GzDw
BN/Yk8VkBnfqa4zoTX76w253W+BtMWlgrYozx/4e0IIfUektGA9yioz2osQtMhL0
3uZZf3dSNcWX3RfxECTuelbbR0MPmTafme9NSDkdbMnDEbLf3R9vTT9AVB5KLPoF
PqMzyrqiiJL55d9mXabeDLWt8pe9+eKyGeEpgepW6YBy96KmH9S965w3oNClmbDO
qbS/emoYXGIg6STvG/mzpOavdckgTgDieiz/g8+sEwQY+WHc3dz5FYE+WgvYd2+o
zEp9sCvywo8ttuBCbFDoQZQwQzSW07NFm8U7803H6iShufBWA6Rr5KWs4hfcKYq7
cNzNLhPdffJ9ErXJ0TjAAheuvSZIrjhva0ZrKwTKNuVPp2ejfV1DBPdmSo/DZFWe
n5QL1e2nMK6HYXS7IM/Y94XLb/B6brG+xcDnnywGFwvjPYye4nuCKGkAiA+/ej7l
N0FXopcg+79h9K8OIH/3Ah7H9+qarMQg7ob0MCtKFlj01AQ/aoLQZmTHjk+L25Ea
qFkGvlPS+rwxaDwAv/bLJkLF+ENq00xicT5cppDxX0EM+2/4BVv2p0RVoX+zSVO4
fOaQVZJmgHm+tFapvEDaVb0nuLBehf7eIM59Y6mTYb+wHCaX/huEdD47jkS0zJmL
cBEyEH098a4y9ZttTs+kyw7kerHA5U+jNJ/JzQTqelaaqS2xWA0zRa9k18Y9wocM
s4H/Ou2p8p7D4F2Qrcm6vkgQaDPejKeRF8Bp3wU3PHc+RhKogrM3VEwuMeQiyqfT
GYPpydBRLesViZxyn3mAa99Z3J1AU0GQLDyy7hxmQY3dOJ/zdDwoD85MZrhpFpnN
MftNT0Dug6GtS2Bg1Z/wz0ZDCSd6epjNM0bvaKECtr9RQw4KMmLzggACPCsO6VHe
1KGD9PbZGcUHbGZG6S2vtuM3NGrHFugHMg052WKacXvfFJJej0BMf3XaGFJ+QB8w
g9tbDPERm0be99VYmOvbPPCnBz3ZRJ3St0hivqV+PyNmK47QtK2JoSb7XlW3cRk/
wS4I098KcOmnQCYFNEs9yeyHxsSh3nk/AmiiLVN+3WnOM92tXBQyJTo8oADL5HTT
PLj6eOOL4eZFoOlqytWwIybZkEQoIPj5JR+4kiLVaR0trVT0p/K0jtVpAtK27eha
Foi+T4IGZu9XeBmeZCOLnVY54Q3iKlyfx0h15sNlHKqTlW5NrfDgJghUayFhLmL3
HPSklmKWdSzQPhlQ7EG61uScgB9hYOCXmUt/85z+HJdZci+vQ9O+Fcn4Sr9zJe7e
bTfgGhZHizazE7UfsixFjf1cGQYZnhxTHFaDffhfgUS+WMOiakjes3Wztw3Acetk
0MzbwOXcB/pRqC+5n1ljKESwcgokPIibnJCiCexrVVH8jIg0aybdIiD3TBpqJi6i
cTIHqwIsabaJh2CQmQVZQ/NpzsSC1e/O/2bWa3Q29/yr46oAPXsuWezFMShBpUCD
VZgRCjOxmlUJLZm3kKyB+ZoM7SOe//7iM+ydgDwR9cul60D+wNBKaPBb+vhlqwI6
3QLFS6ohFOq6hcKWHKi3YB8s0+/iiBFHhF3fidEcAvCPHUhYpsnOgSF44udrisNm
l2BsUIdToDmRxQdc9/gAdIre8ucrgdwS2Ub3fWvCPXzKJtCq9lMe1uGYn5DvG4l+
9ugcKiNrmD7g5QiA2k7/OsiDZYU9pDG2FJdS+E+gQoBMjWaBJqAArVhdcpBBpV2y
afCHUSrWIsbzwsHu8/1B39veHPeGCVbICnPmgSQuagjY4c2dKxyvYgXcm13jnuLu
WfWZhPoXnyPlFA3R2a+ivXIZU83TUu3nnJ5IpN3JeVo0zuLnRiLfX3MEMkJJgMjZ
T3+07VA1wl3SSRbPLksxwG11CdIkQezVgyAmvqfnf0zc9VT5/Dz+hO8pMRpLU7wJ
8YE8qmsiACSM9Myr7It+F8lLRIF0sY+bpUTGBqxt5h9bK9g0ZoqzEOYjawysUG8Z
iNVu79HR9JlMcfTndDHa3x78WCEoXOmRNjQdY7RJY6oe1UJ00iVaxwI17c5kpJTc
Pq6gV/hVdjfEV0d990ue5t82GvSC+qTKNfwTMWvWYjDJaZqsGqoXTPsL26Lafz74
YlBFtmpxJmwLPW2lSkODdCv2cN34OF8+M3FgTC2NgwHe+aNA5lsKIbi8JYJ9MV3+
wFa6FY9J5SJEATpAQQCM7NgJnb3UP4/y4d3FqupJcpjO+zNjwVJyMtPh01HvLtsm
Je34MJ7ETM389YfvDdOGiV1vP9GZNflodC7YHkhtrDANDHT0jqzSi9Ud4eECmS+L
Ng+wLD5jhCFFKX0rLFXLNH3PYUJnGa1h0GNpUGU+tscvBTfqp5NO5A0ZPFmFGi9N
3vNsf9Kq5PbNZcruW8hgQeA2+95ifVUs05I5qOTudu4nFdvZNvPOvMXmoBwR2+ou
rvjGK9v/6J2lz0DjD5NzhrmOoMMSvyZOmK7NkCUS3mOOTG8zdLBuFrIIIocCa3ai
CyQy7TBYk3qbVw2rQ5EUrmmDByyuf0n2O9wyF49ju7iD0kI7xxqLB1G/YF54Qxd7
RibuI8AWiQifdBg5DvLlYjD2F6ay/b0OZcXYdCsthkxv1txzB3D/uLFmt8qfhMNZ
gFem4UQGahNyWq6/zOW7PQL8P064IGW/4SpnJpfU61SHNM4z5iwSIgpCNuKRebuA
AiLtydZNkzko5kZEFfklz0dBbl00eRwNgEbwYW5kt27PrubiJyGeVorkXjJmLhAa
sX9XkLzNjSOG4woFNEpCiV39KKSkrkJOwDWsMo3r+tx/3HUNyAsoC32YZ+sLdkoM
Z0z4oTrbUFBy+uZ47Gb4pVXQH1FxozRPHakr28OYLVsiJYEYhsmVgBPam/5teF+h
wXWpIbWlqqLa94apvcVlOBqJOvT0rxv3N8VMxcI8vH2joBT48X9A58mldKgWGd41
zXgj3/3g+VLuiDmKw2fbYWDX/CnuFfW20kV50uerbbXOjEEzTitMQ68/EEdVJls1
lLidkFMkLhPnRXRc8dcV+J4PAgThwTwjsDR34G98FlHbm65DgcFNiegn0xtyIEQv
++8O3Og2LbRDhH/wp7iqjqskKVQm84wjxpH8ZW+dHytnKJWVlEFmASKWoelyRUmW
PUFo6nsSowXLrUVOPYW3loymHj3Le7y8VzMUAkPgxjPGtW70H2yEB2cT8Q0urvZ8
IWqJZLNp9vRvSAm898CcQIUzRa2xp9wRsuf+bRCfhYywHuMQqCEN5MSRhwEO5OMA
WXJ2xMxoequ/qHu5X4EVeSQ839NCMusZM5g09O7ToOxBBX3BZiGD7q3hmYJGaQWp
eiYRs+wKRbg4SC3gvqlbgnWQfFwhlLJIqE14ta8FYOOguyE1nhubCIwpeZcRd50E
tQh7w4TXQNxpisxpcWbi0MIck2RZLsIOwUs+jWIa5Zkn32chehlWi1suG/2ch3xk
XD5qtHH3mmep4TFbgG2h1OrqLbGzshyWUBG1CGhUwuSmHCyLo69damCzMTAPqS4r
j06x7OjRofhyuWUAG/bpM27H8vqHU9golw9gaH6H0R+wuk1AP7GZBl5XGKoJPMCl
qxutKIUvExtTKTEKhlRY/gQx9B4oITaHS5IJeMN9KmGC9eC+nBzfCOoytQ69bHqU
Ip5UbqT6S9/PCgJmxd87duVe+VsahuTQ434+Qvob74blR6g4LuvoySu12KIXFviZ
Iv1+vY6atg7zolsWPHZOIcA1QqdN2T2RjtucelB6YrYC6+Oh2CvS/xuICwHCH27P
LbrvaioahS+Qj6vJOPPJGcOn1dLnXXcinQWXVWr8ZmiMseIrbAL83NSoDq3xlS8b
2/NMCXWXimtaLHKl66Fc353+1yNjAC5Q9hWZDB2F6c3c/4q5Zv8uxrg7Z/E/o/EZ
d9i7vpvBWENSlqfG+J3FhBCE/kBzwCaaosYy5lmWq4P1LPqjCDJMN4xhJUKMV9x/
lNCQpYr03KhlK2x3JIOQlvfOHhySKGXvykN9BVQlHMKqndLxQNb51RjBzlo7mLfn
COb/LfUoCXCAlT/d2JvooiEIKUccBA6sB1ovDG0kjLs671LhMwSdbWm5HGcfSykc
SDU0iudkb1Opi/XNF21/k/8j7zjZx0+6lFpV29MLzupsKTGaeQKoI6BKQQV1/X4v
NaI97309utPYcAmXwN+L0MckucGxjk6NqXLChNZhqkIJKm53DntNbnmQDznIggLw
WnmSLY9l79C+bTdt0IJB/FUOUObiMbsvqhwd6xh2Efw7sPJb1yQCY6RdgNGIdsS0
/Y2Ubl2MJTZ51UhTOSsZ8tBbF9sauSLlOxyqtdYH/g4uDUra49WPTvN8OWY0r+fw
I1fDUieBwz9UvIKAR4RV5ddlBCG91h6j+N6iUx/EPZZ25ERt/8U3psITocQT2dO+
/wnlyl2JxYMdVSawWEJqOSf7F0Aori4mUP42yTVUPYDRvbUvnUQCcJUGKsBeXWLH
SGmqOt6oMOr3hfdUZ0NZ4KR8GhJoXZagi4VIg6hBOpVtg8gbuXWNJO/ZCtN/xHP3
QHs960qE9lI6m1GXjwgWSTi+5HtjVMOAiKpBn44uDPyWp74JhBaCGRjV9vyetiga
OQmtqeR/4/kptLnyx/dIQQrUrB1NkY8zW/WsroaX3J2ZmDr9B0L1z+cxoR3QiF5i
xshwOEY6pzhjeQksagNvWBV0KnyD8cn3ZXSLE1GTD/SrqhQZvJpLlSgQ+Eiui4Py
9/1iRxZO+F35vdB72iTOHqjEkXZFP5kyWFs6yhqiEANTcY2rCZVanDq5klVDcSH5
et1SiYqGD8dtYr+7O5Hsa4Tt0f8PSefAjfGamKWdJuPTlORow8jlN7SJ4Q/0XEgW
1kocvn+BQcw+25DEEESIj4uMBvn+Ft7Rxnm09AkMbg6nHTLDfytnUuAhcqeo3PJK
RhSP1DPVW8Jo1KlNouJKLVTOoc3bZumk6Pjb/fPUmJxrEIQNQirTPKnBu8Qsy797
ItiMRzMQRr1EcPo25U//vvdDjP23jw+SOS3xg9j9h1Yk1UbfflHB3uDh4fLbYMhH
NkobO//HhmkeiGGVr3G4enkaY3bGFLIbRFtoC9tpi7GmCtafwgRKmb2wBtx6WxJX
er0zVn2fsR7I1FcxwrIS4gQVPRFOgF8wiHe+DYVuYjofbsVz9bCR3jcK+O1WAcOw
rNmiDtgO8sZbhJPlLJO6g0mKbEFI9qgD9f3DA/SdXnBO7fm1P0l6IE/X3i9YDtcg
2Awu5go+B7d6ovoDk4NqidX16CUoEvOgbe8z43Wy6ABBRklWocF27ChsL08+997k
8xJjcl5EMbXz7aZIKuSr8NY8ReRHGYISk0gNcHKLdQI11d+ZEsPlYKj2XhNrIXA7
+0oZF95HJKwW31yUQO8Qnjf0LWpSZxxL/NHiYG8zmFukKC8/44b9Y0SGiPDSQ/Of
NG9Z+dXzcH7AKOZPh0QwlbBgjdf59YYLDHKeilmKAwenXsrLaw+L7Mc6lQzdk8Ak
hKFTEoDXPnmGeaYyRrLSzhlf/EB6iXy0u4Qtf3Ker6ZGSPKZPAcSw+q0SeoSed/q
7rU/cZJMapPySXQ4O6vUAUiaGSzu9dQty5I+EXOnnMsuc87w7JLuGWx87FC7GGBO
FLpkJj1G0ES8y5vAd1LgXxrz3tAXt12fDzQddmJXxuBU4VYbJeMT7in+yvrcva9a
7Gb3gvccTKY9AwKVqy9Ej/h5IjwtyaLtooNwIdkK48LUpkgMTP50QWvscXRHjIWJ
11WEXAst5v50s7myrDEl9lb/PypvSVE5fnnE7kdSSoSm+Qux7bpHhsxlZJIsIKnE
31hl9HBYMEKZPVmwvp14a2j9TL3p3TMJY9Z4MSmjrzDWldYogeBYUnPlaO7nRJeV
k1QkPq5nfQECZlV2Y6f1D2kCXRLioyqKTf8rRjDZh+zGnwWmKmTeV4XjDg3IaVVF
03FhNXCNWwWW14uSHhDkmi5axE68AQFu+e9ZDUaPSptc46z0oeoZOI3m5CnHHmhv
bLRnGTu4UWELzxIgTPK4ecM9CTRmra24lSFgwKbSyyQDbF+cSRrn5OymMGxRc2O+
0BknLS94KzHaLZBS35QUZHVaFij+85WSbzSH/l02nTHkAK1XzT8DYu2sLVZfZOEz
ihLMISm3OXbgQTGR941XzCGFBtfPOYFNYHB3RluK1d/Cx8KVN6K2DE7p+hif5/AC
EnZQrQJXQg9XoqkGDfb2CXugBD6mizQ/oECkBAL5/uWzbIZVIHuZpaV1xc1qF44q
riAUaB6dhgEn02FDrTPxYm/yoB9VY61STWTpGB6FfVZ3h5q/0HoeribZwXZBYAns
deOQRN1lX3Xn+c6hghnBOpvwVRzqIDAQPNQIJyMLaOzm4tJ7YYMTrSJpWjGltYvR
rwRrTiYtdE3NMLMOL9CxLmC3yqv4hVctahEW+ZXfmJkJA6D6vssHAXN4DQPDNnCz
U/BEs/nIw3MAA+/HZPLfb/5KKt7SQBIZmN7oiqlaqEGoDJ0/Ec2HxrxdAw08f4XZ
wFKHr1mOLu03vCP32DNaUw3EzWEQiQTaK9269WvWbOdyKMUgKl7lyO6O+V2hIS+M
bWThPQL8wqG8q7cgaX2LRr+gkK6j7ovGirGoYAHuSK8mE2PP8JCs3nGEP+BG/8i5
yhcjeLng1m0nv8YpDNzKPIIoB1lioYbDesrKLSRnxCYTmNWpgIdzAHd6BsntYoLl
WGNt2ct4n65uFR3BuutwLoAlEY/CNnzpmpi1SDlzWVX+4D+Bf0EHAmUlqs2d0eXR
ue/jabaTifm4mFi7eH6yKrH3RL1qhzb5Oq42Thuka2VsQtbDLOY1Zrq3Nj/DhDCo
fq5JOWHAveH4moi8WfpcCpHNm1pUYvfwu+xpnOh7RdJNiDEYWIsWIGQdJ7bFyGr2
rWsZ0PIB0co7/pEjX6eB3KbfL6IF3rXleZikuCJ2CFe32x099TcO+I9DLf53X+ip
mY0WkW1orRqi5XNlDhhtjK7TEqYm4lh+day3mAAfnkw+4InxcFw8ucOFKMQ5PtkI
zBpXpEBu1EO6282Xan1IfC14L+WDDBy8MxQSmIOatdRVM2gr95t5Qt20osmk2vT1
jqpJpNJZIMfHWBsOCSh+RcFgjgfCTl4DESfwqu24j+wlYPgEv5axdtLvLzi9z9Ou
fOrmDPOlbZEECkDisiSkSnCZTVfVhCxS3FgQLsYUmQMYx1eTJICUYHveUxwhDtKD
27H9HuaGzOoVJHHMxTOyQXMZ5JtPcYIucYRiRXDgZDOraCJsGNNzGqZ74c63YVvT
dyYvvvRdsAObvDjgRknktGDyDFZouORDnBUPQjKVIAqiA1AzmjbkH8Pq4wAfoNNG
ok6j1X45Np1dIfq/PFrUi8ehvXSAPBe8AJJWHbEp3A8sy0EgtIz6h+wmG/EHmpD5
UmsPNurxsOi31ARyiVHau5g0HAcM0PbLxIbO1PYlQVHSsf6VRriI3qHVJK+R5+jf
W8+0I9Awl7jo8p5MgWjeDWPdtVRAjJePicUmeEeTTuN2YAwQk+aAAYoCbF7LieT1
tZ2rek2hWYQ2bpmR0eMhGkiVF28ENybQXIB9c4mX1Ue5PU1VnYTxIjpHRIf8q1mr
qg9AgzymrOm4F/abqqyjNehAp+bMdA6Q+SujtU5R20fnAeE04UAGs2Rj2yqY9Lrr
7VkZiA82/ON5OTfK1rDh9+r9cWeIvjIilh6U2NT6Z6LyN+RUv5p5A85x58QCUzdK
MPBcmvgcvc+YETqzRByVb0gGRSbke28GDPtMAYiZmniNS3vP3HrIu4b6MM1SE3gq
r9CT93lM54eoVa3dnfPWODxkqXwRax/aFUWke1hvScRY/jzMKuYTCTrXO9PxTv1l
YqqOTyUOPiTy/rFFXimgTN81OXExhjyGtEdTY3ooRAOIdbGofDfzSldgIZCFeZ/1
F5Ecy9JtYksWkohSgp9xHvcgLAdVAhRVR3XXM2IXngGAWyo2/9HqaZy9WwjqMUq+
wSGJeBZKVcKaP5j+v2KtGB2SSxsgldi7yi4aQJUJbhYefCLwoKgwgZkcaqr7Qj9G
00FpaOzUayF2XPeMlaZbMcpFTyJrahxgAupKos20Cx3EA7wpYqgJJR1RnuJvl7XZ
XcRLROu11TNVQrZjqkM4fhCmjSEVsoAdJqLFxFiqyv1LX8NeSeSdBVv3M8xSmyVs
GY2kLUFwY5y+PjjpQI+5g7IdVStMyd2BJdYF5l9k9jPfldt+GhnkjerqmtbxCIHC
WXr/MvD0hDgry42i4jPfdLxMFXgs/8Ykk9ojzdV1UEAlL0WIgU1Q/fWIzZ9Ev2jR
/uiW6xtZZtrVwCcpOk8xeEwk0v3wKnzTw43+Px3uzvVwYKDG1rur9d9RrIW5qSVK
sRlzkbfSBU3qOhxoY2vMYZYNWwQDbLpADiwaFpH2ZcnLWo7O6sbgaA9UC4ySdHg2
jC0l4oJIdu1POnsKggIa5Ms6y9/OiYnYPP8cxV2VtM/+uNoIYJ4kB4ZEfgpLKw6y
K1qvNo/UGkX8xeoUtTrvVQrJeZ8laUy0OrjC9abkjmWlosF0Th73jSDJVr/JX/23
b4Eh+ieolLkrnoyjN8NkHFacCTaJqSb5t7sIU+eQDnuNMVxcMlpxgqr6eGEsb+Bf
OKkanrynvAQqE+ticDXhOxrbyav8sZPflKSFmtNO9ESoTSHNaf3iTzRhUlXaZpJC
nQf6IgRywX1lOyfWZJMPfs8f5GmQHGBXliGEqfoqErnLHF3lQTOVTryZhovLXH07
lNdb05/be3I03ifQ7tORY1LqhgBsIG+hx3lxLe+/HlfdkJn+F6KXtPwcI7g6dbb3
HYhmWF5MCArYVh7MG2NsLLHIJGtt6fxbYrGdGP5kcnnxANbn45U1KMMb/yhVwSqA
PmCCkmvJe2Rl9YewzR13jjbyffcL7fyQsFiy8I58GkfOnm7bvKVc1lfPQ5wfG6SO
3mPc8+YibiESqpFqr4Hai75ACFpcKbfSb9dafcOgvLQllACzId+A6KdnS88w6j2Z
aa6omakyoVhfsOAcbZc9SMUIREt83llErhuXHFsw/GnkU3yh8Hl7npZSqLmEEfXY
AVa+Dt9QlkFbCifVwkHRsEALAyJTrwLFAA2IQ7NuyA8NJhkRZPsvQzhVk+gV/IhH
kKZ9LwlUVNopXpbT55tWioVBs/TWZp+y59pU0mTX34MKAvyIze1AiRDv5UpGcne4
GElkx4Wz8K1qWgniEput2WOfmP0mpoa+tqfiOXvAGH2indVVKQ/MOaf7BAYa5F1i
g2D3kJgFqF0ZenOCMy+HzA8zDx2+muMBHin42aZom9Zk7moYhkMg5smy0JYWF/g4
/hiDzuEf7GJ+kY1BsmlnHVWE2Pz++Kk8QFCMPQsHzL+IBSMoNAfByh3E+n6+t3PV
q0Ge2lE6ECb0lf6KQIbR1G5qLzHMt01069Lxx7lCmHWarGjVG4LQc84BS/IztsRn
Cy+9ttR+kRT2gp67KdPzLGPVjadMZTexSMzkJaEo6AMl03NUsrQs/2Xgf7wjFu/X
3wWj3B3qqYgkJdZurNu9A/JBf889v1MiJbzoYBMhQmtDnQnSMd+E0ldXlUzGyOdU
bKfavYTrLTe5LAvyHBvbJT+m0DajBv4SdIRWUWLWYP7L6++a7UZ2pkjKrmcU+u/r
DvGQLX9yAcDBgoRXv6vnm3V8h0ew7gPNT1gsazxIH8zz9arAQFhyP4d4eSWsv7GD
yMPvwG6a8XCxjuNUZMSBLk3i3VJBSCRANRspR6tPCvpIIiSAPl8pNRi2bm4QXAzP
Bb2lR3BY3dceyWTt/5Ik3komhrpRH6nB0fXHXft8q6UTw46EXpJEM1A+A+T9yiX9
Oik+qgEJc79jG3D7pDHAMm0YHnhrUUUtgiS8K4QgCg2j+4wz/KtCNk5AsBbXWs/7
kkDGUWtJUeLjAlG9yO9yXupz2sq7t6/3huFqwc52YzuHfuEAcS6kXZfTySOBGgJg
JUxrYsqHike6DYpN2aMoBC5c3MdFxjji5m3XhKJAG7q4ybxoNvcNp9A9wN+LJeDH
rTWhb+CzAIblnqqUsaCL97R6ma0ukacbK7u3vUBtEeEYzJcpf8usnBvIOF+/Esit
uL+0oKUCPVXKvPo4D4ufwPgf++uC72RhR1f8lk8Yfv4lYoeQB4rVNpmsrPHNmObO
lIZUl07owPB9ybmQXH/A+QCeW+ZgtE/k2nRU3oYIu0hVZqOtTtTFsi5DmXOmirU5
ip8c3MjPsle+ROXkIs/GDQWsXiMx58zAzfiaJNyeKburXQjY+I3VGXDSYEppJPJV
p4tzZa8aT/ZwreaWc5ls8tLOLh0DauSYb7VI0qPlhXfDT18+liw7V4xyz4akAyjM
Yt2e/AEON7Eyjb2GnwqkHHvw7XGt0Kuc91GzWKNLo5VzZFFY0G3ZSKN/ji8eAIt1
tA06Jf2f86ZDRmVXVFLQVfwivYLtAuNlmYcdP/gDvwNFUyY5IX43NTRMIU3diC6J
b+8XWv4v3LsuCXx1h6Eb0KWsAj5YVx8JhDE/DTheNBPWyFryNHxZgWwqktbvkRel
6vevBPxh2apSOlguKkma4h6fQPYWZPKQ7NZ77IflbHHEg7hnzY1aDjJ9TH0xP4Yf
PYDbOJpVj+WpX2HUmYimxLSMv2AXAsEFGvR5VLOACe96TzdEl46ybK7qEz+FVhWz
5qZ1UCrq8tTxjc23xPOLn7K04vQuHhIEQOyW7Ur55JtmmwZHl0NbWYFoyVLuvVzv
ggt4oaQv4x4z77hUDqHMhbZttl/Tjxjbqg7f+T1toqqUsZcrPawrbMWTvycAnIMC
aMjcJGskYCtH7mgzlzoIMR+4My8IhJ9QqZN5olGA1ffTikzCd6W+Sp/1R4+VE/mb
yyUHCX16CrCSJ3gEVqfnb9azfH98QXYbXB0bFqi4HCOvjvZPCVrpUGQ2OI1otgcT
Wht8iqngiz7Uc3sNZSxSdjhhD/uMqWRg+3jfny1U6EB/pwTvjcvDH1zlVVuMI6cR
ZDmR3IEeJZ9oxUk+pbI1xJHeDWakg/uBlC0NAPKxJWBld24Zl25/WxjQczF/cIGR
Ku6thivG8ogEi/NMTcH7vQi2bYIsG+rv0u2ilmYeWU9IEgxON+8rDfGXX3J0V9qA
PmmBwmEqTK52u3pfhCf6ceiR1Pfc5ajUfgHIPMm+mMzIPJHtPIobl89SNyRI6yCl
fT3IKpo5pcNDmVPJmYARiJar46YG2ylPrQcC0/apdVgob0MF0BoTPUx6UAnHczBI
TRJ1uFPwUBqhCcODXkeI5Sq+6Goh3GsNrAZ5uJ5C621rU2NtGX2lPYmpd2BO+znx
2UQFB/JWXmxk4APp5q0tPggsRRe+2XP0id8nh82xkADO21w10VgQiH49v/RSp6uJ
4Mnc9bccwcGCGgYE1eEZL3cdLev/+9uff33f1+U0lqL6Z47sp72ZiskMntbzKLCl
CaLCmtYyv2XztmLkvmmLiiJ755HEAaor1wDqTR4kgJWbOIrHCf9KbO21RZyMHFRl
d6TRZpyJxsoEXCpqyCJtMkbRUgKaupO7JDn9Jm1taaXXWm1jklLVGPgl9dbCGAN6
gUUc5FzahZaAxaWvowuIsFdiwyz0az3+1dncfwXQP/4lGanW4AzhFv8KZ6IC4j9Y
KLc7oxk67qBckrlJZ/mkmcRW+N3tyD0cu5oslQJ3iEV1AneXSi32fvV2osJfBzJI
x7/AsSKcLJg2sbQ5KIwOrv/+P9aTrXS8P6SjBwgJ3mMEnOPb+3mpNa4N12a/Viep
1+mUzqz5XtVMsfxkdjkE4kIpMKp+TopvKNuNAFtMeiEDc2mPKgLOqMNfPPhNR0+/
4dSYqdlxM6Vqc64NJkm682IcxpiT7jBiDAffaUQZvM9jQPMt7w6BcRhLJ8wcaBoL
oL4zcFejqXd5IQOv+llA+aPw5K5BuqJPGuMCOK4lnKkVTnPHQ2ojrXHv4fetm45Y
fCllyGY55XESI9mdyRJe2kejbDg/3zYONDNluHc5hLEc0N4k3kGixka4pkihokF2
WhUBgXUAqQw0YBzAVCPwdaK9u3PWJlpcGTxp7cRw2oG/KV5N1j2KtXleu8imrW/x
XpweO/oAyNGH0i/58BhGd34rTGH/hhgxKL4HsoRy3haUDBfACnDtt6vFzKFzfnbd
C9xvoZyJDEmvYSbQKZ3/Gtp3TceR06tckHSPyhm77NUbfirbzcf+VoIHaKELqqIF
lmbVc/GajnrVucMM2jp9gC+l5JiBlOcvbP83IZcE6XSfz+gae4FCIM9QVJX05VIq
V71hSoh2Fm2L3F23rVRS/6emnN83FujmrzJNyuYKGXEFEWyY7ZS5wQx7HgVVonXX
8CSaWMnWhwakeD9inRCe4NP1EimfNcYLFkFHPTOgfyFPLiGMN7clktzgJuN0u1bq
eEjhyL5rh5qSs1DuC5Vw+FaPQYDd3pk5IjAKxnRkZmz8h6zHCLf+SFJwpcf56riK
7CdtFpYNg4pINbusc2bWS7B09Mi0hCQi2cgJj/9UBtBTWdicuVW2zz9RM1kJVgjr
oA57kM/emDDzsiwxVDLq07gX4Df8Fb07kOTygVVzT+yuB9j5NxzjWJgjRZGDLXKH
WHcb7pzYAxNvuwOkrEz/gTODyq2XO0JKVXmlbCXEbf6pmImCsG+2s83G8KZC2Xzs
itdkPNcdp6WVyNw2xsv2H4TOLc4HxevHal4bjWCeqt7hCzIzeUu1Ui/6BKwf5p7z
VxtYkONHueuTkq9TXvJXrs+XsyPfJ1a88txZwDVTQZCBpuTRHllLpiJII3Vfhiiw
qUw6nsSZUyjoGWA1677S4KVlw504Yq1gjoP4U3IolduQBVJ0/BNJZ2rHm4odgLFD
8FgmjZNsLPIAHIcl1dwwwj9onOtBEHrQEpAhW5njBe71860tl/3bS1m6f5J2I2ND
IWFpy2Ft4VwUVhAjWKT6myld5q/n0dJyBKEbR1CHjzAeLlnQJkWQHhjyiRVxk7Ja
K2hr7UJ5I1/5sXMs2leLX6KHM8KizjUIYkE2hcOuFCHBaG9ByIPxQDoEPKzddTeA
e3ArCfWJkDCN3OXGECJPE5tweX2NbT9oMvX9f57985n8F1EFvKDVIbeenXuQJjp2
1TCgHmpz3C9bUnHVdmBJU2fWjgs18vUfWao92/cyZXKK0euoohd1vWo8241jNY12
DGCxxS1oIKeg22YRC0LTN4dIrDZJkNdKw9Ly1Z/DfMH+CwZqoZQD2LvuThv41jPV
clDc2VroGA616gkBA/cSprX4vcK0TNnKr1PzxbD+crN2YQVH8n+DCauWF/XKNUkz
IoFRrYHaMr+8pQV4CaBHmJd8YB/GQKtMGrzWoCIYppgM7EENFqxg3bi7oXM7ZR+z
aImCFwRQhyABj8am5kpcMJa5fyf3HvboWTnmQDfQ0+yItuuw3kVKRmfSeI9j8I+3
0y43Ti6Dz96vv9v5UVEa6CDx5CwQSW4iT8QP8EAzE13NQQPLP09G1vtZg8unWRts
M2pPIQ4p4YNmJWnNpUgb7Yg+CAfWMkYTfSzsE/bEiFaKaN48AggenmJvmuogdBSy
EfS027X9OR0DGNu4wiaGPeSvkjDaKdu2SARDwnaQNOatWwOfsTSVABc2WYmbYQuF
bs2WNCCbFhyClRlNVSVfh41dfCN1qT4YN6ndSk0MWnRoeWUknLdzVikZTIxDRH81
ozinwNttZt7c7bhXmtfaz34JK5DvaQ+CGNRuF6x1t+32IJ3VaAo29EgnG/93V1bi
RN7eAAje3t852RLue5hlb7GNSe7bfQTK0joNS0mh0t7jtvnQ62E/QS3IHovdQxpk
ipLfk2B2zh2cSp/JhR0ddfitB9wkGnh6GmMK4XuItb00qjN2A49yZofR/Nnni5cw
OikY85wW7EhcK/5yJzMG5wb3+OvJhlbRR8fuFmnIiE0xEr1sZP9iW9zg7sdLEM2S
xECaweaxf67xBcIKA7Q+/53ok6lHvfmWt9xVaZ81jcTb5eslIwIXWcDRdIeNjDKy
3kW+7BtTc8n3p7LNcyiqxDd/s7T9ybZFK9McP9P19X16x4HDzvE1vPsYdggyEvzh
r0xeLzbrhcN3KQXZwMoZf4iYoUukAx0EUUt7D/VYA54rGhgpbdeT98CgAs4nAp4Z
55vQ3ugGQf+3QGpGlzRfzKz9HjoWhIWe892WJNY5K6y/i/41VUIUUDbOXztW4iWq
2oIDUr2LY2700pj/wkdqNwCULw4Mjt3gyjbkfwtyqcvz3nbe0npsjoUk8Y2aBMTf
Qi6eiTPv7B5uKJvu/TEU3TUckPlDYcVd7RMb86GD47Q3HogqWdpey1zq8WA1cuSX
jpWXBssL8AulnaJZIOffv+kuY87xFLfCKgApTJCzwFu8WGCzsj26gNQukRmMLYeq
ut4n9UQFm4n4btcWEWafCBIRItISBT84YgVoQpUPlKlfoJB8BVF5hBhnjNLbO4Vt
ZkKoyX36ORjhc9VI+tz77HfWZ1vS4AwJEiDSt3xlLzTKYc0AMIg995KOZKKOWbgV
11aEP0E65176xbL1pT5XEXPjDiCZiC8QhRgI2xO5z7Eq/Mus/j6YxY4NQTbINaxV
3mZSxRuL+HHUzq3b3VGNE+qRhR1/+xvOcBIH+/BtXfDZWNVevixpKAxm5Yod3DJn
582C1ml7qjq1CWW5eKq+VyGf1jxuaEQFaYrZsvcr3ynKNaWsSXDVwN2d6IymM7SK
ph4jaM+jM06KsJdaCJfjUmWH62iCyaY3AnkOBXyBtpE3vegWOf0zJziSqcrdtU6m
2QV0XFWKzlz+hTTqIJAkwYSWk57ce+ZMHXufmCMiDUrRwb8S5+Sms3OhfATSo6BQ
x0bb87scTQcgoE2wHbETrwra55SYSS1d273rV2gAb/7Q+ORpWdEezIPLtWnvQq85
u5LTblFh9DThMj5OJew5h7AC1mq9bMKbpSvbll8couaaBjF2GwM/9oo8hG8nk3Sz
qdHglYIqJXqBT+/2vU3qhRSrOfS5ZRFLARgG2p0NyD8IMm+ZC9ik5xcZVkeQv1/9
6WJbstjV8zvrTLh57vj3E/08SB7Sd+yHG6g+Bt38Td/K092g0z4zP3vLR2bEHoft
8XTbwdFJVEjhbMvZibaxbqzB1Vh+btufXHPGUt4ROtb1ULvmYizXpltqM8zF+kFs
VL3TnKPEST8ehbjOiF3QOJdsIhGBdnlD7+fkzPAwMpD3ke7ze0VcmhxttmVhcO0+
Cdhef39p5+g0poU5L2YXoDnvCjnFWFCm0XO43z5GOjSISMQ/KnLWJJsnVEhCfLCK
4iGHI52xXnx4gk6oGxwUBh4YFH54zE8RkCor1JTMkcd9az0bAI8p9qyUHUe9IBSW
126xl3klQ95b6mjDkBsgGiPxcIW/PcNnm5UFX9QUdRls0oPLIiXyHtNnpPW6OBOm
v7MN1t7Mxol0YpBqUF2KqHWOc4QdhMULQH/xqgIZRI71hd2f4yuPmLJBPscVBLsq
M3JI8OmIxjHIHa+GVOkpGEtKMjIWZIMDeQWWni2i8aE1mB0KeN8/JqWxsG2ssyCd
sKy6NpberWe180eFaBDmC0+6zs4t6PiEZFEkIKWkVDpuh8GCd8dp5//TpU7BicdE
4rTmbMUuWZtWX4algfrpONzFWUnVId3F8kGskkQuqfixuHqkZ2cwDSpefqvwQKqk
5lkbrVcYdjqrL4EfgrFNcpPqj+nbYPHLPEkkpG1KFxHOT//FqjlJrE5faqImluqF
jO5CZZ19Q0jZjVdZjhZplPVGOVqOpW7PeD5nLODrOAWPL4kgIUZeX0UtoC7Cektn
lETWsyZmiBcBcH1hlHgpkmYjCh4NE2PqW90Q6KuloLkxthm9coxQAOnJqXQ+Ylyp
qP8ZrXrm8IjuzNHNLdE65AkOC/grnAPjY4xJaQhyUx95ZalHrQiH8jQwBc+LEaQo
GvEcdzn1FgDeeni68giYn2DJk7xk1AytD52cbnOYS4Tt6KAK1hpfVZm0IDao/9Xo
hQKGV0ebYIoZ5hykR0nOhHkBA5UAzezf0KLGlLGoE9DtThCRh/GXtxI5/w4Maptb
OjJLTeSmnOeQsfyezP+MgQEKhFLaQmNPA3K7S0ya+xiFn2klfHC/zwd4cdMyzae6
4jlsa+F7CYVxDgg8Tr2yd7pmiUbmVP9n8Gt07O7hbrvzHVpCOya7d7trMH0kSJcT
YpUWIaTi5HMZODidOnOZ/QKMp3u58+rNQlcQCkqpaCfN2/p5Xq1KlezZ7DBxwdPe
lqXasRdvwlZtMnrJkXIJ//OSIOUWIhtx2gKuYFdmgb33lCPuEWzR7pxL6OejugC7
Erp2thzFWPgei9lk3saLsZ/2tkO/bfydN+GEF/YFVi+y2jZGlxXgT8jrCenWdPH+
J/8wyS9wBRie2bTGBtr8nxfr32tl232Zb3H3b8C4bYbwvYySM03jmFH8mO/Uem2A
yqLcLnUz49gwU/nWVx1omVA1xBNHYrUbHxlKNU9UevlMO1og5T8ulBOOPoh1C8Zq
h6IHzKC7FQnUGcrJfqmkEb6pruju8yfM4YQKUxcUbB0wsv7NPmiHbPr85GRasQFu
lgNNrwwOHSTY4qs1qlRqPLg5QX6YS0QsbvpzqinQHtIhsn5qbsJ298UYVBzy7Zwk
NU3rl0cVIdrZ17y701DPGv+VyWqzhb++xyA4izg9OPe9naOE/T5+tWuQiEyyCaWJ
c94HMWdAAosanIqH/zMHI9ee8H7qEj74WNSolKWE3XTT6oaycqU6z6Cpw3E6LjLP
s9WMhE4XtLwSgX3yoQ9MlUla0Tu8pSFAH/X4wH5wyzoFvAr+2hUkA4p7ODUO8jsw
D2hxNh7t49tQUp/Imad0/UeLjRDM3dW7NE1Gn9xOe5bpjtXva0TfTDOCrGev3yAo
5i3EAOJT/yGAzIJ3pr5QjkERJ86zUn4btru+Q10qDR6p1G8tn1uRBdfTDK5NFiOC
B8ne9PSc4UALZae2S4lk6eD5312xsAA8eSIdbQ4gFwmXx+jNs6em/eIWHSd1FGRO
eZg0DlaeUrhf7s733tU8v46j/nrk6rOlsr+XQwtbcHRMfhVjwWdi974v9X6OHx49
AFM/+9lVL1upvOjD+QSBM/I+Mxe2yJVr8bI4QXQU+mDZcCJJU8NqM0SYcRFxytUd
O/Bx3sDO2uUTjJJ6qoauFIqhGSCgz5tTt210B5XP19o5q3xGczzHNmEXF2DHFnMc
IsV/vDtTPgaCiiQshkzWsRcmNU7ZLWx8GGY1hYswUOwDmNIk8H0fvNMNhy4KBC2t
Agmm/jjMcsVD6mbSLrgPRf2SqnnlS7qEffVIthLsJE+kfPfeWtYGriioCrShbFap
xZjyHx0bNkUj6xlJdJKSq0EPGpfdOMphfWIiYMwlBo/3zZ4IcjrumVeo+DXsU933
P8Hyu84nrvaDMCHukAiEwI6CtRrlkJeEgQvtn1TRhTOm3Dls/V5pWTMNk8KOUtGq
07WGk3VBIuQDQMXEj1ZLy6L7/9b3HjMYAIGvy0BrIzYY71b1tX2WpDYvGtQKSAjh
/UTwopAdqtlMsBxkU38aOb0LdEv5AIxcJy7bDwFsot2Q3sFEFgENWmNhhlNrnfZQ
bPzRmNgPEB+rMOaJYW/7oONPbRy5eXCeuyIlu9B7OF6itfXPylXJZJXc7LvFvqgr
vSxPUPXhJ/08aJ8mlnshPzR7QPwBJZCxH7Owa6I5/ifVj5nwnr9Kn8MuXLAGDZmP
q4O6Uk5XnBwGPblc/M5Htt4Y8geccj9kECnCCmnhVowAtHVijVTG8r+Cls5OHn7w
dB7qVZDB53qkwFzqtMUa0zdlQD+2J7+CUuZwa+z3C2WC7d9hN6EQLz4QMQakezeL
mD8+2BWT8zXA/gbOgLYLNuBG7irB18/EIjB+MrkkNrMxenixQTtIOheja6y8BvW9
cd13CDHmX/WYKW0kMCQGOtKrqYwtZwwJYOeMTfy3o2jU6OzZCi+07agDW3CHAMfI
e9Mni/vyk9tA4WKNcVvC8hc0aFX27Ak4ql/aNayvO3/6fP6k7sG/wkRTXyK2UZGj
TTPGUux9D7nS9y6YaeiOBG8HcB6rtT2YkCaUsSUdZZs7jYdfzwN34bR3UWrgACc9
rzbUBu4DF7aL8t9SAXMK+xeLitT0OoEnPqcMJf9P7wi1er4D8KJL54l3MaH0rp+i
nsaDg/3XfkVmWU8LAxMRCKPzP41wtb4wwy0V9RUPYL5IDwO5FiCbBOAJT6Mu6ELV
SPjfXAxydEHtpfrETMLc5clvtxHbI4L0UaQOHTU/kcB8CFsD05ILJKoaWR5NKN4y
ZQvET30A6hv++pagfPLxecGDX+CV1R8BmrDyW7ldTyVjK2OyKT7UrXId9ueNGgvh
iE5/pIdPwsu9BBC0uIL1NPgnbu7IeHdZOmprBKUhR1Ebn6gGNmW8OceE4qcYD4ND
2iI6HwpELYoE4InNxTndnD49ZClUQqJY3sEZ8SqduzZeMLM7B6OLit9naye35vI2
C4nLv752Mf9aG4Q9bU4HEMSRfjINqNgbfhPS94z1g1tAx5T5t0gkOytWcnc1v0ZL
i7Gce0AWlIcaPtLAlErOai/kkFccNRqlGjaqrKcQO0EOzb4E6eyg/b8VTBEAIEdh
N/b0CyJ4JgmviDuS7XqeWzqrwNho9jaffFr3eEI4rRi/peTnKwCEwz8mHfjmgZ0x
wJfcjOY/j0pj98dkffxyeeM6iobj0qUwuowNg5qu6Yq2BYND0HFO/hlJjq0gQafY
1Cx9IqEy+N5ZX11RlGq4MjjSN18eaUMnVqDWdveTnuZV8tP4ZumNo8tueL5fGW4j
bKeXWOH0Lj0Q0FWG5cAfaUbFe2/axbMaVcX/vTVvuSxZH//WPj1V3Rz1iPsXvFhU
H2w6cpr8WfFVhjJZ4B4ZzGPjHpAlWWlDwThaxll3/jYSsl5iySb/E/xrl9KDwESr
ym3qFaeTxZfwTRfE3KpwdY64rr6oMPCkWVKqWtc5nwbKjY9jDe1GFpM0sPFP+KHc
QoFqK5JBa884SINavC+6V2eABaRGo/Zr5w47whlE9KFefFlUYsDD5qrVeDkA44b4
u+lejeK4LjFezQsXrLHcdcK6ihtpufQgOk7mF+bPG7w+daevymYJu+iCi/Cqv+uT
5vWGIiuOEP/nQ8iZL4WcBxoW7R+IMSqq+8fPlp9zO2aMa9J+oRwVbicIL0/9Sl2T
ZepMhVgqzmt3lg4pT//5sCuYTYAoWIVkwC+/+qbViLhRhnuwmvBkA4X7STCmyiRx
tvmh9PK7wFA+XRwESxBtHLUPiACn6+tZAYvgwvyDnYLsXMfJHGyqePxPrvTy43jw
jHkrCyVzfogYjn+g4K9y06lYHAf0A5SSsu472Hz/3wsFc3ztNc8vSXG6MwnpUeCr
rCNfrwyHIiP9csP0EECw8CUdIebteI1jdKO8ssWYBL55J/4pCmxV1p6MnYLMOfVT
dQbT83Trsh3YgdfajVJIoB72y0yeSB7LjBh1TKkvCDnGcKNwK2ZY0auoXIp4AQoz
u8+tMqUa/QzyrxksQd5yYrBBWaBsp+KIIHhw/DCFuDgwa02EpFF35m/hJ2sABc6p
gUCIDAnzcPjZ9DaZKn7VT0pd8/fR18vHB5bl6nM2SNrXDxSZOqHpjYm8xwvoRIjs
qxJZFnHIRi4c7pdx+B84/jUwoQE39263/S712+EVzEpqerRxBWvEchCAcWcsPbf/
9ZszqvHEy3I6CwhsNcEFm9XH0tBw0l7mWn4ZnN6OvxP9D1iE8iuGH5y0+I9nsb9G
hH49P8+Chj3B7taU5SlDukTTcZnAJIr7xvgudX7n/T2G8NiOKOgJCArY39pjF5B/
hy9114ySv52Ck6O8jReXEFIoGg9DHdMsRxQI661a0pG+UYiDVHRJQ0B/fjqxuGmq
f+vD7qo0ZbOsTKbPaCSY2qPmOo2FFtfZJwc5hxWsHunQn5Sisy7sTms5L6ZF7GTp
m8BamDv/U+dp4mfAoz0NflFjQ2dD++jJwzM90jXCJIwv1Beg/vJHkbWcW8Y3BrX1
5fsMUlbuGlKyYta8xIF8FZXcbhToVskmVZglNRT/Ezrq4xZ0NJzykRdUFlvjCgwP
rvPzl1fKAdqzVEKVUczUJSgBqln3dBRTMQNa5GBFC7KTfdk7L1KXEq22tzue+/HG
cML/L+hdsbUcFnq8//Vpw6f//qMjNm+gKiW7KVrYd9a8uaOqTvRnRZcEWHfO16cl
XuQxemggRI8xTU7/zPZ/C9VCIdwNfQxivLx7iZAqeO51QmkyCokyIGbYNc0LbzvM
h6yA+ezyB5CCuqVkjW7R/qCVBp1+udPdgcfOMfMrR0ZQnbdMPMnNeGUnL9LV/RPZ
amE0nPvgt8Jvr0XZSOw27gD7UqaCYtKt5r3KcxLpvE7dMR3gPE3CgaXi5qNz4v4f
qoZ8ELK0V8OX0bZJj3Ve9cOLa4vQpGmyjGjahKEHC3/+qJQMSSZhkDEHdvSoli7U
Pzb4ER0Q6O9KrB4nBUlFstWCKOupdfxlFkjnagXzrDk7xJ8cfbrRPAHb8JWawSQS
mzvT3sXF9LlcYzMD3+tcX2NUGoiuDkYvKumfzzzS598YBboOjILY/8sXhJ2W1UwW
ELH5RlXYptyXey/OzJrwEKS4wJEziZbSQWkG22rVrTX/U/ZP5mwjDizge4EDrrM7
g4pEjeCVljy0pH1vmYm8iMelf0LK3+XdgHHs8fzY76/BWQYp4Rrse1qMUKFq69Sp
8RfRxf8n/sNzYcSlgBdmkA8AtEAzrU3kMI+mrNTPBv4DIfIWO25ikBfqTs7mmOg1
nWrlXGBXM93T2jY8yB2Q1bojoSFaslr1Ffkx15crF4DqCVKoq7JMiOREU/nIfzBQ
BXLxP0qckloIRYVhU1UPuA==
`pragma protect end_protected
