// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:45:27 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fMosCnMbMZPZBWADNQsM1BAvHqD9TWO0xwLfu0vTbICu+HcLQGQVFfuA5dOhYpRn
R8EcvsnJa2dxSZDCWeORPm7IbokzSF+VpRiut5BFs+ykzxc22MjedKKuqSYJsKOM
vWFX0Ko+rVW7Ma7nZizb3Ai0xXDC6Sv//di8yUBhqmg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5568)
gOVwqEqxml2WVbkZZ51qsaaG9PJPgNIzKrDpS0F7rnQKDlU1uxLzSvIGUluDYNL7
LsgGbgL/UdFIR27Cxt37rNEmDtUeRr0rJTvlcQ8MabixvyM9bYP6SnC1HASmGKFx
k/mDxA942KeVyOaeX0VRj/HJnUBkO1P2CQhEc+v9DmNI69+hMiTIUooPa0pNIUI6
olgeVLdqppWhV4gh61fFzJEbH8IIpsaLy3JPfgZkE19VqZNZ4M6o3/TLHLkPuhgq
Rdpk/0JOnhDDCOLf1Xc0yaqTDPgFR5N3yCMuJYhfANrNfqECvr8LZyiinp8rRs3z
EGGpoXNuRnM3p9BqNGYUAOOfYTqaaaNQaDd1J7pclqSQwXBdnZqnToYPic47OcGG
y6rg/jZ2Ua8Fb4mduLGU8x003xA44PgQ573H9E5/X78447scEpdcQm86OqmDKYEh
a6Sh2bF213e82RStPy2Ga2Cj9mDFspWVhTwjjy5QIx6atV7kawB7+eGIjCMBWYIR
r0AOVStj4hlESQqEYskcz9B0OA4NDEnl49pINOzKS2jF1mgfZ6zgnx3MSfZYJTPw
nKSHZTUkZKCTxaLoN2iGAQ69bmyQDxHIOXgCyujz68x0TGJ5ZFOzwdeArkUnBv3l
QSDkmrPkASxB+4IDwhXFdpuCiOplFrQ/itOvckNCsRKiyhs1KQm+5E7EzkflH+ju
tA93Rck9bhwuiJFBdVdQ8XL6efUvsvJvSbaQmOKCIf3WF/T3AHsALq+wwouJ+uvE
veoZKjsMN/CUPqsXYLfjpMNvfC4VFiGIZB7/dus6IgIHrmsRUqri6t5pfSQy/fEs
2figemEAQmDRtSB60/Rf20kaE0RC0Xny6ts59X6qnNSAfnR78Mp9cjvdLhEj5xzv
qev+cI/Y3nxxBdZvBqqu5ID+EGNpY6o02/pswNhd0sMmboF6XdaX7KivmjYf3cwF
HKkD/AsmyDPDKhDEL6cTUIuKqLx4IOmPIhYThjhoGxBQKTQ3sBpmIvbXeTu+ZdB8
jEAs0IB/AnSexnMwO3OKfK464FHhm015ic8xAdODHDPyOjG7NX6FqPhVp33yuDCO
oerojWuiYDKeOny+Or15xL7xNtFXUOjsORA//uDW73uWFwpc98KCEmGxWR3zdLaM
Y0ASXmXQIt8fcZU/WD/e8T/D9zRd1Vp1BW9HJIAxkYungF0PLQuBw+0MeKNo0LEi
sihWQfd2L+AWlX/iULtPEHEGEsFHnoCt6SS02GTmEk7tXc8brLONvnGpPgh8URXo
hfuULc1DDQfDVOKic7YnLgdZ3x87tSYQaMo3/HZZ//7JvU+c3P/cnUG0kL+X1OQ8
XdgyDpjITHQctSGrzHNAAo9KPA/XY6+iUUJ2e8F6gAZZOCLyafFt8xe48xJiqBH/
lZ5J1EVmu4oa95RFOxCXGX72km3rVgvB6xzN1F7tHcguclW5+7qg3yyVMx1KmwUN
LCJmAoH8RTM3o3Yk/5zZx9kPpD3I2RUiclYakPZ7GQ+W4P6ClCH8NctzYhvpZBgl
fGeZ+iC1OxlzTIaQSHRxJ37ND3MKelKIJ5yesx/TdaoGsNX9cFh3cFJp3ukjtdsk
weVy/We2Q9tyt2wz4wqX8Ly4tMJZWmA5tRGCQ1JFIi11S60BqVWXRoexbPyZNXkt
qZfY3dOn1+76QQAfuE59FK9wiKT25lxIt8jiCsnzlpJ2ug+zLv/8/Sf9KkVfFjQQ
HIj58Y+dJb+TR6Fp7SEQbyq5tTtP8H56bCaxAv1469vYsvRfWtfpHh4quSIsmNxl
ttQe4GgIwfe0FSKA847O568EADn3wLpSkRox/RxjXHZiTn14nL9uQmFT0jutmhUI
KPefgwxWnpRcpNqatpXN5BhPcbhYQC6R+GnDB301g+0nyWe/WDgdXcbvGK6gfUa5
ADUQl9i/KuWfeChSxPtfIeH1VUV5sIX0AmpS+qrCMRMbzQL9keHIYAgOAQzRAcYe
EQfIEvkhIvKhgBYXbrzPhAEtyN0utl/yX8jk/97ouzaA2IiVMSfGmj3blwdxvxlq
4qp55TpizysdD50nhcDTex2Zc70i8yPxRNuaIgPA37MVJuqiqQJr/vW+0frNtEpz
KB50uAiVCa8C3rwqNqWFBTsGiCzcos2lLJLcFqEzDC0srzRwIwwDccZTh1kBX8mb
mb3yVf+/pMGIO07Lr1MbjKU3qpua16edFwP1QmXe2FHm+Ji5VR6XNYgz5JeGifgJ
wfHcZ1kh0HrCgqnT/QjEL3rm2zmsKCr6DXHVqw7PNe6nhnkIEQjMVnhmb3cVuAsw
8E4voRsK+tqclsKogwDWUnQHC/e4Lk7tqkFrG7V10TvXW0CjX6tRLihnKfmpvTz+
0im2vTGaNLIwuCEut188jCwrVjayyfN+DYfathYbxIyhsFBUR7HcC0x3hXTbqah5
r3vxqmD73mo/Bkpy/4FQ0clhUgrfC0MrvM28eZx9JHCixCvz9iHO4LB8LcG5SKna
+uxox0JF9qgTelg3X3hZjgav0ho1DflCYNQoHBLbPYzROxodg4RJjyEgW++NAx9V
uZQUUXzPB1XLJVAcmVNstzlpyEWzZNaGHHAX02xsLFtIpCpO6K0Fuw7ixEMImrDZ
w4GX2pg77sseq3nLpocw0SgyMwLt/tGVk0wTvinQLaNBLWwkQy3fOoicxW8Rbuqn
/+f0hZ+8JCIKkyVJwpPwIbPBlw/TeaeV8OeL8dMxvh1mbhOx2mtViO0Ex2AVAeqW
+QMxEBEvq768BqrGqdhmztEcisbj/QKrOlUN9tFA7jjzT33Y7QgPK8OQV9s8zkq1
EMvCkHoq9akwUPQxxmPuLoTzy1/JZYxshEkcgzp/bcq9MDb8aCkJBYxiAA1Kcu3A
AKqcstua85XqCpRU4w6bRmMd9rG88XPtRlq6I7tKadobFXC9ea/YX9FlbSPyHDsg
RWsqX6GiBcF8HbeP4d8zLyRbRNRkd24uIBXFKhjKFgiWj8Qh8/LYdjkLP2fAlGal
oix4Rpm4lqSSLmcaTbMATJ2vW2kWn8MmqL0her5H6EJXplOR6GW+HIufbtmPaMJb
9RVqKVfzStL+Bx2/4pb2wYSppJ6uu3NBxf5gngHKOpyL2MWVGbX1FrPW+9D+W+Sx
Pa3znRhLdMhvLAmINudqTfUOVoqu4Zkr33mujlloeKXKm03oCENdT8icOzmOoTHF
7LNx1gSMwUfeY+Iiy07oo3zRSTZeWdeEgWFq8YYmj+47WFxg0n++Y8HvtMEwA4sE
qMwslyisoiZZ++TtOxMEsJO22AWtVgGp2idTKW5Sl/dhxzhxEXmuSbUFzw+JFM4E
1n3yulsH9ouHwqY3w1ukCPjoI9wCD9UHhvPUbRWqKzuJy1aeTWwCiQBQy8XlhBqw
O5LGNC5ea1UZgEg3/3r0TleLZjL89zxz9P+1wzaFU2jlhQK7vR30VCDXiYgZ9Yi+
Iwg5Mq0+julm5Q+dS40ga94UcgTJ5iv/l1YcfRgIdh+Dz1Qj206Kwv4sHW5dWG7D
T1AqBYX9ZCwtYRcFkyvaB2C4X/GtmSK4JuDp+XFt0sOUI2GRVT97JGrSBKlILVqI
xVT3qcIUTlDTH5kyBYWydGN1ewzxCJrlcSYrQjHIOVJmE5+wFJKVRo4be6kKRdvI
2n76pT97iZxCmldK1ut75AqY/e2kR9Pk/f+uWWciMIg36vcMqyl30YG9scYAEkC/
2QQ2qrYZcgmRNetlmX3nx/4QayArvfeebA7tyOFKm6HX37fxTxkAwn0qskQ9G09M
bDwKA+V26KYpHRDhRoBe1opfoksysC+aI+qkHMcstsLORGbJ4kMWEXLlAn3VgHgv
s6aUDcQS4WJDowfEZII4gFYocmNWxSQcgIEBmAUe9wCCriBjuAxuhr75bACeRqXb
WYCH/LeibNskElPCTT1CF96/fHywaSp8wpRhlmEdPAJeTELJyRL4/VS2c4GXXNdm
6FKg7DtfqEALikvj4XLMuu2G+MCjP5xEsS7Ekf9aAO9qGFk99SLRCUnLGucNAyyo
d6mRH082GKratOhCF1nixroWY1CMWWuzE7KMssm2OCAD01G9uq5xxgkZoag/aCg7
Y3o8FqbeWF1RtxSxWDXPQixf0k1ufFwP/uAM7NYjHFC008d7CdQ2/Ib8PXWOQo8h
A5Cd7sCMhxjKGPjlxYBZa1vTvHqBZKzwt6C07TReNmsYtsIC88uT5CLQo00w/uhB
qQQmPzm4CjAi0TqRz0XdyneudhZtkn4gFz0dBLpp4H1WY2FdPnFwLba47lK1hsN0
x1w+rDiBWNGEpE+Gz72+KAJSxZG8qEW7HcKhXkMpzhtpWvDJfkMkwCrGT80KPh5r
cQEmMA411EQeeRoFfP4pmGcd1JI6mfBMV85G2BdAVaxFv46obNCoJ8nHnjkMdpaS
sf/7AoqJ27YeezBahE+Rqy5nUcDP2RTzw2NPUeQJg1H1GgTW8dP2L13JoDpA0Uqn
L6x6eM1H/Y0XOqm5fEvEM7VgvV7UUSBGgQZNwUb1Idn9HWbF89DVuDsaEGKp4Ao9
A5ZXkZKMmIb3VQOUbEEJ3t5KdM4ZL5CqeGKwqCWce69646D9ZoiGoa41FpLzGrRM
OJrwq6YUZ/go3bOGqMkxPp3ROKdhb9C5w+vng92xgLjmCagn3H2Bjx4ITcDaopaz
Tbzp6AchjBFicAt0Hat5nEfP6pexhLVku8XIwzbFsgEXg2EJ98vUyL4g8/tw0PUa
iQ5PldvETYtiNDCUbyNuEGdWyYpDJmHFtSPFKLIWKa/uudUquasRisGv5xqh07W+
IPaTk1TCH9kMJOwIuHANCzr1byY8zqwf4dxZod0ocPHqngiAIaVDFaV7e58tQTxC
NsIxQ/oF7kHeg6x2WBR3ZFr+w18Qq9f649nvrve46TKz3vnm3W7R/VRZHPXjJ72N
naQ3q4VbBOSIxdLXl7x1L3lXKtJBJz4gJokkTHacnqVhkQntcfoQ/JNgy9Dg4wdE
RodtwsnnskvBAtRDV5hFQS2O6hJL5UZGUoe/H3M4ooUcBqP8bI7HooIUa+RsfNq1
udAebtPQPrZFpL5fPmxOXA7H5pvwT4jA9dW0HGX922eM2l0JM9izfDED5YQ9HD6z
y6bRwtfbDVLfsQ7bgyjIJUthiGod4Bh2vuT6NNgb+fWGbkwEUdROyS2doxZ2DqUc
O0q3N52nD2Whi7fJ+yvX2gXWw3fxdq7Pyj+NStssD25wvPzokEMXvuc14wPvqcMR
H+HzLZk/w0Oxe6r17h5ORWg5rmmCmFT+oZiCOu67HO9DHxQtWe4vBwtBs/9vA88n
Qp+kiOCt/rXkEXkoD5SIMHj0eio8I+HMq43p+qoxzq0GsFP4gaMXTz2b3E1f4uwq
+p+SKM4GGxntl1hGw5KyrSfbazGIYspiJQ3j/CMKA8mKNK4mkUVtrEcECWczVSIl
MG86d86xGWOB8TwHCIjalZ5X3+3PDOeYAlGhwA8zL0vlu2NxAYUnbDgrTMBS1aoZ
6CFCzSCS01Ise1GsrItaSNN0yFjqDTBQohtDA+gMfmI1H3WQcplYTGaOTXxdISbW
MjQkE7pfuSwo3M0B6S31P6rb2BPsMt2PZH4KsXrZK9slUG1c6YWXyXSI9MANs3EG
2x33YdMgrAgh5qEHSLYhooAjLEZQ5oqtlqeB9J8v7d6OFfy1leILPEFBJ2PNFbzI
spe6ELhFMfRmwyoGdH5ZUifPWWtDJ49j43ipT6DcVJw50FjA1e7OzxL5BWFMM2R4
Q7XXhGcTn+kQKc6aErxAXT54/NgS9TD4Me69sBGqy6K9OK8TvQT3YrtBeioTarTR
U8UBhP3tO/mghShYPinrtcqR4FWSn9rbYq6/wWzRYRRCqyHNSvYfB3xKQwEOi56+
H+OfT9nNmdd1TEmrO8V6MGq03E4cPx1KkR59nl+ok16R5iq+LlTOqZNYm6tLhtDz
RhVZsXR/jCbuXAfsUkt6h6fiMK5LdOtUDtQpu/gxTv+9EXRK49ds3aMtlZVjWBQX
jZa5LX6R/T1Pq9wIxSyaEWkBqe2cXOGRqkVXh+VHwYp4gJfYGDtPR7QfjjiWr3tv
SPPiHXV2jF83mDw8pwPzL8jUsOsxaUsgEpjepcu/fSXGUtnKIt0HPV9KlH02NXsY
Hhd5i7OC3ePsL+B631cQPedD7G6LS53lbCwlBxJEvUC0Qhg8us36qslFRDTcNbR8
paLGu2jP8LoBQPPNeM+3FaLBEieQq2lAUbV4QBpM1AHcBd3tY+v2BDicKjGoY/nf
sT8lXQkBsqY0Hl/F777Kr7gS19IrV3fODSbJttEE0J0dMO2BTBDYnclggc7ACdX3
06/6urEDnorE5SQBQ3AQeuw7mYz3+1VC8adJCj4qqTx1zwV8ZFI5lAQjgjsxwgzR
rVOE2LAbHOOd/bOk7QgExTQ6ZBU7bbevQacfVu2A1ko49JlsUbLvVxa/FtW+LkMP
s3/LChui8wQjIBLGXIyEUZ9joYUU739k20OitS7kSk4S3Ac3XwTIprbkM+00IICM
N7x82tjieJ42MQgCSLkd4QGAFD69+MLysiYIFVyFdLGOmy4kDIs+JJt0Fry2K76n
rlVcqehdn6lvF3GjY4NlBt7zXSXHroIIvYIALeY2P1BF7tQi5QKRdcn7oUhXBHoc
UXCHlckMSRbM7QQmlw5ygaUXabo035Dw1SUoBERFxhoXCNpVk/JMjqv+M5bXXKIx
FUiHUOJ4DtKu1H/JMf25EqTy54EwVi4HFieeGQ4KNjdlyep8Bk7mRsMRwR4YbnE4
vIlkhl/tAy8xcqDF8yfhg1i9+5GSFtX5FlXCCk/px442DUd4Lkul9UpTiICFZe86
lQwsYPERTU7uvQNxPk5oTRrT/Dtr7VtiIAS9tlqGWhuGJ5UtWtMWK2pnAIdTYV6G
gSHUIP4tVlS/33InCXJNdXOlVKOcd9mox6CL++aaRDRNglLml+KAWt0RxjohggNh
DJYK3YnROKEtouF/ZTBamKk4ap1w6FtLUSQ3LqsPz6p1KA2G9KMkWYJ2Q8dtjfFb
fUjQBhRKPJXswq6KlFPEr7W81fbXsh5ShkAJ+NAVo/9XarJhoKRqQteYzOAFK008
SiHfb3Gnpy1r0fx1kD+tvccoAttr5RO6v3XT+W15MKuyXklO7IhmxrbosfIjwcoR
d0e4wM2X2PIkH5zWVAB37/Atjw/r1nSUQwWzLdL9Emxre4Nq5Lsjza1ITLyJEwHX
F5Vbg2LTkCx85WSigW3JWxi2I+HdJQFC/ruP1CpCS/LwMCy9oEUJxLwLwIU6xhsN
e3OCSPWi2wOQG4oTPBNjia+0HiE8J8mLxc5egCFa7kaBBJEqkfOORxNd9NXg8oQA
P/2Q91mtEVssLc9l+aFAHespT5n2voJHp/o36D9lPTGQut2ipsm60a0ljkJUO4eP
`pragma protect end_protected
