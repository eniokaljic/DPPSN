// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R0NHSgkW3U6XoxvfxJSCusklHLpIlUtsFF8p2W+M/6zxkVFVLWlVFeJtme20tYDt
oPwJNK8e1yj0s3DV7lSzZDW2/bUMpkdVdtHQwV6z7wCadxOFnx8UsR76AkgpGLu2
kpYCNeHKf8nmXGHWt8tdFse9RAADZ3GeQvaB54oaRQo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2352)
Nnm2JMMmgi+jmitnwyUmZ1ICNJlQNzD6HQLcD7BzlOpQPB21PU9V7rVN76YulViV
vMwU+5rVrjTSPY3VMeHjghc6NBdQIDtqNPr8jxN3EUBYZMzrlZ2M3nlHq6oPpU38
XKc3bmSxJSzONG/Ok7GKu7Oo3Lbm1HlGedc45P2wCJtizghC3fUaI6PqpD17/TjQ
6oe2nvXSMrS1xnSm8tLB1oBGBjRSGZyTnC5ZUkcLAO5wSV+PEyMbihhnUcKLo2dW
6hgGUVTXijKxrBfP99sYRrZVJufCxh+ZtSH/1cmp0VbYzJQriFMzto/BlxWFe1Hp
cEqVO4mHzwSh3AV9O6LXxon9fgQcQDuiRfnLF/fi9tVMfEz1rLDIA7S1j2JqJMpW
NZTtK5IArUTYL3l6t+sBbqUN3XIfL4xkK4bCgKhj4Wk1HPcXdb0valbyPs43b2QW
+rqD3CXeS67IDjpTGGg7hcBPnegxKxL8+KDYBx4GSTdgnH+xz0J6P+fyXYE0+VHW
Pzpk66mJhCLeYmbC2WTMZpge++9kGvUp0CKOViV3RidZnXdw9muUj8CiUx6KSz9W
ZHwG7/qut3eEXHh/h5t4nvSJep9pDu9iUgIYJV9GBG+QisZo4WXt6cz8gMNB2mIZ
B9esRGxYmbSz/bo8GlhwlCQDrBqXDQlhWOeGQfN9vpygRHJ5aJiu0FejgyyY2Wt8
Kq6lzXepz0a9MUiNlBRgfe3VRxduu3KrHui2RhEb8UpgydduDt87ivSidVWOI8Xq
aQRKMOCxSHZbHiHq8YZqN49KyIyK54khtEKVLYI1zx/H4EvDrqOkcYz/fGXMdMSS
Kg4vmVemOH3iYRS7FycUTnWCBgcVMYU5d/yuexMCrOJPjkaEjWnk83m2O9ZIIjlt
08ERpvHpfMQ1c2jkc+X4jTPWAH9Zs4TJ0lkNpmrbOGfrlDi8JWsDZS6XYlD+A5lI
61Wb+jqswSyIsponS0lD3DzkXnM2imjqsnu+sPT60twk9/4HEiN8xxgQu6FmfWpd
YLO/NPcjuhOm3lZ31XCTyOZssr/bOnmzWPn8nfqMxstejPB03T6W9PZWz3CECf/c
cQs+xKoYZnpPbU1VwuOlS8oRnYvJ5kIN1DwOBMsudpLgCkse14W8t4S62YC5T0ss
lYYr4CfgwCtW4mXG53ZGwNowkB8X7/F8sFvFnVCMkdpAqIaKtoG7VwKDwQZTxWyT
pANVde1E/aeREt48fA1TvI+wrFSCuc8NdzQYL7/A6PnB2H9UBnGYOg5OG4oqvbN+
hQtGJn2SOuhmduLfkddmfxOsmyY2j3cvcHYDNc+CDZRv4G8vALbd1Y3HDl0yEspz
QFtuXq+cGxX0BsgkzoqOzYktTVgLCfUXuKtPaopPG/K6WJTVOINYHKPOv32N8+JF
BXhMcjpEetPZoSMdhE/TMrMHFknXFYOgk5iLEuitlj7TZVDLIjH+TN/VinHdCzSY
Uu7slt/C7DsV18d9c+D3FQwV2QLyS7m1zM8NhQZ5NEWaTD3zUgTNq665GBwo0jAk
D4+ZnO+ocyfReTyMCe8rVebEgDcU2R4X0iqmLxO3iFQk6uUk/0Of15kM7gb2+0ky
cgU1SOGOwrX+vAGs49RZgAUzqN8Ge8SCrM/IDdhn18S9qxDOx1RhCK6SQshRzmoH
80F9k5iTxwtiYvghxqWmHHP+M4EnwZD3cTIczW/hUQ/f0WvP6GmUWq9bMiIp7KMr
SLX+jB8Vy7uqLgVzSUrS7bMp0I3EsxLb7R4EySlWoNJo4hTdJFW068L+hpblaV7T
rSrOTOllUXYkJKeK1X2jsOTMen1rAWJ23JFHcjgkv2DHnBMKWomQ/+CVg1fIAuPg
F1GoD352I2exnUij2L1Rm52a1IirLNi/DmWaQV6rmmK1gS6A2Hc8EC7NMmLgToRQ
3S1YNP5W4WMU8QBcIn6GPZFKz+rrcx7wmLc6LmrpdUshPr/xnKFSQgzYegAu1qOv
AfSo04a4Rq/iBE2BaevS1FPwTyTyrkAjwgWcq+rIXcKmSKPjSPuYtUG2cLyy5Us2
wlFmQw12xMminz36RI6KR72xUtbAoVrntwjCcYsKt9BcmoRfNddbRDthGK8gui46
4DkmF4XLKMsjvqvISsWHHCpl7mMezPv7xxUw6G2L55/+vbGmBjxWJQ7+j/PABVHt
NsDILCtlgLqX+bHqJFOD8UnAhWrlQmdlimpM3jRSdL0nqkTioIRnL4103n2vWx3q
s6zWfi9pTLdutLpEmbYqwytwIuSCFYKTtbq8SmkaXK4KV5YFbgI2AVRSC3vydqx9
1dCQhkuBFOHyOJnLKwN19OYfLsfJj1CJPPYV6Gi4wOymdSq4IWRMMrzOg+IBkovB
SlVtqgxc0XnquiGJNG7ZUIOQ2voYaeGMWm4Tq38c5xndKYIIbii4FXW3yNBz+0mq
9Rb49NSbWWNohlaz0EA+ChJc4RqxEbeblYVsyvdfLxz09b+5d4G16OtmIX6xju7w
/lqEQGyRcgZGiwI0LCx1K88xz+kKPXC9++KHBti6lmgBYpjCwZ3LvITnszhcUxRF
lh1Fj6Lt7/tHSEOgFxO+VUejoN0LpUOEg0Va1YTIxoo+wlbJ6pXwgGsf0oQOcZoC
t/VwCUoQIN0Mxeq2Dr6gshuftAi1+6a1F5k8GE1QzMz2hvtY0/L+bj8dhdLpfDGi
sjOflrVYQlDeYY2ETlvqzCe+hEfhHls5lbbwTuLfa1aZQD5S33pjjMLrV8BH5qUC
LewDU/AEPae0l1fO2XbTXi/oUdEfI5RpImVr+79UMRr55vg5RiUvce+bgaZaxUQb
0Jss3wU62+7rjSW406S52UsPiRmCWGee8uj5fkkNqaC9FYDeLebLN/h6tBEop7yk
RjFmnL7UVYV8AVQtDRYj89Pp1fpE8GxR65al5jaeFlF920JdZjhhhwCod6Slp1Ft
I/XQotJHz6IZfhTXRKDXpSay6jS+wj9wHTpj7oXSlUnEMua4+NLjZAyJBsPlx1ng
6vpw5WabGOka3xhy3g2jOjSLJ0yq8L+mthmo2yAUth3bsCJuLQke5cQ+/avpEKsL
NEheRdjLZjPwGlJt7enqrbzIZzgVIu+8hn2kmV8eBVEZCuIZK/Hv4LwyRZmA53op
`pragma protect end_protected
