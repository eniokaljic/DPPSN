// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:35 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bcIhK3N3Rn8HsHIYZD2LVi9Gl2iDKvLBXUg1bySE7VhwaLqyGd1CuOk8duE70V3S
3rmBuVDxwEjeKBax6eBpDCCjfvj3H1TiGYe8OZrfbx15DTt4kTF9NEnLfRVavvHT
0+34+IMA1JN/Y9OgISqjhuHc9FxXcgozJue6lcZ2NbU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27776)
Ly08WY0NfWMmlFfASI5vNT94+/PmDucIzhNdr32ej+4hzUw0nzzi2wX/svdCOVHL
ONijovWF6jzw6HzmszwI2JmSWLjz12wI/yB+dNweGlR6NbQddFEwqb7PEiaLCu2J
ZBxWapI8Jt56MhXTC/Vs+Dn+MA71PbSxwpf3SWGkUPDMUKPI6ItyvJOTxTHyLL0a
yY1TgT1ZS3r9P68/byXZOrnaKEZIp0/5WIAHpussTG7THikuCLHnCot9NfHnNjTo
W7/S7YPx32BoCEBVFMhLXS6cuTrtDbMoLDPjj/PNF7jkU44mbbWmGrthPtrr73GM
0xgr7KJzWIpfapQWYpiquvvOQC8ycfSd03Lkf8rQ7ktTb/zuG45KveVGIicwbaV6
zkvy7Af29EliwBHjA9he6v1hAW6yefa620afV4e8ikCQIr+0QQ6cGIeZjEjorAX4
Bu2VsJ+Mkchl7Iyu+5IusLOZXCMPN2d6mXNqu+8CYXHvRC9gGYWAKA+OJJC8n6Lh
E0Dy7i7qs/lhb99Qvx4kPeA8sK+R156XBFZQ0S95Cf8JHelWPQZjNip/Of/tLeMC
w4oQ9MhsXd9+1djcnocjncAEpAWdrTpxBAK5GXkg3jtY2sm8+gxcjIIyiRLiZZmI
Vkwh8XWtTnQ8v05Sp4PVRuz89poqfiZeAHzQIK8wIqOIRCohSr19voGIUGt5fw+l
aEITmpvcQY76mgplwYlAcFltngtxSnpCWg0BuwLo8kbLZSYD5XwhsDnTB+yr/GE2
DgbtREu6N9Va27ibbY/wvPM0RvN0MPLBNbM++O/hlYGxT9iFFxZBjqSaVVNblW54
+4JsiaizaiTLvwF4V5NlPI8FZ1USh6gq68D8vA9spB0JLMwNG5aqGaJfjTmH6jXe
sjEdNnYyl7RqKopn0B3EjjK0lCV6f/yjFVxYAz4y0M16rTLWOiuwTn+3FB9BSziq
Wz/8Amy5Jv7+V9XGxefrBg/uVQDz4va/HwnJIX09DFPb5dv7iQMv9L9x/rHmZnPX
9gKKLUJwtsCP2C5W0T5MB9jKTib7UNGSBtf/Nz7t7xkIO4xNBbTS0wClkgMCsLk+
I7UWxppgIq/mAVhtU/FOl3jpe2uzp6WEUZTlMFZhrbkaFZn08MHOsq9+bCsElait
rEPlKMcYFwCU1bd880GmOrpzJKpNAXmPkTFFezzHmY1BJABZE5Ib3rZByBB+k6tO
gEOD3CoaY69VYPk9sAOsE0OyEXVpW6rwLi6DR9j5kzE2w2YI6Jd89rTN8vl3ChRi
jwPkRTolOr2GPfOZVD+r6Vwnj75pH3lcOTQq25CQOyl3lLOdg50Uav9SA9aW5Uez
83Z+mCmuyqoiSXFGhqv1Dv6t9/qDGUS+rsoYP+5bR6N8Qqh2m5VsOKvgCtXAbN80
P/g7I020bgRUzWOQeELZANpEm4sQetvmItOH0us2z8oww7FFQfAugfpyfXenun+I
Oo2gwTlEuNnkE7KT4cVDHTkQQxsPswhadT30x1vh2px2KhoeX1oze9tzXTCI4H3W
OsJ5swajSnm8eq3fMr59Ahn4ZjAM9chn9Her31O5ahOZoC3Bts6khpxSz/K3CNU7
kSO7UmHL39pPw057YeWScjTf07Vllt2l0Vf2iZlY2wg0YprqnaxNcSsdPVHUGBFU
hw7evl2T9OFXowBMAwXp1fXvpi/lIhfgMFTyrV323u+kZMXoyYFYPbPzoGgTkl9c
Bl7cZCjOKs/QEHzc7sbBh/B9LC4+snP3PQJgPg5dlRlV1Kfmlm6IO+3Eg076MSU6
pm8NRHvOqWYDrDnI3CT7xMgIhAqKWlUoXn+bXhVb4x7d3gD7Fh1LJEs5Vfeny8zM
zrg1sulKElpiisZDtsJ0N8pyiyNsRkxf/6l9GCt2r7bicG5SEOB8nc/0tIGyDhND
3ItwVsv3dJFACCy9zI7CM9G7PXQNlGipZtCeNPfb541xUtV7OCqkkln5B8v9lWSC
qR98Bp4FJ4ArDmuf0ivtrOVCtaDnSqcZ11efFvBFq4xBFT99IaFdXe2ks/38ysH6
CuUQBLKu4QYA8VZSjw7FH8osst9N/STvibOC3fpJXiNzaAroufmQc09sy3Izqxro
8Kddt1vRS9w6mvmwo9UBIROItLo0VSCHdNypSQkz9jPC+WXUMk5hZFLmnNdic0GH
GERIBCyByetwuqjbCJHVeCiic80fQQwCNE1yEXZQzsszCPRsv5pp8ahalYecmdcW
/wNO/5Zyk2Ojyq7VxUS5CYjwe8G9ShMrOeJtlUQiy0kEDwpmx5q/DbKI6M4kKfiY
AArSM3+nCrWiS586sHoKAeH+4ut3IHWJN2ZYlmI7/0iOEumHZ4EGWI2eL3XUMlxn
CePbOiGt/OvCV849zInoU5GEUMeZYNXTXJdS7Hb5SXiPbVMsvUUehN3rEzb6hzcz
P/HHvbHOWR3zEAthmqAI1T6Pyz10umRWBmDp9qFHsbFbvipY0exOjKtu5J9X8N7+
Ie/5BGGTARA29F1bCmV2hO4gDQktajn6N6y3Fq1pswHN+a49mmGUCXyQN0x9f4gl
ivuAP6p3UIb10SZ9xR1h+oT5Gt9XzJHSqb4bTFswJ3E8qmw21K0bv6ceJdZq05Re
nAbvbbayPj0f07r5G/EjsTWF115HUn2+9eWesO3DMBKrvJVpCsjSf0ZDNE+P5rj2
kx5bGjCh/kGdk/90RMiALydDjKh9Q/pX2dWDwdFVnlNGiwYEG3KnZNwxGCaG7w6U
MwDnDqSn4IOxBvYlXWeb43a5V8FfjMG17ljkyMTsekt6AvsMxiXJqs57f099eNjV
96UvpbRYFOH6TDblhuN1+gt4hbKAtRicHHwqVbzzfzH8/d7Of/7Kg+pMRI7mtD8O
UCv8xzLcWGWKNi95/mhWyrZhjIcnr36Kfx4MU1QSowsH8TxDqAPxs7OaqUcpGetJ
whG9SB/4WgsK9XtngtJjSOa6980DdPM4ts2k/41C16OSwkw8m6zElpygiGc90v3C
QtxAVdESlYWUsz3+kAELGQbVtYAIShObhCFCBWgnBKsFg8h1nV82pta++Lia127p
iQUW2iQSSuK0jA+za8tFa2jugbdeo362WWd7rnD3uFgWoyBfCJSCoqAei7Iv1E+q
LEu6vIU/TaKwTDYoyVvaaZBjsHpxHrClUvmCnOADHrrpFkyWPzJ+1KFI7CsP8H9K
Z/hxkNo2DFEos7iFPRXFz+2e6RyRZ3I/x8i6DaTidZ9+CVVFEWsMZf/QIEMbySWa
R2m8GsxhIdEYIsU/wloYZLTkQdm85wQrfUxxGo4lfKXyUy+JBYQzVtv3WAJFU7V6
e3zwBTLTNVsiVcBkrmdhgvuxpIz8ZO5pMOekU5Q5Fi5CSfLAabiVU/9PzRTKOZlS
IkOQkV/xYOEdlnykYqlEEush1kDGKXswbpgE8bvQeNv8pzHe9foi5dC1+FgizPi/
QSsa9zTeB9iyeyurYCpxevg7CF5wmeqMksWurIzn2xXuy3jG3pFZ3RhgVVKKUvEy
zdVrFKhZXp+UWEC+pS3Q7Sr/dl2LNwbBYUCXmld4UFDeSaaBuzZ7gvIL5Nv+DC4o
LexeF12MosvRBB/QAJYP7h/jp6h8X6JNRn90/rWhzOHUVWhL2i7m3RcTS8qQGxOg
5AhWHzxAgB263VtmgHoCsEh9/6OtsGdXkDylaHS2AFSnTtdVg+XdqT8yUgJbzane
ff94b9daIjeZVsozlOv6QXcQFPstzZY+gsc9WjfSI0Rv9Mqdv6qjUQ27/7cEL+3/
RVORobWjt3T7pM1cgAbHagEVQkHO88IaKrOAjpLUxk7mUG1PH29ro7Rf1ILXS+6Q
UERjygvqSSSCTPA+0SjXzLLZBAGKYXZZzCneapcXl/mwyOcfby53SfgydMqQrrQr
shD1McDsuNLIDYi4dU+K0DRP5bj9D6hHaCFdecTDC+LFqy3MWPr3gmEurvIToxTw
Im49IA1Ifoa4hfjQTYxFEmPtHehwT3cos2/rVSMqZ5UoKp91d9nmQL3GmN72Gui3
IA7EtGcqMMq1ss40tlg2t6IQMYMrW1LEZcyS2Sjmv7EV6h0K0jVtRxwYraicggLT
UVXsQDKAgrxMkQCIbplUwqzNYVt1nehYu9ZkIxNb+1+B+sHaz99dpTwYGEUz00G8
xdzIyVLcN3Usdo1OkX3DpjBTvfVSVX0cC21deW+VW+8xc+NQV7/x2YC497j0EqvR
O1JZh30p3APMM3/xuGuMJoN0znRn7UpfG+ouVkEmi9KWozTZK0CdFYGK1KNIp60j
/qbT/rKK7t0Y/odQPhqyF/uWACsE8xl+8EC1YIiSTT2iUDSE+dBfhT2e70Y5UbgO
iULzQiY2Ptex9QxULZDhC0D8YYOTLTZ4ey6RGyu0JvbG9/jIuVhlz8gO/w/VmcVV
cT/SXVaNNzOHHIGRAv1Y2HFLCHTGGruVnzsS8Jg9g5DbrYVCFVjOKlx8Oe4o8NV2
z3WIIcJvSDcIuy4S6NhYQitw7aGLZd/qmgMN2havbiOU4M5H3IPiC7TFNjbr8eRe
RRYfasP5Oxuh95mP+9vS3cJQAXYL8ATNAPpP/AxYMw8aEPWNWPccVyQ2vtEOuJIp
YBRy7qUVnTpdBSkW8jHOZiSpEPK2cyoqQG1zCdwHwkHJsZx6zBFbEDQsoi++TtTe
oCEDafa3DHJgo9e4CCFwqyEVHRIVHAFoEA5r04BcoG37s8AVy+AYMDwH/9JUOYDR
kr8Y+B2reNNZT0Gl0zxvFXUoQz23BUUCrSZptk98IerGFsU+F3qdtiehutggsHAK
X/Vz7NGanTEu/YdRPhuZfYs5JKDmsYKoECBWYwfXW9otn8bqzDtLl7odvxNLzNge
UWIaTApzUilkXZi3UXvNuh9+kEKjMefjCkJ29Z/VIdskmUjZWitniXMoFYdN9hNU
F2cbobmOOPek+nES+vw7FsH8hw1AsRt3dXIzTMB44tzCsy7/O9TNoDq2mFb73eKY
ETL4qusRDvxYKwuWcJ7OBPF88tGAAtHGPaFA05zRAi6L+jfxYryr7ubyASrMup50
GulovLCHb0E7bw3Ggf2uf6dN5SOBMbezbnwiIgFiGKPrERYpG4PqCyrTruazVCdh
hgr9C+Ee+iOfGa2T2u3cSp6Jt0FYvZrbowJHyX1+OaTSW2POeuVgWhexPDNOHLcM
OyVzonsBXKreAeBN+YjhG9kBe2+lhUs76KXdX53P0LUGO5AWlvSrf5TnBACjLrHp
SEMcaUu1FKKZryLcRUqr47pCOuvced1pJkr+pr9QrVczyHBmPnd4S7qN9ulKOaYw
NvcpcTiPvIbhNCPgApnOPK4kBEoRpzk23w8lYDihuerf/gQZMZzoELx7E9VPZ0+l
nRa0452h+Mx+eWMtmCqKdgfaLPtb2sXDG7VR6XtGudw07spWlnSXaww4UVfAkYiw
1DxZlXteZdbg19EHeVpliN42amzNY+IyxpQYx01idBP306rU9xLpVy18OCUIDSYo
8hKK7LiCn03mVrnU13oZA0F72gXYh1OMhY1Qo4iM8pG5yBcF30NJ/Llmh6QSdgWH
cNWhPW62Iwi4xSM/rna7DNw530I7z/NIJXSjm1uxDlpApkRYifmKerTXg/0FdpX+
Sjh1OEOcodCjRqKVYOzlTKR8PJqRcU2jQt8M6DvWsULtL/+iXlvsyH15ivgOKEAZ
S8Nyg8uETo/KNEEvltZPQb8sLvD07EiaXUUlAiQmTpilyRPrmBC9hOLsr0BsvWdb
96FM5mOztv2DCGdyhj9iLhXTojC7eJRpMEmFviXuSH5yjLlE3ulx6ey8X1Mdvs6q
rhQWoAwNKHXtTa0+VKVy5DoEpw0XkPwyASCdt0PuvwcJ/rPba7HkQVhNnlBndf23
fx2rTq61gxzdetxFQYWjUC0GEtBCJ4qvmiUptAPoQDHGJdzqv7vyEG1OtJpgloEB
FJN2EQIdwyIeHYm3js7B8bBaSGz1wSsEBEmoVX9WKaC+E3kCx6BATpf8G9fxI6ew
KM4NgUEycjMwGmqLTJJdUfPKLYXDhtUEVVdWRfdbkKDnWB/K6yPKvWw4knfcFtFM
AJbiyYZO7as/3EfT1cnGddfBPHqMCSstITBPhofWFna5qgKo1KIW9BBcGiPGdC8E
Do4unWE4R25JW0GDIvmR2QbA8jURUIq6YZnobTOPMtTh/a9tctjJOyYCak/56crc
kNyB6o1txfPhDqB7MzjEhduLN4uHtfzlyXJwj3xDZqUFZdfyzHkn/FFLdR7SkuQC
gPfeU8qyTteec+qudMI7WP12DLk3aN/RJAhODyNG2sWjF6jBknyoOaiLSH4ZtxRs
IMk/+V2dH5XRTtLFQLBjYuU/lDeb2hWr/jIkw9X19GORcF+3q0BBc5DBR2ib+MPV
ydFCLV5kWXVTRQA+kmzqk18pUZimqnrPdDatcmkumaE4me+GhVXMfzInJ2lDHNXI
gmShyYhrx/8mpNVesocp98AZfJ+GYC/Dx/8UB9pFSWQ6MzSKL3UzJ9Z+CNrmsZel
N+php7gwQvEc6Y/RP3ze+qbKa40hHAj6tBWKCMFS9BS+BSlguV644QHmUcrcZcht
84L3aXfg2UGzqnuOQgczFRzUIzOkqUw1LXFKjRYLQIGwNkMRAiZOgVCAp/zIg05U
s0wlVmMLokm6OCQ1prW39g6YjYKaj5nAqWcknID2gPTMVK418TWTtca0pBDfM+Fg
mNlDTOH9Id2XMv5FrL2hj+17QOJEDF30RJuFLezHfXsDil0RCPTD4SfBxJEhJAg+
9TCT+WBC7vIhNWgn47Cc4Ub9OPhogqYvtltW5Wpw9FxowJ3kgphCxhPXRy0frthm
xCgdpMAX5o1gF5NFXg7jpZSU7Y14npwXP8c4hq3Z2fQHMI1nyWA9kEOy6kabju6F
LlboKEf7K2ROASfvjTJUM6s3k3nT8UYPPM4xLv5ffNHqKBXs6+DxkYXGSj3TPBaF
Kru+9bcRJp0dc3J6Bh3editNa4XQXajDJATeA8WMLXWpvtOL3gJedX/mATCpFALY
zlwOGenBWgHULypYIIOgcHE5HIE5SbJl7gjN+kPYFnObb3mi7MBbralB73YpyZ5W
sYQp05Clss6PL7DKCS4jRBNy64NoKNe7ghXAihqgZnkaCw5meB5Avp/Wm9LJxfX4
efu1H7UkmzDLr8kYJ8Z6Y3KvaTLjMxoqu56Jvv7C64zlvNXoUTkwcxO1dOLIIlh1
ICyVcIPoV8JPL0ZxOAMmLocHbEniJN5QZnNPYwfzRiGbL7UZAgF85eEpyhmJqgDp
r9JC4Cu4jEADnhsj6qfiKoFYdmEcI9gSpxkHYexxctFWDdQo0FjHM9IQVwIVS2cv
qakwH5vF1r4+ZSXXAP8W/rO1L5ooozNojvCkFPmkB4k7eovoljony2q77GmrAzTS
cukm82XhiaOVdHi7New1rRQ1FoK+am4/Gmd79FUiSt6RJThYGqvGnm53RqhFc3g7
Y8oGrBbPfzVpM857bvnR+b2+GnJGOwstdWyEFUAJEQDZdHXXdf6MA/eW+Dh/p8xV
WWA2QaYHWySmFYtzSJnS5jG0ZVOFDfSYY3EZ3kNzo42MlMQoHzjm/Hqr/YZCmKPU
NlOH+SJ/mzkTArzulzcYVOYKhzhbUkDLRuSVLNNil5w5mj7gPWf6jOwlmUNZWLD4
bTpgOSfpdRETB2cTQmwTpm/lSTCCPSw+l/nfn/C33kSfl4D8BDDALcgmB9PK/TUT
r9eBaaECZJboIsz8uoRXqSn0eVcCzxv5CkO0Qlter81ACKVZuczQ7XI6hqcZoV/n
YZS2jdSYAi2KEI51Ncld3K9xHlOGsf465eJQ7bKenLWhGxXtfutK1+dT0I0aG6BP
Mn1FlaNYE76zGdocKQlxr8jl3Ux2IBkdgNZFp1dZGHQcFC5Su62jcmrH/NdY9cDc
U45YHvoGC8QLbhxp+BYwWRCWAF5vMAT55Pav/qltLOEMRl3fbBwJRMXpphzXRqFU
IeekazyZw8VR4UG/uuF2TDWdW+POj0GUX50ouBOgRdKtw9gDeNvuor9r5GmW5ASj
btEP0E7CA4eh7DjxIo+D37feysTVIM/1GRLyoDtZlET4q/Ra/7RyY+f5rD17Tsy+
AVYBpto8ds0zsOumEghMvgKJOBvNiGkX8vUeYrkI6H+WAapfhWEXf1ktD5l2FzCx
cJCJDGhFETewYQ3rhWkyFr3jjIDBTS3RG77aTQ4SsUDWncLM5LCBFtLgVl2tBE7h
jSixN7aTInGkhlp2VUD9kQCH2JSZq000jT3sOBp+eGwuiPb4pOvqEExmSrviGOOQ
UXmWqr4wnU9bYRdNxAZiEAyzzHCLuueXNNCnWPP6TAx8sCOw9qZ3iy7JUlPTxcoX
832hw3JLANtPAIh1d/vCjHYFRooYh7uffej5NehI6e3VvPjAtbbODOo6c97N5434
tCG2UiRfhdAJ+9SIPbIl9wlStzz5dLqnu2u+ZIzB909gHlAvXpeklleHO7puCp1I
2xnntWFI0WTVr7uRMIW7/eU4oLnfQgMMrmZqRJc9pTBEhF1HSunqxQqTCdyiEzww
p72pCie11EyG83RdeyECKuVUfz5TOzzIpn2rXVyk7LCRda3vYEnfqIvomHBKNyF1
bRZP9NNFmjxhvNSe6gQU8vaMI2RQDMa6BJmi8qOAc8YZmGkfyAHLsRfk2k4O5xzN
cMCQBxrhldjzCqd2hvSdqba9/XhiUs0BW4DkmB8l2jyzlRbX89+nF2Zc5iE2vQCD
tguIXaWysM962K0cPwg96jgRMcoUwFYZxMixD45R7z0Ei9cz6UmSriNRB3J12oHj
d8EOYPDszRgU6/XtNedopttwQWTGnHM6oGRM1SKxwEbc2RqJTZowByW62adM2mkJ
HyKnzmnGicpzn46sbn3yZeM0VM8XYApqCdOqoQ4e7+QhmDwzj3TVAjwNU6PjKjH6
hlVqAaKGqLc1fvPmReNu+PbHn3TgBoyP6IlPLjb4Gfcp/otahrXcSEbvTFf0s5/F
zjs5QCQOT3FNspYnszj/K+13dfRL/59YPnaXIq9N6YwAbXFVsZT1Og09EipnIh18
9jQLbJ0U8/+bRVsMqQM9q+URlO+vZ0JvqsTtaNRg84Lv6ybSkqhbQXfklN4dNcwl
Hihq8AbJMmRnI1oakwoJri7kGtoZiR6bJrYxs6Pyr1ILFv+5MjdBefjoovfhle4Z
NTU/JEMiuEMVtvlUk1hi2LnP5Z9gpL7TB2uYf3csw0kPPvib7NIM2PhZRfeDvUAz
rQYv5qms1zIRF9WLdY3wYkhOMcXZxTb5YUn3WUkPFgdKGjP3+djgwEhbZxGvl4mW
yMlC4juak5OZGJVwpAbridiNoTOZlVy9F17YYBgf0PgFok3/qOqPOJk8zHkwrna0
AJy9KqX2p0/6ktk4paTnZH1k7sUcun4tkNhQjBsJr+wONttFe2VUfVtLuxlPcyFU
OI/Ifpa2DK0eMoX20LhqePvIR+jsuIR9y4DnzbrR8kyrMIybZju5CloRPyNEpOqf
WmHQu2Myv49zLWtubMchd0WXQcWDmKLp6b6/6u3jf56yoAwobsc/vi/Edl/0puzl
C4nRqCJKFDX6MXxdb6BgKXG6e/4mFEJlKnTNT6yuhjoVxOtmma6j2YFR9FZGaRx5
xrC3gOApTSMukmlx/h7MIz4nc8G1V1U3Dxb/21tZQvgzjsxOuXFWRhb0wMwg0eN5
IQZe6WQUxFkCRDzAXNbUtNBwDU/P4mUGdH4XvCHLi56zhGxEANIqIsIKX2rsiODt
8mCCpiD3qc7e9Tw5XG3ymx5jBr6xG/Sij15xgVU1xKuDf+P/v+f1DWIvBHjJSNel
jmurdKQyQ6PU2zjbfzhGeC9xBlSeAfv9M+XG5yX7MvRyFkbEEeutIss+wdR5IXVQ
E+8DHYyxTSihzaKCncOLd2SBDnDx4xDLvod4QG42c1puSPc1z+Sdh7bNZo//Uzlr
zXifNVO5jf1MpQ1T3dOhqlBBnPZhRyTRaUAeE6pZ0RNvoLUbtQj8LGyTJxlZQ6mZ
YcQtFHvJ1/7Dqu6/dLsZ7Qt15Vrc4LcDhXZU1vL7OxBBx1PkKfR+a2qBOAczCb71
VHGRla8TC0qS+XeThRIn5VU8mQ3OogVlnsS5UgXFSlgxN2d6XJ/4D4kBAZ0IGqPX
weyeVm8WVO8W3fUXtGWle0fZhGfa1q2RB/Tuyy+pqMvpLjMaPsxFlmkkKrmQdfYw
JXXZ+5vTHl1aFDzF2iDAReuu77unUWfmWM8bCd7JehJBKRteoBaS9Oc9zaL3wAk7
/f3p2V49s7lsK7kh6M0FS1hELqEj4SzMIPdUc6p69NkukDvLy5pSPQWUNnhYgse2
9bY+3Y9PpXBQ6XjBDo2olNTtTECRfjNq1DVvNU8JgTE+xUxA57HlVAh0C5umAAdx
Wl+xR4ndNLGtNOhN6Rp1tqkrLrHnmN+IJZPpmeBsgqyCL9ocdA6fuNuz8TI+fCbf
oDVQeJZ+sFiifXv9LksdcujYbp3CVbnJtYSRnRdSm3nVvbW19r7oFKPHK4QjItbk
Trao6RjJSjyRJWHJpQdHESnZStucr8UvkM1PVw0pZc2ZwpDRz6BVuSiZTA62R7Wn
GGKV/8Jo6h1bmjmwGUGeP+pHBrKR1E8ZtOlQsYmx8cYerle9lubheGvk2xlXGiey
5hoxvJbBByOzaOLL7E0V7MZqC4puxDLaugln/Q7nfIwPGd35afkbz6LZtqXAUB8s
IluGVPSNZTTeTG5mbHfPCfvzFS3/ArlGN0VDTtdZ5kL9QGbVHkAuqm1MGhBgzL0f
otbCTE8lq+X8SuKNFhc6dObBWL+3r0tIjSMuVISTl2R76tIg9kDDKw5qG8JG4dfm
P6vEqXi+sRbP5RX9kzNYGFVhz03eFNBUeFAMQhJVTaveZYbYLBbJJ89CHOhyNRFc
lEgzInB4DodFyuuvWiA1wHMyiDeC4gPy5pvoKWjpcCR2t4b2u4GAzjDB87m5VZ6E
+r5RCIwQBiovn7uwXU84Ue2pqPTK+Gq32nc1qhtqaNeKdxpkx8J4Q5N14D6LjCKk
zoNmK+vWJxoQgO9IIU9kOlX25Ap9HRZeFLAIn0MohFpUipPPSQ+9FIOhJudW7Y5x
U4RyJYTM5EMvJfUtLNstuocQwVADPBIO+G94Sdv6S3aDsLAgjmzoIUN6ksBm2xWb
2WgXwGgW1sVn++wOZoBpRfI2ibk0DGgPbMUSGB1F4shSQmsFGa0dEZc8/2MHWzyo
Myeei0INaS1lYf6u7nWgrF+u6kLaED7Ue0PR3L4HJP5Ahzg/fg3foNGU4RGai0aK
8DwE1E1P0yUzc0aX1k3z2QyFWukE6X2PzT2AE86L4COs3gQZct3i8+NFmO49SmuX
0ulAha1FibLGwIKGIpxXJ4uDM9uU+mwLGcXQ8lsmG+r02oLDjssnF9LBZH1Mwovy
KxTJhEaq6LhFQq5TuIo2wjnQ151iT8aRB/YCceIiaEwh6KHvX9VU8xWF//41OWdX
xqlUaUTTW1pTp0yId/dLm9kLnV/P/CZYs1TgsEFKQ85I63bzIVx0RMdt+ikm7yYB
rt3PIbbCMJU+9VE+cmD5w0pwy7B/ipufEbRNLYLdFzzCaWjj6bKgHt4f55dALsuB
CQbnWzaXF/Pj564IH36w+OFsvfZkBZxZykgQu3W1TayuP2Ny0YWRF/1IhLXErEqG
41fCtMBaFCNygGtsT3oGBN/M39Lt26uvc3NcwZ4t/9LE4dbaULZlIbZggCah6grR
7rm96qVneQsUN2C4yVghBk1r+Jzd2sYHvCGA1E87FBE3k4wEQ1vD6R1tQy2j+7oj
EIkuyQRrPKurM+MTgQCGXlRiN6fTy8lCTVYWX/Q5Z2KyxFtsjULX/sjxs3fRZLeU
vQvc3Favj5MdITqcpR+OoDWJa6kCh9AXCMPahMj/Mrh6qiqKV9aEOMyzT6oTl0rv
OpQEudh7h37QDbv4cs7yTjt7cRrMEQhr7TP+d48w18JzjtCU6Aq7yb4cLl00KoPE
okvk+ILyL95ok+O4uqdsOAk2ltrTWV/dgz7ZYZre2QOhLYxZs7roU2ATMqUNT4V8
cl+C4HBRKPaDj5MMiEq+z0QBZT63M13yFt9glSTq1o9g1mTDpnCpkBVrAPvVJrOK
5eRv6Vg6+PhGSzYGiJzyTkCTv5VZAyx+49ZRgg3oTbX7Q0pg9EexSC4G7j1RzXZ4
I8oBYt5UbF03ksvVQEgyanXhjYSuoGdvvUuPAUra/yNETwJFEcR86E9FIGyrldNW
ysIkQdn9koMZCvw3vJ023Dd8/bH76ALZXYFe39q9bZzHnPSnocv9I7qSEmFcYs7g
rMQCPeKRytUR7jpNr3vCFbeZs87dHf06VrBCcBT4R+14iM8iIXi0FGoKT9ES099W
KgVS3czjLr3Pj15ozePe+aNS/fbMZmnsR8uSxlH2Xbj3NvnjaVOqWg5lrdrqcM1R
dSxsHiir+C/cORwtBIE7DBpFbseXY5qKQqZsC3oUNFu0B0txhX3AL0PTybIkz1qw
utRa7Wzz3AxktX1ApQmxy05NfclXwmc0SRfK4ig1bE6Q4Skgr1soQKmSrlvHYeVu
WFFlkCVYwxsw/dQgIA2P66FfMBRmL3trUKDbOrW0uqbSDJEO8PX0hpKMAAcJAlIn
zo8h3WH29ubxfrPpks8RBEdUrTdmV607CUpwlixJ4oxjTVsfz4lzpOhHCwgyIFe7
qdscT6HCumscw54qu9d/Z46Dn+BWHJ74dUogSgY79Wt5O6HV2nQJZLtbqyoJe1CY
JvLX95eukmD8RzPvbUHQnHVZ/1liFSWkHIsNUJ2GAdUCRZuxKJegfRHsyIGhzCQs
m8HfsT6MHIQhtvIteiGktPVs5tZlrwcyMN6k2rn51AoC5b0QgS+s0OmhpuOXDpe8
cqOmWYH2qQjPT3a0M6SMktgR/N0pz4g3dXlhLit1mUaCoQpNlMsM31PzoaTUAVWs
a9bXpytrlml9ye0ZH50NGj2wInh13d4agTCptsLoq8KpzOadan2RGCTzwLqNzAOc
F+RlM5fl8cfqZ4mvh/wi71qlq/MowqkhBIALaQJ+1Zcz5mq9ZnCBX75D4Be/TJh6
tkwAMZEfBQGQgnybqGn6/1I7dvKtHbkKEeqOQ80DJRNZvpxVPFOux7tGoTW7YaIg
mOd9k79RIQg7Uska7eAXRoxOKW5tp/6owpAxX738EuLVqaYcpbI72tDztcfr+X+t
ga5KNZMy4ySp3GGL0rt+qoWUQ7lmvZb31j8BmDtcXYETXxXUt8hw0RBDDPOnMoiF
V6N498jyYX/US5unMcUXj9kWAtKQjWNRf6ZKyACLCXDPJnQfQIUzUOVptz21V/gP
5N9Kp5XbhTTk04rSvv1BQvr4e9ctb9fwCLhIFO+5sKS/zCUlMaRvBOsRO+ezVmUr
F5Sh6mLs2ilWZzv4i/eqAcUCaQRx6TeRWl1H8tHMsIVdxkeMVWWC59h3cRAA9uY0
lMf4uJ/ZlM3MeN5JLeHvJimEtSeXuU/dvtbdNKfdoJ1yg53qbGceZFg+YGpCqNI7
g5noJ53SAFfoPLEaSvJihPL8cRAMB7+uCFUr8pCeAhMiAJlaWZL8p/ySZBY1wVsV
QxSr4NKKfgzDUQFIYWroMzRw8AJPgajEyHhNewWIXAjrQmxzcUaXhW/7msp3dIqP
qzQ4UWzTKUmgduoRfDPUC612CC3aPLXRoDSigmuxGrnukyUAniapzCd+FK8XgMpY
dH5dhdkKdcfga7MZEUC0/oKBbbxExTyG09Oell+WsEijOXf1BH9g7wMc9GdkzRBo
dJ191I3TSEq2PdJwqOyYsF/OqkqJ6c7TeDftEKB+OYUhD09BA8/u5DrnwcQ9hZNn
rpaRrs51FgIhmOGp2wR1KtuiDPnAV8gAPuopuV0CHCtnnCK1u10spIKVAGgXGkuX
qwxElmG1M62xPEyyG6JYtrgeNA0Cq2ajufM2b7BhIDQzRRVE9HOwKR09YQ6RQWFq
8s25X/P01itoiHIP7y7W+if6H+JF9qPmWel8vHyBi+WXEFfLgZqjH8OdPOAYPujV
xtUVfZ9S/Dliy6jdRrFL/yyZC3joxzSKLO7QkrJD1K63lcc+K9mJofi8s167Dscu
dhGR3pQmJnImNVazr5zXVOPr+VR+ne17MovOdhbzA2pG9l0gnFSnGfR/aX/mKnGC
K2BREdSr8pr8lagq7AZto3DvU8pSuZtdaMtOGyZ8Og/7lB+YtF7xmyZEFRBW/6TY
ifAJOHqFSm6DL2dXc64qxhhJL3qVLDt/y2lzVqypgy81RSBW9KMyhT34AP+owdC5
m4dVYzZG93OgqZUhaDeO+z4vvu1Tx83qloMLvHRuGd2vAb0tuatz1EWuw+vAVsQH
Wc3rkLNhCTMSL+0FzG8DJxUDE9YGS/k7DkdSW6HNT6LFl44HQHARoqsZoTQz+MBB
2dtlwbHY9uo4C0jxLC7/JyAoWe0ZxPI6ukt52g99WtrfQ18JuXimSEiJJky8gjiv
Xm+l/7jjpr4EvEXTaurXBRUswoecaTbyyI5UA7YrC6GxG8LuhDzdD8iPgFRHftxs
8o9AO7qaMW0FzfEPNybYRadgo0iin4Ec66pYKjIiPbGD7dD4AyQEVhBxS18tM1mB
u1QfS+3kCFoCJDO9pAafcygWAXWlicvZtgLXurSDw9DaXVgHEMNQAtn9Ipex3LZC
fvBpp7BGojQJxgGKBqpnFLzAEkjclv4kP9tixpJLYCJyyl9IB1UlZP0XwkPZOURN
4gEl/oBL/Ol56Lma3nfRiVMfRRS8OESVVJGzMd+JoBE5kbJvuvq25za+DLU1sPca
Nf5QlXP/jpBjcnfr/qTdFlUkuAONHfmtsbM94jag4pkp5zVKa+hF+ns0gw4CrqAZ
TMH65rz/MgBdONSLpIfI/BL+b8xVas10skMtCgcq25e+kZr39YkVxIvkpZpPUMTT
TZD6N3lldbDAScZtYprPhegCa+UoBiA4Gs1rbFKusreIea1YZZEYk5Mo9V5UYBHn
DfLkQRjYRI3uuR0IN0Dn3+Lcc5W7s9sU3u+eOfjMdaSN5UqEW6+R7cCZnL+z0ZOl
UaQduq70R2yIJDCluyzQKh6SxXgZ/wok0iX+DxsAUMSsiX994xu3buu4fbncVx+q
Eu0CDWd2hBiHcjVHfoFRjsCplaZwqUlD2ytwDt2DvXD/mDc0fGQRkalmgs3QQjB8
JtJkYSYwJgmNYBImSfudPe5vAhikVW6sTU4pOQVcK8iNDD8oH9F3dqmmN3wHIBOJ
XtbCXC1M0kTraCZoZd8k2Xg/8PwLIHWn8MXDKkGy708GHxs7B4IUZGMgOAkz7dQ8
03i/LcGk4JWkJfLOEFz6N8JPBS75AmAnmEHWg1gORUeedNY2eIAm2gIhsc8KAD8M
92nGghp6cSoKl5y1VWQU4nqzWR3peR0QvoKuzo0Lefby1msXd9rtG41tUunBqq8D
hUKf0bAg3015dtWnafu5BRbiAs6gyfzdQWJWe36QZamK8+6YtPj6mF7PCxXhu8Sp
jFpRcnGMXmcEtF9rWuX75k0zP3OQa2wZ9+IY4cicprZz7ZqjA7f9EfQOivtby/yn
8zalcbZOnH6Exd2C6vuWu/4F7rYuxK6BfAZjYnt8+kULvFmFgm7ecNBK3P+ro4pw
iOtHcgzQvCFmMXCUR1wrhj3AIrOvVh/QSjlyypIRgfyKNH8dd2Vsl++R2pvstWzy
lTq2mCqSCTEHzXuY0NART9DCE+5uIndq5v1exLC1S+yHN01znEHTvphwlw9G4s54
dz8V5JrLh8FQojKIDtOrCZjuQjKHqahRC8srO1paR/ZbRp2NMJUDDW3rMpehmaVS
7rhhpNLyAmu2Gm/+sspWgazwA8KV9KphTU9D1+YsylJKi3IBEaxU182fPvdZ9Y8a
8JKgFQ9q1BP1qt/HG4fW4fb/NdokaKrXtHbaKhLlI5Z36zU+/Xek+ubBpZzH8qdH
23Rsf/YL7gyzY3fL7unjOubwwRmaDtQA87U3DgMqyvTxKAF9dyx/irMHy/L3vMi1
EFsFYeeH8Ib0s2723G0GctWa8WaQDcanou+N9HFRQowciat0wA+Rzuu86HZP6Oc/
kG9RFi3kk4jKopjVF42M0pcsIfyHYKhdyVTlPMMUdapQvunCrr6JxclLXJpmOD5e
zwrjrF+7DGO84tRZLq6hMPaV9UWpVJK9TMOztpvDdkXLxDVFbx4iAT8zZAlvrf/V
zbC/boFBmk9WAnyq3uxWR4Ufk+4soagIBoe04HcgfxaTYcQA0TTOhqqgb//V7XFu
qxPe4jlPkS+f/JNeypE0RCMRPiQGnT5zGkAYuA80PRdM91kAVHY3F1cTckDCVJlX
YeENfDZ7o8abAFIktJsrx23AfTQ2Rgg6W1rHezAKzEz+bPditt1IglLFyf34C6n1
2tBoopmVhrh7PAx6zpqncTDZ5zqok+sqyLt7jdK5dpK/6zKcUHZpLHdBeURXclVs
64YVOejytiZSpwQt/Y+EFSfC1Hx1GsMwYdOfz4O05OqgAirn66kgHxuU1/5HG4cd
Dqm8P78I6oYy1dsa7aH0XrM/3uFYFsyfQK1gScBVK7LJ3QARteXEjM9yuAp5jRtM
IIDUpB1IX2L70WHsYEGggqMLfR86jJDlBS0QeLTaWxjqUGePIRoSbXkVXwOIWxEZ
+0VCV/nayR6L6sqSdagBm9dffxUXrpZAPPHaTBY8SKdCfVvdsPu2ZyDbhsm984q2
Nxnunihq3JONg+G0D3wnMNJU+9KLQbLhPXIL4u1g9Gwq9/j+jvLXNOw3LAHvg+qo
2dHmc61gxWy6KaydfZ5MDXG//u6yry1NVPlumrRdg0hOxm0LBGuV3x7UOJGgSzPk
NBWxAWogFaFVbCG5nSKwDzLjRUNfsLIcTGAF+JDyIzpM+6kjD7H+X7ogduuBC/B/
A7Mn9T2QxEBZibC+kS383i6DVWfekZE1JmeNC8rIje8FPFIuirVqFWGvDLFxpIiB
b00+rcQT/LJQvI5ToR9WmMqfoXXijvRtMTvJv431peiGLHuIFLusrLdaePK9ehT1
Mk0nI8mjACd48kRpfi5qOHwuEZQUPHWPW9pwqrF0WKqGWxt1APhZDNAvsjI9DP1i
hyui1SsH7te8sUshNP4ebWuOuWN9chPfqIYrAfqn43t006gtwZMP9t7pWAnEu9SE
KxwhdCMK2/sgPp61j3toIHypXR0M4YjFgIG38j8Gy5UBwo1qJKm7Gu+987CvByEv
NYWd1kYooS8x5c/u3sojy+vBkN7SDdBbr/g9ZZg/OqnSaegxMLtBLyOEZs4d9k+J
+Cd8jiySskYhwslC00a31f91UqFsbqBAgIErav2JXCipmlnbH99f5Fge08A0f99A
zhsRbnjn5wUvBuvtJTtXWHrnGfCZkKdvoE94EwqgbrqO60G8kxn78pVEed/00+uR
WCvpxN7f6Ngb685GoGF2NTc1p4atTdx3v7n+SFq8PFcRVyE5qV9KGID2V8hT2040
qvUJRVCNBqH06/8ckgv3rsRz7HelqS2diGvMfdN5UN3yJ3s83x5IiHmXWEl1SY2T
KT8GFpBQbaJ0+1wTjoPxRh40Vnnes7Ut2RIQBRTdYFcAU/s/FU8Bkd1HEhMm33gz
JLKA27HyuZH0jbqTfO21Sv1CPIWENSVGmv2QzTim+Ft71/3JtQooK6Ri6916JtTx
fwREy+H1In3frr7ozian4Sh4RaTqDuJGO3vyi+uzauh02zazqYDOssb6cyE4+mO8
KQmqlAD7ptHzCTargBd9yGXxkMH06F7kv3E40xSuxuka7tMHYkKRTUhh//USHU2/
j0f+ieZZ5VmGpuprEALwahM9In0H/xyZi9hb313cCy9lS9wTwkCb3V/9B5w3D4J2
B3e1NymiP7i7jJqoz/eSKOJGT9xh3iTJ09WEFwNe+/LiptaWvnoRsNd5RW52mtF3
jS3JnPaHXrB4csDN7FnO+GP4W4eyFL39mMUJ31Vf5ijdF/oszxmIbLX6O1Pap9hb
yftN7D/JfBU4v+nJCVs2WdwCmjca6rGG6AjIgbyZ6y6Xfwbm706bnNppVQpMAJW+
KijCjxfh1v8IDJqjopVZf9TYInNO2SQaKoOCudtxMrkv0/6z+xS3vebUGmcJpdLp
Y/TvJ/UBEZY+hP5DkttgZa+t5+dfw7a9XstyAM9pGCnkLA8KFcmK3C7U+or4Q3dM
/2PPfw+0nWjrhQpXZxVtCNYUNRrhdVoT0z70+Py3L4aB5ECfcf9tWwnKK92yGlcW
6QzOd8ySdmqNoxJevfIrAdebMzxpRxCrKluPJYlvOh3xDT820fRH+lkz7XLmN0y6
rNzYJtxQEC6c5rK/m8td8RJrnL20PTL75PF5RaxuDzT8WLEvhsy+IpbaycJTPGBJ
wByej5hzEnvdYEabiOUWA8TVm2tT8MPg4A/TSXi53NB3MRekptoYbQHxL3y2swoR
i5GNBAPcF9OM2WXKqBGvJGvzzBZ0gEuSZEaVTTwxnbN55U8DDp7tjmro0PTOOPqh
Fk6CxsPCYZamcymA3icwtFxCyYKapuvH7FV7asskDb6qVZffMSuW384ptdodWLuz
hcw8kkjcD3nCg2FPZRrVL8gQCfoMsIlIoT8QAn0ktJh33L59ujn5fXdho3czRGXD
Fe3YdmVJWhPmi88QyusuDhAGrpzAjyRDDn5MrcRIqDMIgAGV47S6tpg7uEAxuHnW
nnU2d8N/NSkp2jcPIS+9T/MVybKtOd+GLYingpF+N9JD5R2Sa8m8As9UjlXcY3hG
uVJFZ2e3j6D+4UV5QUUvO6LkTtyHCfoQ9oZsVjrXuJd1uRYAOWZ3GS+9sPCbpHwa
avrTYcsxBeUcQxIH+l/cHvnf1nNn+TrNS97ZtesYMOl8fr3yIrIyz5o/QP+Kwxjm
BY1nOoQmXSq6yidhsv9OWuBysL1k+MpKR0B0hKKydFoKAn//38cKPALJYy4kn7qp
Nddl9WxObkybBgqTk0KYC0h59EXBWpfOQ/5Md1n8iuoxnya1ptIdzM5BRRgMnJF4
4dTLgXLMYcI3d+xnJ7dgOFNqn4gAfBQGgwaGZ4o+Op5RJJo9bVaOQhKXL3Fc8laW
QPcdpVpDKSbDqX7NDpoA2mN9J+5haHsP52iW169DfAwthnq7AzfOzIUL5pFDc5LM
L7jPbEdS5IsATMfPmlQOkEKRN8R7VDSeamxM3tPdjLQDE7XxqUa+/f0bhKpxvxvA
fm2ZN1L49JTun8t6/IM7MVBoKxjDfthcu/sH+F672wkoZufWGj2y2Grw9jn/eTX+
X6vSaG0Uee/PIpcfaCVZopu/RwoVcmxFekKSqZqiGU7hzt3rJMGTkbJwQr8ocsbf
z2bUqAWpnC3TXq/vALTekVhIRWqwbxQ0FUwqvb1pST1T7rwYiFycsThxXV1Xeuv4
V30QGtv3pgSTeb1/1BCh+H4HEQ8BsS2s6FKvrntE0WdR00w02C3VRM6lUb9x+LjN
BwaHH65A/kGwz7dTaIIQZW39yfK+M5tLyMPWD/MHbAbgITpTOywsEQmH3jp2H1qu
VkF/cYVenj6GTxpuRjVRLhy7IbPwQvkygyt5HEqJCbO0CoNVABlGoJwPZga6vnZh
X4NKBnogguWInCcfmBgSBx+GgJKpU59ZgbyscNnkolVSI0P2yU7hsTqvwW3l6n23
2uwOKmUqAvkk/fhpHQuglgi1blXMDgQJ5wZHPKV7PsEFD9gkOvdbU14hJ6P5Uzvo
SY1lv041j9TNEyM4Q7V90kfHGY4IEApRki/fBByioAw87fFL4igzhcRsf1N6u98r
pOg1Y2hzUWFAhy8MV3vLy/gUIiSZM3y0vmwyW+ZP+RcmhkgjA32NePcbtldekllk
/V8EXZloXxwpNzyXsKd4Z4c7aODdz450kiZwdwHU3Hatd1LDn8RBnIs7oSHogdGg
1z4pRa786SPm6slIMUs0JnxFlquuknV0P/zMvzrpa8M1cFXYLltWVebXdRaJ45VB
dWrd8ykwITuESZTM4n2raQWOldquTzhwwT83lcxGBeA1cuaKgSy/EqQRqajvoA3H
cTjNQYxodnWnDA9EPuXzwbEvwmcMqAHX1X6t2Oq22y6eDB5GRnq92sYDyfg3birJ
TFQiWgVgoM7f+nUXjCtQ5VfUDhRUEoI2hkpnbC+tpLvxtOjy7WbQJiWfgWcsP5zn
QazlvkDMonqx+pGgaM67zt6czaIu3I/IF6DPJ8I4I7+0c0nS2lzWsXzVDVbhtqSD
/x0SNzPYXgA1k0Cv6UGnYv3bO8/bdDawO4JaZPVqv7K8MnrdrWpSuejibhiYedrX
S5UIhOhGWNK7ZNF6BuF2t46j7aj/CxX2EKGRpZK1ivAlAS0vgVdHMfuD90qPd/Qz
2xsXn0aVHMOwWHklU5hPQWqdDbchsuyR8fl6X5WiL9pMH75M+0vagfuORVnm1ib9
xmBTMAQ+Ap/iYv8YKvfvyC6bUZl/pCC4nfNiulUju9yALO2Wt7wQCSslNE1GL6fm
BSlAaRWc+JBSpdBR70ENkYyoqiNou+TtsZs7gxEKAm7SAcwdvuFqoIbYJn8ho7pU
rFZl2XSJP3OMEKpc9TuDcXLaG3RDpy2JjYyKjoK14Km/jr+dUjTC9CHcJgjWW3ny
zVwhNTnZMcY/YUuFoRRG40PKwNEudGwbjQlqVkwb3X8pqXR6GLFg3fejF1f2ZS0i
+grd5znKyL+Ypa1KfxYAPgVlSyAiVPJ2CtefRX6m5F7cGw5Lvw1fjTIIQHcx5vGm
FrTj/HuBbNhpoSwBCAV/zzDaGa773UclqsXtgC9NDDdli4O8PBIfHVmQ1t4+rYQ6
bZDFEV/Mj0zdvwt+UspEutyONJqYxbDqfJ/2j0abwh7+yGpfGH4KxA5nd4bGuuOp
P5HSdszMLjHskAP5ab6ckNIbxfBmwHNr7Se7LrhI1jnXvChCc+312g+zUL4a9l7F
thVk6iFFSINNKlQdqu8YWGJCOVQhFCNgrQp2LrN+R3LHvjc85xzJy8K45bvDzg42
wrzcvwsKfr1DLmxJ2ei2IAAvfwPyOr8RhWi05s+mlN/Sko23d+Y2jGZT63Z+iqBM
MHlJRQxd6awnmJHXhs21heuZX5wATp/gyzAsXVtAWQzB1DRGyB+0uZ8OLWVfksN6
CE2L5lzG1SWwSLn/7sJcTfjsYcO5XPFRISPGRekmitp/0+LaH8PxR7qlxl7tuP54
G/3JKTZL6ANHYQn7YKMQ1LSBHPNjM+B1zJfjQ4WKZpXK0B8C9u0OzfhYugWz25o9
JevorFx8a4Iaf/rxMJm6H2nj4ussI5bjyEqXj0RMUy0XxtCy/carHLPRBdqAuVY2
IsomEZ1w9AX9L9gmZZTvroAky65rPk4xYspfL54AN5x6KXcqRqG3Y4iOD6bwaxDk
kg9ukUV9lszH5D6ArQM/WiSndeFSmiiypYBl2919HnWYbY+FbrSFD2JY4vKMZTMc
t6T0QJnz86K70xLSiMTe1G0Pik3RWYU7swy57irxWZP8v9nkqbdeUzqvXhI6QX70
Y3zryWWuquioQEK/v9fvhqpLKvd0ff2EDQUlt2nY3OeyOgU4veDiwfZyQ700OQ0U
1XWj2XQEMdPnijseCST6avUJ9pLbLXWDNYFmaIAXIcwfLJF2qhcY7N2D9eQsHTtH
9gn/zKa/XSfbMi8FJDOI21SvJyrJyO4Okn8juv581tnyL+A5+f9VfobYD1yEHv6K
uHQtIvp9/kZOPeTOUUlDygSkX9OYCVdajXRCVN88oK0wXlQ4+WUHMbMLS759WOcG
pHSteT5vXQq19GDoK/AAt4z8udZiGnPdWiul7TASVuM4qyPZcR/L8AvK1yNSV1mm
GkKactLOS5jfUC4VYPLsXJIpa2o09V4N+H6IhB60QrRCjPNiy0CQq2uClzO0cp5a
S8h/bcFTuFHzYqT8DIQyIVhDX4o95nmC6A/eexHZ20Xd5hLKQ7NPxeAyjwB8Led4
va83ZJFqL8ZAh5zyGGvavAepqnZZeqUg9kJjRe3fdmTbChT/2DCh4rjSHaW9ABiw
WiUoP4wRuF6d50C20Sz/rMW/lBlny1oISL2kqQNTlIxIpd2EwbyvBD1zsZJJx2np
wifuYixQNTzUy0l2vJqW8xnsYhRErePlWQb04ecCv2ZUtSGUP2EI7SqF8KjYlitj
YlSyUo1w7aViqClpahHZJjErI20lo/34T4usRQggWIJbToT+7NSl/acd32zjF3QY
S/Zo3KyKcuLSun2w+VVc+ELNoPT4N3rQce4s7S9gm8Y5/mxa70oeYoL6i39buCz+
bqmRfLHTHNnufI8aSvN6HlVCEb3cDok8X2CfsYexwdRXx6ZJot+4MMJivd3NlMhJ
okBs2Spuuj3XdT5kCl8Ur3FDlnwAx41Ja5ZtkMyxT55QtN3RITs7nuTON3ejo+xG
ZJ4Hl8s5W2BOv7JbCoxRH0w3AyJDMHD6W1/+xBILYZnELS1nAIW4TQ1ckH4tkvVP
fORrowVXvM42TDQPNOhx5fHZ7xwZM/ewL1VZaebBECD5pMIr7TH/ZlImV1ZROL5w
xYO/I4MaGvKfg4CWslGZhQDltlouyP/MdmGa2pxJDW+SZgzdZ0knJHW7oUn+SOlW
UziQzeCVvQ5WI3VQZ7CuEaVMsN5J1QqU3bAwX0A1mIYBpi2aCqAKYp6h/Bqi9chs
CjqBaR0wq2QCVScHLpfikNsxSJYQKfOSXy5P9aVhwSc4xyhwEHCXpRA/AvWi90KZ
WqjfoMpnzkTckLlscgX0j2K2EHUBWDk1+KcZwtMOd+g8f2/o1wHsRUXm7nLrnY7e
UXHrTFMqVBzm/y4F7pTrv3g2SpmCxsZCyouCNw2zwuGUC495O6AQIrNXRydnsYxJ
eajHaWB9UMRYj++ZT81FOAFeOUHCTAtOTQt4kF0m0vxc3b/Hwh0BwpLxRsQyI/Zy
JyDNGTpwKKS6ukLRb9uyGDIRzwRMzie5TbxM+c2XHvkFWPlajRtLvDOrzQpD2iW1
N3MWyktuR10XIL+IGofLpu7KxO5H0VEQjtnUBdc0zU22gnFYlHY1cSVgAULW275j
HN9R3KJqkh7fQ79d+XP9v6VFCUKdOnBm4+O5vMLPh47MWRjWUdSPjYN+BuKHJOJ5
dBIEn3ZSWOyIzvQ+TAQX248H1E9EtGDhtVMjrEQw7A5ag286Sw/C/fjYM8lLRZ5R
evDi3crQ6hsxvsWIEx3SRX1gotYJihuzHk4Hp6rWQgBFOwrBbhRqxODZhUnLAEWy
oh2SVYl+jGyFT7XS8qMWRMd5deBxa+VzspsQVKzEdDuvc0AKJ8t6kVrcqwa6UM8T
g7NHkjFXB3nXBYyHCpe2CeqMxSKKP6xjtjoSIrsrRtXhxmWoRCl0wNJJf7GKf2l+
ivEwAFhBb6vgY/YuZe0tJIXyMz0BeaqLdlyWJWR188X3wS36huIetx+SE4tc523r
EO7k+XJtFZxliZf2g89N7jouWM8T4R1fmXtD5dGQKLZp5Y5q9b7Kn+3c8Sk9buXy
I7QGdIQgQZw5T05hrfO21B/lG2yfvoWUXTSMMZBToU3qQg7TkThoqTH3zLPPDuws
3+D+CNEFZkZPYrk2RiTl2fkly5u2tSy8DBPSw3U32twUlMMDOdrM8lVXRLnk9kYG
xlC/f9ZY5lNfxi3LS831uQAISWJHaZhjYSImqUkn+rLaizRTLNnvHqAU1/T8vF+O
UMiBDzZRGyr9TrbApTChcHldo72SXBkVTztB64X/3lFSyXhA57ugps9d7hftMJo1
kxNXXMHtJh3+0NDueqIk+r5bE1ZZxUmI5f2y0lxc+BNv5JiExxgAp4N+IQXk6VL+
yzjLQCPlXKV0PFypbK/W4MXUJ9XaThOYcIgLOX0qeSS4YilN9ZJPpnmCujfLODTH
S9Gjx98vqCEoOpspBvF+29Z+G/lHFh8FonzNplB2gEQUMHQGxSP4qTIZMX6mZp7K
Jyc9r8VcT+8XKC5pY55u1fJTEaotcgg+NOc+XFUdEUIdmgB/svrHR7yf3sZB1qX0
lRdJBB/01eyt3DZM8xRe6BcR3488hA+nnGDTdVdgzFyJ9NibNsXErzSE/Yyr5nCm
h7mzeaNrbJXsscEJUYUxOB4Q52nVAccdEm6fM3p+b9AMW8U3K8zeBvGhCa2ASpQu
CEGPCHO1Z/P8ETxZO60+2DBZ8tbalSS2OoxNpr5TitCW4MrvqGv4dsfXTj8p+8dQ
dct2zgciftO65bxBuwBQKWiIqH15JvZujcWjYAuuoJ0h9vdFpIt5NNlIsb9adS8Q
cWYXRAVGTyxYRl7cDY/5eb21DcWdzTv64tdYcGJdr3lbOqpl6UdeETFLxKxPq1IG
U+uRt+3HiON24Ccv1l97nUxqD8qjg0SPZ4r87EwJv17O+Sxuy8/N4gfjGKZNduGE
VceVw2xnEYzKKeL1QG7hKrnKdB0c/lnHuL3ZrnKky31H5WCau7SWemxPwaPecf4l
IFfuTFswsDjngkRxP318YeGbCVubGO4JMcBf39nnvts7paqf6LQ4yWSiGBcVaVBL
O8qxzvLzEJn+H9mhyMTDnRNIChLV3NazxahJwcAdWuZQ696OYcv2gM1eJvLWREzq
+9ey8zloksmXQc8B0ru0pCloH45A1AgzUGjz2cll9nYlm/gU6quKkNwmWSwnhW3V
ID0vIgrQsN0jddbz7PJv3Adc45fEAi1KlDyfVErMH2q7ngtFFIumEadQ4RSI7xF+
UV9/dl5XZ6j1FC3j005sgtqBppkney83F8+1yiQiFZDgRFaWmmB3jOt3WFpPuLI8
tso6GkyuHMPeU6ddElpGjN7BTZhxGMSxAcDp9966h+GhHUur6QK+PN6zr0NNOF5I
itTltyIpeZN8kqHCemItWnEQNZ9IfRMbzohpQsRzA0dbba2Gtoe8IoKrCHHz/XS8
8AiXc/2NRIBQgBp2sD/M7fbX9DgcODzlCtWXyySu9FN5+9Rs4qwAKRINYag8TxlQ
YcoKYr5Yd4WH+Uo7HAqC+ofEvxmBSi0gMMfMoUOsKLe1euhPW5V7Er6tj7QmHrvi
ikKWJ7r6tPVLT38BLJ4i+Jja9ka5tOlFbudyvO9/In6wX9omgHZQWbDy4LNCASmh
UEVLUinBfvVgupwJg9B8sRMs5YE6feiZd9pCVU6w1qlh/l0poO93oYUwTxMvqywH
DLz63ORsJ/vw2ebV407xRRbwPf5NsqcWggTCY/VRXSmRJt75fRB/mIlgv53V4NRT
TWNGb2gG99RnXzONvfxtfUtk5EgIhSYt3b8bhPu8eHXYjiHXtDXV8P8zXHiLmhF6
SXi2O10GJmGFYhaOxXquWpFP3cel6myGdBOToleKUBK5iuIP2x15ve7XYG2QmtxQ
gIbBHqJuwT+89bB3e9Qeiy/1nJWOVKJsr69YOxfWFAUVYEV9ah4bSOqF/PoaDEdh
WpfVTqz8v53qZKYWtuRBlYSbv5xXe0sYGh+ZwxL6lVAsysZvzwePMXxIM0IVi6op
MRv/mRB/rOvkND76dBWEkQ2W9jx0eM54NJ9txd7xpdXPthbwyqIiV4B+RMVX9FIN
6Jn2DSxPS7NH4GM63V/2f3rDIRCrmMjwwQ7wM8oU0DatKBO9NVfyM/1/0DdMk8T8
5p7L3kQipTl/wIw6JeQ58Pl2pk8niXrdUQbeBSHnjXELvyiVnGDkMxbV6lww11go
+J2afwJCpLBZMQKIfDbSFq9j2lhW6nI2JlbPq081r4BfmVzY6ZJXFi9UsJKlN0Zn
GuCtlDF+hodaru9amhhLvgyE3BbTH+WsyaPKd1cfhSRMnPfGcRKyAiLsJskB2Jkr
ERnzph+5gBOzoUostZSLIKorGUTonPxSd7fQ/sPm2DEUsj3175ibqmjHHVz76mgg
fBQqi8QBvyQupcwS2ireKit+QAQ51p6LtX5vaRhZnUPlUfyc9/rfCf0AExax6Clb
V0KfFvJrATl+T6MyNR2v/lOgOp1VZ0EPt4EH5iCJLi6x/8GLFBiPrCL19NMEs9kZ
IvcDAoQfCMvcnbpmKh2N64jQZ6qJ6TXZJ90Z+TY1V8iq9o4mar9h+ctXc3ebLp3h
U3l2/Xi/UMY9FBq/KdcgwG7oqZ7XJtgVVjAtX4aMw7jv+3EjVpeW1a1wVYgQ33Gq
MSNt6glGwFjLf7GL7YMj67lNUNGKWwkP7ittSq4BSha8+STLAcFGsLEejaSV5JZ0
0Kkry0D+YayHq2/9Jxq3EWDZb6k3nDFbFLwqa7eK8Hu6PJJvoVB0U/J05HQ15174
04XvzkZ6Lx+9CX8eReq/G6ozZO5fWRskjRdHwmSTIPfVcribBVUwvWsZOX5Ci6A6
PpbFimPHEuz3hyzFNgIRw04W3ntKqN5Qy4PXjyVNLcGwuqCIG7aI4n3L23sAboJO
UV/RIXQwSqR/5iXzmIt7WNC8VqIXybG3HylaITIvTHRP5AC55itX7iqJ7biNdGk4
lKPluKosMOV1WvcqE0zmdF+8IivaKteRy/uWd7oUdWKoOIyaSghsbVqQYQ0s/WOw
e4T4s5okGFSTtFii5DlEkDgqwbxRTZ4fXmKgu2qhQocFo37OOEpu6/zgRvKPmwey
BrGC1Y1tgvvojxRVx35nvgq0MZXwndtBPR0CmWpolccOVYatxseZJ3PwstJ0mPdk
tVmVa1F+4AzHuDRublGsp5qdxv6o3OLQVZZkQLEe2FrIPmw3sVhXJf1U3MEnhq7z
y2Ych4EKPmaRTPwzVS1zt5ozwIpEbSGMNLo2EBzYHAKjsQlCuFJGbauzv+hoS9Sk
lIjJWfpXIcHejDoD/urQ8TJUMaJwqzNzgoNaRA6qsP3srbsQgHJWexY093Bh21KJ
bk6cUMbFaVWBXG4u8XUaW4+QWZljx91cWags8nn0OkbtKlwXv+VakTIQoTvMTw47
s8e+EChoIhQdKPnvA+oszeIn19dMYFHK95jhXX9jB0AZciLy987NpJJpsIkpbtGI
D4sUrwx3GXdWegRQFMmNIJnhDJnux9WTpKNv+I3xFfBNvj4QxqaGK7BLhxt8w63h
wQZQ3qnlxBNAEPCP4tRkRAfS0VijbENbgF3iW/atyHCGC/wi0Q7/wdpN6qS25OxU
X9q1PLPQnpBAqOyy51QyrVCdIidOuykURAIupsXTRQ1og5H9qX1YgPQZ6Rq3IzlU
dVX2nkP3hAMFX72wBj6UqvDsXXc47tNiC4KZ9AUKNnUdInUle/5nHCa539+rXcQY
zerPNBmegFAs8Px+s8C2DVjG1xCRmK/CsJBQaM6tQ56nMzMZgsR07H7UDly0cEgL
TScNj0nJnephyt5Uw/TAFG3dcMfKB97LA3MTyIM5kF5JBnQVSBZ7o6p75fYqo4dB
8olljHaRtvnDNHaEX2Ho76e9JsFnU1KXsfDwHu2smLFWLub47o+HecF1ZLuYxLos
EROFlWRumu8d4W5ohKpCVZRTI6NBwVZqIkoqPiDHIL4+uuvkfODxwIqD+NToFwqw
xKPbMkvyvGQM+GvmY3NCpFYkcfDpJr827EMWBENWERd2re05qXQY1spl6V8Vfwu0
i02u7QroxGvoE/cW4iK6krvdp1xg07y9D1gLSLdbaaiKXxzx6390w45JlP9Z0lJL
J93WHVn7Yis4xeAIV+e/sgkfMjbjGo/f0AbzYPebu+nQ4ZWTRjjENLQFdWg0hGZF
jHP5ioLYmJkaS1x+JZYwdtpYwjEC+olddSbAzn5qEpi7JrG1pucL+zzHT49bKsDZ
jzMQSB7A/oLBvtrE5LIX1dcvynS5LzvsGCQNe+PEQdVGU/O8MnOHkNPxaHxIcf45
JNTpUBW+mQgtDMqWVCGOIR1Ddw7Zu5yAq0YMJqBwKZE61mtXZOKZVwCJnar/o/gp
3djCS1gYrMFj5yNp2loPHuftORNzTREPyzMZeMtFs5/tgt3B5FV/AQ5uBvyzi6N/
nwsKQCc3B4rnd9Qfon3SEQq+lesOeDROQqmqoedlE2OIOws8AiCM9hvR+7GbogXT
pgEUPURB2lFasHIAav/2Vom18B28IGvM0J2JZFc6vtytNGoqSGhZHfDhvveIzErr
/zjCf7JnqdldWFNl923eaAwWLHH9MIhO9fM3ZBivAoAoM7i/zf7sfx27sijjD9pR
yGVsKd/yMMZnc4I/W5tk2wpsulaYY2roTRcSroWRuE4bZ0ljua+KQmg9Cy0RL7tI
e1gr1dho0RI0zLBn/J11OJtIm08bVO5QLrajOt7yV8dAjg8MoCGGIeWrG0MpdIi6
R2dylW2QrBhiaVUgBn6XhVu0M8UmkCYjWGtD0x+8XurzbxGabfrNIap0bWpizqg6
bDCo6mzg7xH9Asbs5QTUypjJI3hQ3jeN4hnSfWznwhWt/dmqb5f5VkcNW4IwKxTi
kwBg+JNLSg6ZAv1ZxRmWYpXf241N5ed+5dFm8KKRf/rWGSGJF99RuIitOLwuFHtL
HGknORkwVHeTL872r/df27Acch5vSDEyc0Pv1Gk6Zo58VB3RFszBWGOXIwG9ilom
0WArQLcKX8fdd+0LzInn2abxCRwPCowY5ZM3ayvy0J+VcjQYC7QkCUeI70ZJaTsW
kr0qCgpPrLKAw/vYk29FDyQKojImv7OL7n5oWyrmnD6Jbk6qJwImfEdzrijFwJ8U
ZHuKr/bLUliC8IkVc1OeG0xaWTfA7N594rs11O6xmwVN2NhezlLHJfBiIi+UYalL
t6XDMDTliQcq/VoZQSoQmYcMYxtbYJ56s75aTTfIMymSJ406TRAsshNiV/OFUNwp
cNsHSc+cpKw+QT/n+IejA6ZeR8Ri0Vzg1spYFxgbrrbSnEe/zOpGqkcn4C7HkMbA
GcEbljGV3uzRFYUHyPTv8VHi1FCimN24oma5jqtvvuoaz5tzhI02rawRvwrNbNpZ
KjIHRMGi8bLD6UYSyH/WY67wSYVZYAIgp7UCUqjiiJ8BFqZifd2aPiDnaIu623lo
xRY4qJPhaDHyKpiQxgTK407C017U8tpAZQaDyYPHsIqww6x38xx/08bwguSMy5zP
hmIc7Xk6fdpYeN5ZNfF8KJYc34n97qClJTtDp8ZfXyw/qtGZ627ewagvpG0EqE63
We4EaYulJgGje1To2fEBfyat0PFgNrdpg9PXBWOAvviCW4ORAK/csM3sEG8YiD0i
BJlmkfA7d4IQexeJvyVZKuTp1P8DmqSONMlhUil2EIWE1WpX8MhdRznQVKRZnTVX
BFhtCNlvg4rIhJGSia2sIz6vTafbSklo+aOvq3e6LQWNBprFyz7f3zSGK/hKbfVt
dSuCEtMJXuw2p+T2pys/7UCfZFyNYk3/vNuoMlBid2kFYlmOhkStnB5Cj+kqp++W
QxZshE8tuZmLk4rq1LL+tXxtCFD4DRekWS8t0+hYUBykT98B81oizD3QbajPwBso
xoelNogmnk820b4hkifRT0Xmy420xnSFWCa5la3ZIrDNpBjgkXq2LJTigQ1hhui1
+PuXWz8scqTXXsHix3ynU6ShEH6DlS/aFyGahtMy6npwy/8wda7JAbV39KSmCTcs
kC1UwwBbfZHKRwNTt6Y40YfSH51dmrRYxoKXwTgdTpiwtCLJQw24aow65LyHcGyp
FjoZQwtklRMEr/0lS+WJxKu8q0R53A8Z5i6Tbdsss4SCGkhaRtapgnhpgefmP560
5L+IGCWkxfSzTYTgCfMIE4+f1FeUfodDXPymOynxnGlPlr945/svRLBqBc2uDrgm
QiP2hn7qHcalWjMZmt6JOkL9zSgftOfK6ybo52uMan33UtAPKt/V6Kk0XWhLJD61
WboRWbu2ny42cLkG34rcNIbSlVUbADbhjhsJ/ZuqtFrjFprNXkjY64bhjKfRejWL
7EgOZDKukUSa4oNSeDLNqgJp3CirW1v3pOKns0ets7QcHcJARXQhrbYn20vRGusY
i4B4weUmBv+nAMA36lkTpd+zdWLehxNVl1hScrpoMpaKBL9A/YYnu7yGE7btf+3v
3zrOQBt/xZCjRo8IAVPrnlgFRFt08atg0ZMlwwlRhXSanaSfjOwtciVLmM7d17hs
dMNhPa/iBT9FWs/vYlwGQxjV2WBEymD4Sd+6EHa5wA84zEbvpFdojatbpC/iBoxf
PnXTwPSRJaUCMEmmKS/9rzh4gLSZ/kJHDlCvWGJJZ/cGFttmg/3BgHexUpGTBQPS
e4DKtH/okgrErrMMqQOVdRdI3ewQoBSrEx9SNao8YgOkQc1OilHJdGltMWNESVP7
Mv/Xl164zOwupIMUERAxblhxJ8Fvwb4JBtP77AcoxGe2mzEm2NZX8183Et28Zi9m
PkOKIEcyS96XEdtNNg1l5SYVDL2yh/fOHzgli5ilkIncXe6O/hz5pHccowGH90B+
VoMCUciGzlreiBSsbWQvWR413sMVSYCeN9NvpWnsl4deX+/2BQWcbRWXahyUhAd6
ZrK0kC+Q/h5FWOcNwr/jCFcDeKU8vEkpnS8BqSe785j5hmQ7zEYcl4MpLESlfbuw
58UR+qZL8fzQ+qH11gKBLoDJ3/kR9Xj5jsuQynFTbBmfn76eQI3IqjtwrK8kt7E5
NwDtQC+kjXHCbHfcppkkDHWaF/da0a51k30Wt/BaaIFUxrUpHSQ3QyYqDsDXdmNm
dcSKOTuATVXCHtMBeeJ4/moZxvWXNe9Vw2DrtA+kdMoADfTaAUMSzKWlZRuX03xZ
i4TBcY1BAr/NR3jAsGQtvY4ywmpTScddrQSMR6upiO1+UE04Jg9VdtzTQK3M2E2K
CJy11eYPwKoeAkt+KBemrWvDTqlPHBX7bvKGfsDK01q55l1yke+COEico//LHBZG
8rZ6qkz6wp9SsvvE4+rTl7ndl3I3yeUUTL4feyyivIvAByPZTmXY42sX6D5K8KjN
eS0cMf9J0gRtAQ4zwT1qIeeA7Ml84QKbWMrM/YJqiKGVcwEF10Q4MBglYVAeiM4w
JXY6XNwCaUVc/gBtHDCjfoeiMkFrjU+cMtSsIMxVUAmjtw7l22i5Xfl5k1yGWtYo
+kLUUjbvI5zLzc7zV7Q7FLuLzivpm8vFZHOpWapyklyOh1TYOnK6ri1/BqynquwU
fMbOjVxa6yduGHGbNR8nT2RtqsEpkIFzwRxsUhhNi/bpX2l89EM9bxLewgrKdrMz
iVbnze0eqDnJmL/67UDgIpZ/1N61usl+QiKn+o99vDzLcL7cMGCI3t0ekm2sS2rO
2eHBZhfIuIrmsbaZFWJX97OjOPcPuAkAJHoQoVxH/CUpUYjjbzww9rxCwn2LaTyf
77FNDg0VcH0XhoMkPTbqU7wA8v1pG1OWIFkCICE38kiith1x+ZW5cc20uh7jrsVW
XnndcxwuvDsDmHyUsWYvovfaB9TAkOGaqs52iPTV5RcGFHQdvfSukBg2bwLSgEFj
xwQDx2gIhx0+ebXdESFWr4k0Kpbx7OJB/bHscDJR4RKQQ2vxRhEy41UMvP/a+tNe
gGvdAAvPA7bTvl5uJlIJ2bieQDsUFatdjBPQMc3Y+V8MX4DfW2nhe3z+C0Sn3v4y
a6arHjiwOByjUIC3+t2DlmGJJ0RCkSWyHjg1U247NQRNY7Um4jATff+alhAfOZ11
hVEm3UU2locbTnNpIKELuLWulybC/oTExVIroSJPLX9vavp1j3/1fuApv8tjiZLk
uAhR12WS9rWVq/4PY4J5nKM0Bj6qxcnXUkctZtjqqIET3jpFWX/BLalp89Krh2ib
2OUtz109UqZoAetkCWGzAYpRqu941sRgReeVIEecaR/rWOOaNsTffujxfzSZpnzQ
L30ndXpr51HwyZaPqvUtQlGIE/hPwNJNedsiwi7PaPlfQC0kSAKiBzFdy9zZmO/5
XM6rw2oBQUZAmulJMe3NxHabV++x6F/NPyiKYAx92PJQJneV5q9tdZVrdKykuWfB
fbIilwkgD84YnBZXifl7nrf0pQAoyUY+7nHboEBDVJ4wfOcI+PEtzQI/8aCjg5VW
nBJUyLSeJfaFykGp8Qfs734PgQriG8XxWQBiVoi8uafuW37Koki813A6Qu4/kLVA
GiXE5S5A0dt3T3bTWmLyFmymc83xpYKMJLTPoK+ZIauBxQHEhgoV5UyvKxrdCTyf
YdrVKoeL+8ozgRP/XN3B0GhMZ2XlxpoXPzWd8oMzf7Ij4DwMRp8/et38QF/f86Ln
0SLvO7D16+E9DgSrpHuMkEI4Sc8AtQ6TVNb5Jrsp0mFPXrqoN0o6oxbNaFiWq4KA
ZpDO7KK9544PLkMDiwsiJECXUv22Vh1DrIUTwEcxUA0LsPkv8bnqmo9XYvh+JhqV
5wdZ4mpPDXCg5b63szTnhqY2S6ho9SD8Z2zGXq0K9vHszaWt8U5LmVvVZ0Uu+5wj
20JwPgSPZZ5/p7+7sX/7ktdvippQf7d4Vbd6wSORnU2qQBxboo157oboQk/UVdki
aijuG7zJGTJWPyaawlQ2lJhpXsPzn4KynVYpSmpFD9ykRIhsVya53MavaftVL1FN
D+KBfc+5PiAW3S94lX7jsEHwo9GB+WFa6udCb/hB6i9R5dK9nk9rxxbPLZCSte+U
6IX6Qu6Uhvegx1TFP3Md6Y1oObpjXfq35AGwIXqjiQbdpLb6ddkU6yfJGs1zrtyq
FuGesMhZYLnAZWq8orA9L59cEs1V+c800UC1WGCawst2EdGAZLyYhVpMSm/1/Jik
d5Dm+DzxNtZPwVyRMS26hcAOyGYlDXvOf87EeHhoI8lEBgD5WJe7VKtPxORiFuG6
z53zQ4ZIBuRMyujfav4j4raowrA4ZqcGATFV6xzw5bFk3YegaQf2NxgfV0v1mnyR
7Lr0pBDWzPjOrQ8qzvMPIO6HnC72iUmEbE7BZ4iH0Tgap9Q65FZUV/VBN8AZRdhq
R/fa0IvTs2i0QQJGqFIV2BWnkyWqMN5Fh1wJnqlGOgfnneZwXP+y6OYuOPoQKVQC
yfnXkUrLoUT85od7anhc1okJjDnVck3swTF9haODXFkFBImclVAP+sknHF1kyD79
8Br2fqwxzT6OGidvvgU/bdvzs/iskYF65kdmwAyMCh4msi2InO6Xw4iGmM5jhM13
Wa5WmXMxl3hJFkyNtc8yZmEZtocQclamv74MVOEvHc+/t9d07mNPkPPZuAawJRNL
pibyjgEq+WpKv57lx/kfmIfpHwQptOuRn1fyfswV5EN7qmPAVY31fbk3FN2FYs8M
28GDi+RxtIehC3aguq/McI7Ku/Lp7B51YJTf6TFnkLw/YZb0Dh/DT/t6lPxYMYUO
GhI0axF18EfUf2KgJFS2Yhjs63gPZ9YncCHs14TXN1BxUMCNBKCpRGZoaDrV062K
fD2LWCV6Z3AD9xawghce6Nwtzv12RbUA9Cn8DQg3rQefQOf7UAokbnlkM61S4LT0
5+xfegv3nzedlIYX23sDu7/rrz5mhYndemlt5THXKX1VVNVvrhewc7WgUm0G62b6
FqzIIN9GCo+jyR6W2M+HUjSeyCkx0vKHSqLTQI95+9j1Qq6R7au1y7a1vtM/hoAG
ZP70tsofmiAiPPNDQRWdlWOSiMFba+/cvvOiFB37sw/7OpgqoJoksAMYrdd00QG/
U2smR8WeSlNni0hH99kF1ViYrNhmwfPCmxEj1E01zjfa2s17OOSZVM8YPZbzJKaF
3+jhEXeUCrSaXcvT2ywCUgVsWAqA0Qwpk+t8GDwC6j7h1F4HGWAaelyWdT5iPYF0
8hXlsW//QPm4q2Wyl6t+80Sfvm4dXPcIdpgiHj93T1iIE+mbvioEl1LVjvMszPnI
jWw1SfJ8VAaAgJcHI0e+bG7YDfY5gtVGJwKcxjo5TBVMV3LNbqdbsBm6f1Pw6esc
gKfsOJYfjC7LXhddZn4Ugc68dkrvCzCvmfYvX2e5nOAxCtlemFdATYQUGsOw8Jp9
zXpWYDnSylp5loP2QG/SoWZa8Dvjau1G9KFq8CUk/AO0W8FJYIAOjgV8Ad+VuURm
KqCotSgafGTtsQmKN2NfNj8wwz2vqoyw1/Gyyq5cSfy35wMLtyIzjSikC1ljmTMv
b8O44oLV9BZvLe4xAti2knCKPQn9S+gpmmQ00GcZv3W4HmUfADHrnDZGK+GPVF+/
V6azeu2PKY5EXqbRyna/233jX40KOhP3EL3gpmiIvZDY2ouUKFJfSZqsC1KVcp9C
LgU+ebpcBON3SWiYC3PsY/4cSaYwKYKUbUb7Q/AVZYOfJSCsYAgrsL5OqQvgbNJu
2pcsJi3+mqNv6vuB5gzx0YDRHvI+rajMjmZ48J1s6rfOb+jLY89igHGM1aYsgA4Y
EpotX9U1C/gTmxEwh4s5Gxoh5vx7REANJOIgY+XoZ7BTpq0HckUV+zlKfx1pgpbM
wupPE5mnQFStArjj6BKNQDNgwU/plVCfl3aEqKs8bEh2JZT9o2pSkbco9MVgxXKJ
NgENaKvbDyjzJymEAympKinJexES8OwUIYdGb5qPv4e9KppgVo2GH1XdSF6ynyMy
QNfmA7hA10lw+PuKD+wAg4rqSfmEDUFoRmhKsGfYzutEs+qYla36Y7s+1CVIh4uM
PDgvrZ02CdP7UoGqDSt8/ssDJGq+cQRFSIEM29z4ydt6shQN5vW4rMUOwLDRYtKN
f3r8Z1Tg8iI9SUWyYClYqoHBQ+Ata1zrxW93CJcINVZyWNlsHi1nTvLD4vWeWe69
9Fx2j1yniE9Gd6uxHIZkIu1MNjAyjiKHRNfT4aKvluPUFXmmTGxW2LYotTWQfU9z
caF0GEigVIPhGKRgz2+9mu/Kbc0MR9+Rbv0vIfB4NPW96yPUNm7DEBCmWNxB/o8q
eSYN6ThMezHPUppTggOdL8qkTLNZ4oLk36xg3P7hLakcR2VBODshVrOhW1aMn6oW
4PVsDa+kOg7FqcPxGyICix0uFYBK9gBr1lnNomST6VTHDwx1MDPk4g6CnsmlifiL
csOQbjgV0hSxJomGUracCSvcc//LB0rlD85DC7bXZv7txvyYzJFtLziooPnsosza
rj2eMj3Dv7P8JFT77Wnd4r9uONbQJbxI6y1gkZ2zDjpdqc0OLOphvWSe/WuWv9zN
L9F+YeD9L98SvtzqOpr80WDR+ZHEEbK1EAgdXWOvfM5htetoVf9PB70ChsHRLv2n
4vaecr+fi2bM93ryp4uHWIYJhcDoxtXrBeBHTssCbkOb1kj2fdXLhFmAcxpOszTF
QeZoOjwFm1xRdw5u3VQ/xUSx49RI5o4fHpWmpQ18mCBwAfks+IrAv5Z49qxzqk5J
gt4grtxBIbfGeDk2AfzUDh/oXG24DTOlBDWhBsyvNRatjir+993xyC6kJ7Zt8Rt6
fLioi1GUFkUUlL3yARE7yadsmqwMRBWPnd5tbWjscO34cOoF9VklUaKzdCUwjZ4d
oMZUPLxGQrMFgoQZ+2P5Y+c+4ZzMoGIa9lk383B4il+UhlUOe7xYQ6yXE20u6/0y
Vih9JwaqH1jcRMEmVzP1NykKJr9GItU5j20YZlgGewqsvI50NJQJtu2OH7PtDzKW
JcbpdbT0rdzM5qar6M7VSEFMp5UQMTrxs+LKLCXFKA7f+WmKhTCpIfy4LJKSYJK2
dPY2zi8RRV7VwJMCnVq9h5LG0QfVCvOUxIXPyFUyAhUyj3B/T1aENhNbfqS3+NkQ
wl2ziBnt+bgtdLsklR+rFwpWPCfR7x4k8UOirsI7zVMPbQ6u6W0hSxKf8FPoW2x5
7SGBFa49SYhwF+FGAVVk12LHmO7D/9mTycQyboAHTeYomNYDaODaW95sRPomys3I
NnQP/8KH/AbGaOFy2LMI8xxn8HsxzoJC1gq67ageft/mK2oKDjTOAJ/JvLbAap89
5kEWesYllxaJ7PsQlGOzs1d7osk4L3XahCsK21s3bE4SAD2K51cfpOW4X/iQX1sg
G14AevKs+4VPJ/Z6qKgtHdulX0rdNjyRC66DxPPv77cL2/fAawcBPapJw9kICYhz
7TGnSANkwBxucSjkMH2fUFbjWBnoR7KDrio6rnbukJFDkD6DfI6xLLYwV/C6X0zH
eIbK4Rk6/3ThlyKbBDCnfNGZWsIOv7tSEC2RdXB3hLAEb19Qfx4Jf4HcHWrRhndB
vLMl7wfsTtDzK9DKJjat1J1CvI7VyGIjy1XkgT6qWO00oP0C+7ViAriBNquFbnGA
7A41ZZ4HUMjnjcZAsj90E7qnS2sqt9heFei2148ap7llMNDc7eehES4fZZo1+kiP
5pc3jOGyYQt5xttw09gHZQhxWCZbBPKyoRSRdhZI12mHScNXx0BdVmxiWybxThA+
G7Af8L1UkkjJQw0UObGUEsx+PdHmQ3tMQ6D3bwPOYuM/3Bln1JScCm55hMQrAgzu
8Fper0V9qlg/DjIlxOb/+AgMPYc/z+M6PxvXfl0s9No2Eiuk7KB52GkE31ibD1pC
g/oc5dwEq9ptG65w4yF3vZ95gNhOYT6LXnkP8gi3MBMACh0KyYGdfS5S5q2kez3c
KJCvL2NzuiyL6Jg/D9BYSugFIOlHOYaSerijQsOmkYUhlVbmzRSh+KucG2MTtUfS
xM8m08gRZPOqRZjA7moXSNrLx9OHaq+0xRIZVdRL+IeOrUfeHf+6wi/2R/cEstFr
t+MI66A946YRye3eCKSaYGGuYykuyRAhCFqnESx9/qCd/rAX90nFSMQmCIZnhTFI
WPXtFnP493lHkbT9pb2X9gUumV3V5iIEO2A6vvpag0okR58vyFhAv9uNEG6E/OVs
4ugn0pd+uN4QjEYgVlKXM1BnqK3LCCD/41rd8aijQynn1W9GWJCZNbtf7BhRYLaU
W1L2wxuFdMFFByJoSRMTpSJcC2hCLGxY88Nd3EOdGwRpANZXhmb2vprzTkfhdNaA
7jP1ba4EO1Ln5PXGaZKNf1+kEppGuaKnF3oQ83lFeQh7ticeU4bM3HlPHPtyW0aB
fJkIOqwAU9tOSIFMoAO9+goLbPccq4Wxc2FgIq0GrcN/vcAhRiKBmPxnlUzZJDeC
p/LfC/J8ga96mUQt8oOnCmQYL/j4RBSRGdDJT/HlNNk=
`pragma protect end_protected
